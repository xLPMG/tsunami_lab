netcdf tsunamiNetCdf {
dimensions:
	time = UNLIMITED ; // (30 currently)
	x = 50 ;
	y = 50 ;
variables:
	float time(time) ;
		time:units = "seconds" ;
	float x(x) ;
		x:units = "meters" ;
		x:axis = "X" ;
	float y(y) ;
		y:units = "meters" ;
		y:axis = "Y" ;
	float height(time, x, y) ;
		height:units = "meters" ;
	float totalHeight(time, x, y) ;
		totalHeight:units = "meters" ;
	float bathymetry(x, y) ;
	float momentumX(time, x, y) ;
		momentumX:units = "meters\000axis\000X\000Y" ;
	float momentumY(time, x, y) ;
		momentumY:units = "meters\000axis\000X\000Y" ;
data:

 time = 0, 25, 50, 75, 100, 125, 150, 175, 200, 225, 250, 275, 300, 325, 350, 
    375, 400, 425, 450, 475, 500, 525, 550, 575, 600, 625, 650, 675, 700, 725 ;

 x = 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 
    20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 37, 
    38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49 ;

 y = 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 
    20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 37, 
    38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49 ;

 height =
  // height(0,0, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // height(0,1, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // height(0,2, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // height(0,3, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // height(0,4, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // height(0,5, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // height(0,6, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // height(0,7, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // height(0,8, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // height(0,9, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // height(0,10, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // height(0,11, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // height(0,12, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // height(0,13, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // height(0,14, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // height(0,15, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // height(0,16, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // height(0,17, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // height(0,18, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // height(0,19, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // height(0,20, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 0, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // height(0,21, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 0, 5, 5, 5, 5, 5, 5, 5, 10, 
    10, 10, 10, 10, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5,
  // height(0,22, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 0, 5, 5, 5, 5, 5, 5, 10, 10, 
    10, 10, 10, 10, 10, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5,
  // height(0,23, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 0, 5, 5, 5, 5, 5, 10, 10, 
    10, 10, 10, 10, 10, 10, 10, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5,
  // height(0,24, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 0, 5, 5, 5, 5, 5, 10, 10, 
    10, 10, 10, 10, 10, 10, 10, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5,
  // height(0,25, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 0, 5, 5, 5, 5, 5, 10, 10, 
    10, 10, 10, 10, 10, 10, 10, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5,
  // height(0,26, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 0, 5, 5, 5, 5, 5, 10, 10, 
    10, 10, 10, 10, 10, 10, 10, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5,
  // height(0,27, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 0, 5, 5, 5, 5, 5, 10, 10, 
    10, 10, 10, 10, 10, 10, 10, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5,
  // height(0,28, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 0, 5, 5, 5, 5, 5, 5, 10, 10, 
    10, 10, 10, 10, 10, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5,
  // height(0,29, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 0, 5, 5, 5, 5, 5, 5, 5, 10, 
    10, 10, 10, 10, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5,
  // height(0,30, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // height(0,31, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // height(0,32, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // height(0,33, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // height(0,34, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // height(0,35, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // height(0,36, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // height(0,37, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // height(0,38, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // height(0,39, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // height(0,40, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // height(0,41, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // height(0,42, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // height(0,43, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // height(0,44, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // height(0,45, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // height(0,46, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // height(0,47, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // height(0,48, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // height(0,49, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // height(1,0, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // height(1,1, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // height(1,2, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // height(1,3, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // height(1,4, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // height(1,5, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // height(1,6, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // height(1,7, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // height(1,8, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // height(1,9, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5.000001, 5.000003, 5.000003, 5.000003, 5.000003, 5.000003, 5.000001, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // height(1,10, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 
    5.00001, 5.000023, 5.000029, 5.00003, 5.000029, 5.000023, 5.00001, 
    5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // height(1,11, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000005, 
    5.000022, 5.000071, 5.000165, 5.000208, 5.000218, 5.000208, 5.000165, 
    5.000071, 5.000022, 5.000005, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5,
  // height(1,12, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000009, 
    5.000041, 5.000161, 5.000472, 5.00103, 5.001293, 5.001361, 5.001293, 
    5.00103, 5.000472, 5.000161, 5.000041, 5.000009, 5.000001, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // height(1,13, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000013, 
    5.000065, 5.00028, 5.000989, 5.002667, 5.005479, 5.00688, 5.007271, 
    5.00688, 5.005479, 5.002667, 5.000989, 5.00028, 5.000065, 5.000013, 
    5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // height(1,14, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000016, 
    5.000087, 5.000412, 5.001609, 5.005196, 5.012874, 5.024823, 5.031068, 
    5.032917, 5.031068, 5.024823, 5.012874, 5.005196, 5.001609, 5.000412, 
    5.000087, 5.000016, 5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // height(1,15, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000018, 
    5.000104, 5.000527, 5.002232, 5.007843, 5.023126, 5.05233, 5.093832, 
    5.116333, 5.123362, 5.116333, 5.093832, 5.05233, 5.023126, 5.007843, 
    5.002232, 5.000527, 5.000104, 5.000018, 5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5,
  // height(1,16, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000016, 5.000111, 
    5.000595, 5.002696, 5.010195, 5.032046, 5.08562, 5.174296, 5.284347, 
    5.345138, 5.365025, 5.345138, 5.284347, 5.174296, 5.08562, 5.032046, 
    5.010195, 5.002696, 5.000595, 5.00011, 5.000018, 5.000002, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5,
  // height(1,17, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000013, 5.000091, 
    5.000609, 5.00287, 5.011568, 5.038834, 5.107607, 5.255316, 5.45458, 
    5.654781, 5.766831, 5.805127, 5.766831, 5.654781, 5.45458, 5.255316, 
    5.107607, 5.038834, 5.011568, 5.002866, 5.000595, 5.000104, 5.000016, 
    5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // height(1,18, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000008, 5.00006, 5.000425, 
    5.002811, 5.011596, 5.041329, 5.121252, 5.288161, 5.587032, 5.889495, 
    6.114048, 6.247925, 6.296353, 6.247925, 6.114048, 5.889495, 5.587032, 
    5.288161, 5.121252, 5.041325, 5.011568, 5.002696, 5.000527, 5.000087, 
    5.000013, 5.000001, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // height(1,19, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000003, 5.000028, 5.000218, 
    5.001533, 5.011003, 5.039038, 5.121291, 5.303221, 5.596775, 6.011393, 
    6.30257, 6.444544, 6.550306, 6.591668, 6.550305, 6.444544, 6.30257, 
    6.011393, 5.596775, 5.303215, 5.121252, 5.038834, 5.010195, 5.002232, 
    5.000412, 5.000065, 5.000009, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // height(1,20, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000014, 0, 5.039814, 
    5.109214, 5.288445, 5.596817, 5.95014, 6.326973, 6.498679, 6.541141, 
    6.600243, 6.624728, 6.600243, 6.541141, 6.498679, 6.326972, 5.950134, 
    5.596775, 5.288161, 5.107607, 5.032046, 5.007843, 5.001609, 5.00028, 
    5.000041, 5.000005, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // height(1,21, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 0, 5.108829, 
    5.260567, 5.588036, 6.011554, 6.326994, 6.546953, 6.566364, 6.535832, 
    6.558554, 6.576564, 6.558554, 6.535832, 6.566363, 6.546951, 6.326972, 
    6.011393, 5.587032, 5.255316, 5.08562, 5.023126, 5.005196, 5.000989, 
    5.000161, 5.000022, 5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // height(1,22, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 0, 5.226802, 5.467532, 
    5.892158, 6.303021, 6.498741, 6.56637, 6.621973, 6.765517, 6.920608, 
    6.987292, 6.920608, 6.765517, 6.621973, 6.566362, 6.498679, 6.30257, 
    5.889495, 5.45458, 5.174296, 5.05233, 5.012874, 5.002667, 5.000472, 
    5.000071, 5.00001, 5.000001, 5, 5, 5, 5, 5, 5, 5, 5,
  // height(1,23, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 0, 5.378377, 5.679589, 
    6.119381, 6.445471, 6.541272, 6.535846, 6.765518, 7.138705, 7.442398, 
    7.559381, 7.442398, 7.138703, 6.765517, 6.535831, 6.541141, 6.444544, 
    6.114048, 5.654781, 5.284347, 5.093832, 5.024823, 5.005479, 5.00103, 
    5.000165, 5.000023, 5.000003, 5, 5, 5, 5, 5, 5, 5, 5,
  // height(1,24, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 0, 5.461733, 5.797845, 
    6.254579, 6.551452, 6.600401, 6.558572, 6.920609, 7.442399, 7.841739, 
    7.990802, 7.841739, 7.442398, 6.920608, 6.558555, 6.600243, 6.550306, 
    6.247925, 5.766831, 5.345138, 5.116333, 5.031068, 5.00688, 5.001293, 
    5.000208, 5.000029, 5.000003, 5, 5, 5, 5, 5, 5, 5, 5,
  // height(1,25, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 0, 5.488677, 5.83798, 
    6.303374, 6.592873, 6.624895, 6.576583, 6.987293, 7.559382, 7.990802, 
    8.150589, 7.990803, 7.559381, 6.987291, 6.576564, 6.624729, 6.591668, 
    6.296353, 5.805127, 5.365025, 5.123362, 5.032917, 5.007271, 5.001361, 
    5.000218, 5.00003, 5.000003, 5, 5, 5, 5, 5, 5, 5, 5,
  // height(1,26, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 0, 5.461732, 5.797844, 
    6.254579, 6.551452, 6.600401, 6.558572, 6.920609, 7.442398, 7.841739, 
    7.990802, 7.841739, 7.442398, 6.920608, 6.558555, 6.600243, 6.550306, 
    6.247925, 5.766831, 5.345138, 5.116333, 5.031068, 5.00688, 5.001293, 
    5.000208, 5.000029, 5.000003, 5, 5, 5, 5, 5, 5, 5, 5,
  // height(1,27, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 0, 5.378368, 
    5.679588, 6.119381, 6.445471, 6.541272, 6.535846, 6.765518, 7.138705, 
    7.442398, 7.55938, 7.442398, 7.138704, 6.765517, 6.535832, 6.541142, 
    6.444544, 6.114048, 5.654781, 5.284347, 5.093832, 5.024823, 5.005479, 
    5.00103, 5.000165, 5.000023, 5.000003, 5, 5, 5, 5, 5, 5, 5, 5,
  // height(1,28, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000009, 0, 5.226734, 
    5.467518, 5.892155, 6.303021, 6.498741, 6.56637, 6.621974, 6.765516, 
    6.920608, 6.987291, 6.920608, 6.765516, 6.621973, 6.566363, 6.498679, 
    6.30257, 5.889495, 5.45458, 5.174296, 5.05233, 5.012874, 5.002667, 
    5.000472, 5.000071, 5.00001, 5.000001, 5, 5, 5, 5, 5, 5, 5, 5,
  // height(1,29, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000013, 5.00007, 0, 
    5.108382, 5.260472, 5.588021, 6.011552, 6.326994, 6.546954, 6.566364, 
    6.535832, 6.558555, 6.576563, 6.558555, 6.535832, 6.566363, 6.546951, 
    6.326972, 6.011393, 5.587032, 5.255316, 5.08562, 5.023126, 5.005196, 
    5.000989, 5.000161, 5.000022, 5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // height(1,30, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000017, 5.000138, 5.000946, 
    5.005786, 5.03459, 5.108321, 5.288314, 5.5968, 5.950139, 6.326973, 
    6.49868, 6.541142, 6.600243, 6.624728, 6.600243, 6.541142, 6.498679, 
    6.326972, 5.950134, 5.596775, 5.288161, 5.107607, 5.032046, 5.007843, 
    5.001609, 5.00028, 5.000041, 5.000005, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // height(1,31, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000005, 5.000042, 5.000306, 
    5.001886, 5.010614, 5.038951, 5.121276, 5.303219, 5.596775, 6.011393, 
    6.30257, 6.444544, 6.550306, 6.591668, 6.550306, 6.444544, 6.30257, 
    6.011393, 5.596775, 5.303215, 5.121252, 5.038834, 5.010195, 5.002232, 
    5.000412, 5.000065, 5.000009, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // height(1,32, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000009, 5.000072, 5.000477, 
    5.002755, 5.011584, 5.041328, 5.121252, 5.288161, 5.587032, 5.889495, 
    6.114048, 6.247925, 6.296353, 6.247925, 6.114048, 5.889495, 5.587032, 
    5.288161, 5.121252, 5.041325, 5.011568, 5.002696, 5.000527, 5.000087, 
    5.000013, 5.000001, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // height(1,33, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000014, 5.000097, 
    5.000602, 5.002868, 5.011568, 5.038834, 5.107607, 5.255316, 5.45458, 
    5.654781, 5.766831, 5.805127, 5.766831, 5.654781, 5.45458, 5.255316, 
    5.107607, 5.038834, 5.011568, 5.002866, 5.000595, 5.000104, 5.000016, 
    5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // height(1,34, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000017, 5.00011, 
    5.000595, 5.002696, 5.010195, 5.032046, 5.08562, 5.174296, 5.284347, 
    5.345138, 5.365025, 5.345138, 5.284347, 5.174296, 5.08562, 5.032046, 
    5.010195, 5.002696, 5.000595, 5.00011, 5.000018, 5.000002, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5,
  // height(1,35, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000018, 
    5.000104, 5.000527, 5.002232, 5.007843, 5.023126, 5.05233, 5.093832, 
    5.116333, 5.123362, 5.116333, 5.093832, 5.05233, 5.023126, 5.007843, 
    5.002232, 5.000527, 5.000104, 5.000018, 5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5,
  // height(1,36, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000016, 
    5.000087, 5.000412, 5.001609, 5.005196, 5.012874, 5.024823, 5.031068, 
    5.032917, 5.031068, 5.024823, 5.012874, 5.005196, 5.001609, 5.000412, 
    5.000087, 5.000016, 5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // height(1,37, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000013, 
    5.000065, 5.00028, 5.000989, 5.002667, 5.005479, 5.00688, 5.007271, 
    5.00688, 5.005479, 5.002667, 5.000989, 5.00028, 5.000065, 5.000013, 
    5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // height(1,38, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000009, 
    5.000041, 5.000161, 5.000472, 5.00103, 5.001293, 5.001361, 5.001293, 
    5.00103, 5.000472, 5.000161, 5.000041, 5.000009, 5.000001, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // height(1,39, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000005, 
    5.000022, 5.000071, 5.000165, 5.000208, 5.000218, 5.000208, 5.000165, 
    5.000071, 5.000022, 5.000005, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5,
  // height(1,40, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 
    5.00001, 5.000023, 5.000029, 5.00003, 5.000029, 5.000023, 5.00001, 
    5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // height(1,41, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5.000001, 5.000003, 5.000003, 5.000003, 5.000003, 5.000003, 5.000001, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // height(1,42, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // height(1,43, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // height(1,44, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // height(1,45, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // height(1,46, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // height(1,47, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // height(1,48, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // height(1,49, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // height(2,0, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // height(2,1, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // height(2,2, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // height(2,3, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5.000001, 5.000001, 5.000001, 5.000001, 5.000001, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // height(2,4, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 
    5.000003, 5.000006, 5.000008, 5.000009, 5.000008, 5.000006, 5.000003, 
    5.000001, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // height(2,5, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 
    5.000003, 5.000009, 5.000018, 5.00003, 5.000037, 5.000041, 5.000037, 
    5.00003, 5.000018, 5.000009, 5.000003, 5.000001, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // height(2,6, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000008, 
    5.00002, 5.000044, 5.000084, 5.000135, 5.000167, 5.000179, 5.000167, 
    5.000135, 5.000084, 5.000044, 5.00002, 5.000008, 5.000002, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // height(2,7, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000004, 5.000013, 
    5.000036, 5.000087, 5.000192, 5.000359, 5.000562, 5.000698, 5.000745, 
    5.000698, 5.000562, 5.000359, 5.000192, 5.000087, 5.000036, 5.000013, 
    5.000004, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // height(2,8, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000005, 
    5.000019, 5.000055, 5.000149, 5.000361, 5.000768, 5.001396, 5.002146, 
    5.002654, 5.002829, 5.002654, 5.002146, 5.001396, 5.000768, 5.000361, 
    5.000149, 5.000055, 5.000019, 5.000005, 5.000001, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5,
  // height(2,9, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000007, 5.000025, 
    5.00008, 5.00023, 5.000596, 5.001375, 5.002819, 5.004971, 5.00749, 
    5.009201, 5.009799, 5.009201, 5.00749, 5.004971, 5.002819, 5.001375, 
    5.000596, 5.00023, 5.00008, 5.000025, 5.000007, 5.000001, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5,
  // height(2,10, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000008, 5.000031, 
    5.000104, 5.000319, 5.000876, 5.002162, 5.004771, 5.009418, 5.016093, 
    5.023739, 5.028931, 5.030761, 5.028931, 5.023739, 5.016093, 5.009418, 
    5.004771, 5.002162, 5.000876, 5.000319, 5.000104, 5.000031, 5.000008, 
    5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // height(2,11, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.00001, 5.000034, 
    5.000126, 5.000408, 5.001172, 5.003046, 5.007127, 5.014987, 5.028435, 
    5.046975, 5.067611, 5.08152, 5.086449, 5.08152, 5.067611, 5.046975, 
    5.028435, 5.014987, 5.007127, 5.003045, 5.001171, 5.000405, 5.000127, 
    5.000036, 5.00001, 5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // height(2,12, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000009, 5.000036, 5.000136, 
    5.000466, 5.001442, 5.003905, 5.00958, 5.021203, 5.042273, 5.076715, 
    5.121716, 5.169673, 5.201324, 5.212531, 5.201324, 5.169673, 5.121716, 
    5.076715, 5.042273, 5.021201, 5.009576, 5.003897, 5.00143, 5.000474, 
    5.000143, 5.000039, 5.00001, 5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // height(2,13, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000008, 5.000033, 5.000133, 
    5.000481, 5.00157, 5.004634, 5.011772, 5.027131, 5.05641, 5.105655, 
    5.181499, 5.273223, 5.364344, 5.422204, 5.4425, 5.422204, 5.364344, 
    5.273223, 5.181498, 5.105653, 5.056403, 5.02711, 5.011728, 5.004572, 
    5.001609, 5.000513, 5.000149, 5.000039, 5.00001, 5.000002, 5, 5, 5, 5, 5, 
    5, 5, 5, 5,
  // height(2,14, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000007, 5.000029, 5.000118, 5.000446, 
    5.001536, 5.004781, 5.013485, 5.031936, 5.068588, 5.132482, 5.229629, 
    5.367397, 5.516597, 5.650199, 5.73082, 5.75868, 5.73082, 5.650199, 
    5.516597, 5.367393, 5.229616, 5.132443, 5.068489, 5.031737, 5.013205, 
    5.004946, 5.001672, 5.000513, 5.000143, 5.000036, 5.000008, 5.000001, 5, 
    5, 5, 5, 5, 5, 5, 5,
  // height(2,15, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000004, 5.000021, 5.000093, 5.000368, 
    5.001338, 5.004398, 5.013077, 5.035445, 5.07743, 5.152986, 5.270136, 
    5.425341, 5.623005, 5.808567, 5.954159, 6.038265, 6.066943, 6.038265, 
    5.954158, 5.808562, 5.622989, 5.425284, 5.269968, 5.152572, 5.076609, 
    5.034278, 5.01373, 5.004946, 5.001609, 5.000474, 5.000127, 5.000031, 
    5.000007, 5.000001, 5, 5, 5, 5, 5, 5, 5,
  // height(2,16, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000014, 5.000063, 5.000268, 5.001024, 
    5.003561, 5.011195, 5.031907, 5.083897, 5.166404, 5.297246, 5.471339, 
    5.663941, 5.881144, 6.054009, 6.170801, 6.238191, 6.261086, 6.23819, 
    6.170798, 6.053992, 5.881079, 5.663725, 5.470706, 5.295689, 5.163324, 
    5.079466, 5.034278, 5.013205, 5.004572, 5.00143, 5.000405, 5.000104, 
    5.000025, 5.000005, 5, 5, 5, 5, 5, 5, 5,
  // height(2,17, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000008, 5.000038, 5.000165, 5.00067, 
    5.002472, 5.008275, 5.024992, 5.068762, 5.178341, 5.314689, 5.498798, 
    5.701071, 5.878989, 6.057094, 6.174425, 6.241654, 6.28508, 6.300066, 
    6.285078, 6.24164, 6.174369, 6.056881, 5.878283, 5.699006, 5.493689, 
    5.304491, 5.163324, 5.076609, 5.031737, 5.011728, 5.003897, 5.001171, 
    5.000319, 5.00008, 5.000019, 5.000004, 5, 5, 5, 5, 5, 5,
  // height(2,18, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5.000003, 5.000017, 5.000082, 5.000356, 5.001401, 
    5.005028, 5.016359, 5.047846, 5.129076, 5.339933, 5.523062, 5.725195, 
    5.900149, 6.010222, 6.107472, 6.153584, 6.174073, 6.196599, 6.204854, 
    6.196589, 6.174033, 6.153419, 6.106858, 6.008182, 5.894237, 5.710595, 
    5.493689, 5.295689, 5.152572, 5.068489, 5.02711, 5.009576, 5.003045, 
    5.000876, 5.00023, 5.000055, 5.000013, 5.000002, 5, 5, 5, 5, 5,
  // height(2,19, 0-49)
    5, 5, 5, 5, 5, 5, 5.000001, 5.000007, 5.000029, 5.000135, 5.000575, 
    5.002245, 5.008015, 5.025926, 5.074886, 5.206708, 5.580922, 5.772137, 
    5.930871, 6.024444, 6.039964, 6.04226, 6.020387, 6.004436, 6.009708, 
    6.012484, 6.009684, 6.004327, 6.019951, 6.040654, 6.034697, 6.009424, 
    5.894236, 5.699005, 5.470706, 5.269968, 5.132443, 5.056403, 5.021201, 
    5.007127, 5.002162, 5.000596, 5.000149, 5.000036, 5.000008, 5.000001, 5, 
    5, 5, 5,
  // height(2,20, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5.000001, 5.00001, 5.000042, 5.000171, 5.000613, 
    5.001966, 5.005518, 5.013143, 0, 6.070654, 6.10031, 6.109229, 6.073961, 
    5.989838, 5.897338, 5.812802, 5.764136, 5.750331, 5.746961, 5.750273, 
    5.763871, 5.811723, 5.893331, 5.976495, 6.034697, 6.008182, 5.878282, 
    5.663725, 5.425284, 5.229616, 5.105653, 5.042273, 5.014987, 5.004771, 
    5.001375, 5.000361, 5.000087, 5.00002, 5.000003, 5, 5, 5, 5,
  // height(2,21, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5.000003, 5.000014, 5.000054, 5.000195, 5.00063, 
    5.001772, 5.004181, 0, 6.513035, 6.426273, 6.282675, 6.110457, 5.917133, 
    5.702082, 5.514227, 5.387189, 5.318944, 5.296926, 5.318848, 5.386738, 
    5.51234, 5.694969, 5.893331, 6.040654, 6.106857, 6.056882, 5.88108, 
    5.622988, 5.367393, 5.181498, 5.076715, 5.028435, 5.009418, 5.002819, 
    5.000768, 5.000192, 5.000044, 5.000009, 5.000001, 5, 5, 5,
  // height(2,22, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000004, 5.000016, 5.000055, 5.000182, 
    5.000515, 5.001205, 0, 6.890601, 6.696692, 6.413081, 6.125101, 5.847679, 
    5.523096, 5.231614, 5.02129, 4.898302, 4.858558, 4.898164, 5.020628, 
    5.228783, 5.512339, 5.811723, 6.019951, 6.153419, 6.174369, 6.053992, 
    5.808561, 5.516597, 5.273223, 5.121716, 5.046975, 5.016093, 5.004971, 
    5.001396, 5.000359, 5.000084, 5.000018, 5.000003, 5, 5, 5,
  // height(2,23, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000004, 5.000016, 5.000049, 5.000141, 
    5.000327, 0, 7.175317, 6.901651, 6.513165, 6.143483, 5.81144, 5.400992, 
    5.024344, 4.753988, 4.602839, 4.55656, 4.602668, 4.753143, 5.020628, 
    5.386737, 5.76387, 6.004326, 6.174033, 6.241639, 6.170797, 5.954158, 
    5.650199, 5.364344, 5.169673, 5.067611, 5.023739, 5.00749, 5.002146, 
    5.000562, 5.000135, 5.00003, 5.000006, 5.000001, 5, 5,
  // height(2,24, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000006, 5.00002, 5.000057, 5.000128, 
    0, 7.33971, 7.028852, 6.586917, 6.171556, 5.805634, 5.335411, 4.902411, 
    4.603594, 4.448595, 4.40392, 4.448415, 4.602663, 4.89816, 5.318843, 
    5.750269, 6.009683, 6.196589, 6.285078, 6.23819, 6.038265, 5.73082, 
    5.422204, 5.201324, 5.08152, 5.028931, 5.009201, 5.002654, 5.000698, 
    5.000167, 5.000037, 5.000008, 5.000001, 5, 5,
  // height(2,25, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000003, 5.000013, 5.000041, 5.000108, 
    5.000237, 0, 7.394997, 7.072412, 6.612961, 6.182293, 5.805012, 5.31426, 
    4.862948, 4.55748, 4.40407, 4.360934, 4.403889, 4.556526, 4.858529, 
    5.296904, 5.746947, 6.012478, 6.204852, 6.300065, 6.261086, 6.066943, 
    5.75868, 5.4425, 5.212531, 5.086449, 5.030761, 5.009799, 5.002829, 
    5.000745, 5.000179, 5.000041, 5.000009, 5.000001, 5, 5,
  // height(2,26, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000003, 5.000014, 5.000048, 5.000146, 
    5.00039, 5.000851, 0, 7.33743, 7.027562, 6.586339, 6.171353, 5.805575, 
    5.335398, 4.902407, 4.603593, 4.448595, 4.403919, 4.448415, 4.602663, 
    4.898159, 5.318843, 5.750269, 6.009683, 6.196589, 6.285078, 6.23819, 
    6.038265, 5.73082, 5.422204, 5.201324, 5.08152, 5.028931, 5.009201, 
    5.002654, 5.000698, 5.000167, 5.000037, 5.000008, 5.000001, 5, 5,
  // height(2,27, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5.000003, 5.000013, 5.000049, 5.000171, 5.000519, 
    5.001362, 5.002976, 0, 7.16783, 6.897426, 6.511255, 6.142797, 5.811236, 
    5.40094, 5.024333, 4.753986, 4.602839, 4.55656, 4.602669, 4.753144, 
    5.020627, 5.386737, 5.76387, 6.004327, 6.174033, 6.24164, 6.170797, 
    5.954158, 5.650199, 5.364344, 5.169673, 5.067611, 5.023739, 5.00749, 
    5.002146, 5.000562, 5.000135, 5.00003, 5.000006, 5.000001, 5, 5,
  // height(2,28, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5.000002, 5.00001, 5.000044, 5.000165, 5.000557, 
    5.001666, 5.004333, 5.009483, 0, 6.869401, 6.684888, 6.407736, 6.123141, 
    5.847076, 5.522937, 5.231577, 5.021283, 4.898301, 4.858558, 4.898164, 
    5.020629, 5.228784, 5.51234, 5.811723, 6.019951, 6.153419, 6.174369, 
    6.053992, 5.808561, 5.516597, 5.273223, 5.121716, 5.046975, 5.016093, 
    5.004971, 5.001396, 5.000359, 5.000084, 5.000018, 5.000003, 5, 5, 5,
  // height(2,29, 0-49)
    5, 5, 5, 5, 5, 5, 5.000001, 5.000007, 5.000031, 5.00013, 5.000485, 
    5.001624, 5.004813, 5.012438, 5.027185, 0, 6.458423, 6.39655, 6.269349, 
    6.105521, 5.915573, 5.701647, 5.514119, 5.387164, 5.318938, 5.296925, 
    5.318848, 5.386738, 5.51234, 5.694969, 5.893331, 6.040654, 6.106858, 
    6.056882, 5.88108, 5.622988, 5.367393, 5.181498, 5.076715, 5.028435, 
    5.009418, 5.002819, 5.000768, 5.000192, 5.000044, 5.000009, 5.000001, 5, 
    5, 5,
  // height(2,30, 0-49)
    5, 5, 5, 5, 5, 5, 5.000004, 5.000019, 5.000091, 5.000392, 5.001544, 
    5.005568, 5.018255, 5.053765, 5.13902, 5.339774, 5.824156, 5.992731, 
    6.068674, 6.060568, 5.985876, 5.89627, 5.812539, 5.764076, 5.750317, 
    5.746958, 5.750272, 5.763871, 5.811723, 5.893331, 5.976495, 6.034697, 
    6.008182, 5.878283, 5.663725, 5.425284, 5.229616, 5.105653, 5.042273, 
    5.014987, 5.004771, 5.001375, 5.000361, 5.000087, 5.00002, 5.000003, 5, 
    5, 5, 5,
  // height(2,31, 0-49)
    5, 5, 5, 5, 5, 5, 5.000002, 5.000012, 5.000059, 5.000257, 5.001028, 
    5.003737, 5.01235, 5.036781, 5.097425, 5.235366, 5.544514, 5.750298, 
    5.92068, 6.020491, 6.03864, 6.041875, 6.020286, 6.00441, 6.009703, 
    6.012483, 6.009684, 6.004327, 6.019951, 6.040655, 6.034697, 6.009424, 
    5.894237, 5.699006, 5.470706, 5.269968, 5.132443, 5.056403, 5.021201, 
    5.007127, 5.002162, 5.000596, 5.000149, 5.000036, 5.000008, 5.000001, 5, 
    5, 5, 5,
  // height(2,32, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5.000005, 5.000028, 5.000126, 5.000518, 5.00194, 
    5.006609, 5.020349, 5.056161, 5.140028, 5.324083, 5.513662, 5.720868, 
    5.898491, 6.009674, 6.107315, 6.153543, 6.174064, 6.196596, 6.204853, 
    6.196589, 6.174033, 6.153419, 6.106858, 6.008182, 5.894237, 5.710595, 
    5.493689, 5.295689, 5.152572, 5.068489, 5.02711, 5.009576, 5.003045, 
    5.000876, 5.00023, 5.000055, 5.000013, 5.000002, 5, 5, 5, 5, 5,
  // height(2,33, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000011, 5.000051, 5.000216, 5.000844, 
    5.002991, 5.009605, 5.02779, 5.072512, 5.172647, 5.311225, 5.497193, 
    5.700458, 5.878788, 6.057036, 6.17441, 6.241651, 6.28508, 6.300066, 
    6.285078, 6.241639, 6.174369, 6.056882, 5.878283, 5.699006, 5.493689, 
    5.304491, 5.163324, 5.076609, 5.031737, 5.011728, 5.003897, 5.001171, 
    5.000319, 5.00008, 5.000019, 5.000004, 5, 5, 5, 5, 5, 5,
  // height(2,34, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5.000003, 5.000018, 5.000078, 5.000318, 5.001177, 
    5.003963, 5.012051, 5.033063, 5.082146, 5.165304, 5.29673, 5.471141, 
    5.663877, 5.881125, 6.054005, 6.170801, 6.238191, 6.261086, 6.238191, 
    6.170798, 6.053992, 5.88108, 5.663725, 5.470706, 5.295689, 5.163324, 
    5.079466, 5.034278, 5.013205, 5.004572, 5.00143, 5.000405, 5.000104, 
    5.000025, 5.000005, 5, 5, 5, 5, 5, 5, 5,
  // height(2,35, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000006, 5.000025, 5.000106, 5.000411, 
    5.001449, 5.004638, 5.0134, 5.034968, 5.077124, 5.152843, 5.270081, 
    5.425323, 5.623, 5.808566, 5.954159, 6.038265, 6.066944, 6.038265, 
    5.954159, 5.808562, 5.622989, 5.425284, 5.269968, 5.152572, 5.076609, 
    5.034278, 5.01373, 5.004946, 5.001609, 5.000474, 5.000127, 5.000031, 
    5.000007, 5.000001, 5, 5, 5, 5, 5, 5, 5,
  // height(2,36, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000007, 5.000031, 5.000127, 
    5.000473, 5.001596, 5.004863, 5.013367, 5.031859, 5.068552, 5.132469, 
    5.229624, 5.367395, 5.516597, 5.650199, 5.73082, 5.75868, 5.73082, 
    5.650199, 5.516597, 5.367393, 5.229616, 5.132443, 5.068489, 5.031737, 
    5.013205, 5.004946, 5.001672, 5.000513, 5.000143, 5.000036, 5.000008, 
    5.000001, 5, 5, 5, 5, 5, 5, 5, 5,
  // height(2,37, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000009, 5.000036, 5.000139, 
    5.000494, 5.001589, 5.004607, 5.011755, 5.027123, 5.056408, 5.105654, 
    5.181498, 5.273223, 5.364344, 5.422204, 5.4425, 5.422204, 5.364344, 
    5.273223, 5.181498, 5.105653, 5.056403, 5.02711, 5.011728, 5.004572, 
    5.001609, 5.000513, 5.000149, 5.000039, 5.00001, 5.000002, 5, 5, 5, 5, 5, 
    5, 5, 5, 5,
  // height(2,38, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.00001, 5.000037, 5.000138, 
    5.00047, 5.001437, 5.003901, 5.009578, 5.021202, 5.042273, 5.076715, 
    5.121716, 5.169673, 5.201324, 5.212531, 5.201324, 5.169673, 5.121716, 
    5.076715, 5.042273, 5.021201, 5.009576, 5.003897, 5.00143, 5.000474, 
    5.000143, 5.000039, 5.00001, 5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // height(2,39, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.00001, 5.000034, 
    5.000126, 5.000407, 5.001172, 5.003045, 5.007127, 5.014987, 5.028435, 
    5.046975, 5.067611, 5.08152, 5.086449, 5.08152, 5.067611, 5.046975, 
    5.028435, 5.014987, 5.007127, 5.003045, 5.001171, 5.000405, 5.000127, 
    5.000036, 5.00001, 5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // height(2,40, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000008, 5.000031, 
    5.000104, 5.000319, 5.000876, 5.002162, 5.004771, 5.009418, 5.016093, 
    5.023739, 5.028931, 5.030761, 5.028931, 5.023739, 5.016093, 5.009418, 
    5.004771, 5.002162, 5.000876, 5.000319, 5.000104, 5.000031, 5.000008, 
    5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // height(2,41, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000007, 5.000025, 
    5.00008, 5.00023, 5.000596, 5.001375, 5.002819, 5.004971, 5.00749, 
    5.009201, 5.009799, 5.009201, 5.00749, 5.004971, 5.002819, 5.001375, 
    5.000596, 5.00023, 5.00008, 5.000025, 5.000007, 5.000001, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5,
  // height(2,42, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000005, 
    5.000019, 5.000055, 5.000149, 5.000361, 5.000768, 5.001396, 5.002146, 
    5.002654, 5.002829, 5.002654, 5.002146, 5.001396, 5.000768, 5.000361, 
    5.000149, 5.000055, 5.000019, 5.000005, 5.000001, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5,
  // height(2,43, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000004, 5.000013, 
    5.000036, 5.000087, 5.000192, 5.000359, 5.000562, 5.000698, 5.000745, 
    5.000698, 5.000562, 5.000359, 5.000192, 5.000087, 5.000036, 5.000013, 
    5.000004, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // height(2,44, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000008, 
    5.00002, 5.000044, 5.000084, 5.000135, 5.000167, 5.000179, 5.000167, 
    5.000135, 5.000084, 5.000044, 5.00002, 5.000008, 5.000002, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // height(2,45, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 
    5.000003, 5.000009, 5.000018, 5.00003, 5.000037, 5.000041, 5.000037, 
    5.00003, 5.000018, 5.000009, 5.000003, 5.000001, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // height(2,46, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 
    5.000003, 5.000006, 5.000008, 5.000009, 5.000008, 5.000006, 5.000003, 
    5.000001, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // height(2,47, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5.000001, 5.000001, 5.000001, 5.000001, 5.000001, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // height(2,48, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // height(2,49, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // height(3,0, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 
    5.000003, 5.000006, 5.00001, 5.000014, 5.000018, 5.000019, 5.000018, 
    5.000014, 5.00001, 5.000006, 5.000003, 5.000001, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // height(3,1, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000007, 
    5.000014, 5.000024, 5.000038, 5.000054, 5.000065, 5.000069, 5.000065, 
    5.000054, 5.000038, 5.000024, 5.000014, 5.000007, 5.000002, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // height(3,2, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000005, 
    5.000013, 5.000025, 5.000051, 5.000089, 5.000139, 5.000192, 5.00023, 
    5.000245, 5.00023, 5.000192, 5.000139, 5.000089, 5.000051, 5.000025, 
    5.000013, 5.000005, 5.000001, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // height(3,3, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000003, 5.000008, 5.00002, 
    5.000045, 5.000092, 5.000175, 5.000303, 5.000471, 5.000645, 5.000771, 
    5.000815, 5.000771, 5.000645, 5.000471, 5.000303, 5.000175, 5.000092, 
    5.000045, 5.00002, 5.000008, 5.000003, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5,
  // height(3,4, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000004, 5.000012, 5.00003, 
    5.00007, 5.000153, 5.000309, 5.000576, 5.000975, 5.001488, 5.002019, 
    5.0024, 5.002537, 5.0024, 5.002019, 5.001488, 5.000975, 5.000576, 
    5.000309, 5.000153, 5.00007, 5.00003, 5.000012, 5.000004, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5,
  // height(3,5, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000005, 5.000016, 
    5.000041, 5.000101, 5.000232, 5.000495, 5.000975, 5.001767, 5.002935, 
    5.004404, 5.005916, 5.006993, 5.007383, 5.006993, 5.005916, 5.004404, 
    5.002935, 5.001767, 5.000974, 5.000495, 5.000232, 5.000101, 5.000041, 
    5.000016, 5.000005, 5.000001, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // height(3,6, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000007, 5.00002, 5.000052, 
    5.000135, 5.000328, 5.000727, 5.001502, 5.002871, 5.005065, 5.008235, 
    5.012152, 5.016148, 5.018981, 5.020005, 5.018981, 5.016148, 5.012152, 
    5.008235, 5.005065, 5.00287, 5.001501, 5.000726, 5.000327, 5.000136, 
    5.000052, 5.00002, 5.000007, 5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // height(3,7, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000008, 5.000022, 5.000062, 
    5.000168, 5.000426, 5.000994, 5.002136, 5.004256, 5.007876, 5.013505, 
    5.021459, 5.0311, 5.040833, 5.047673, 5.050141, 5.047673, 5.040833, 
    5.0311, 5.021459, 5.013503, 5.007874, 5.004254, 5.00213, 5.000989, 
    5.000427, 5.000171, 5.000064, 5.000023, 5.000008, 5.000002, 5, 5, 5, 5, 
    5, 5, 5, 5, 5,
  // height(3,8, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000008, 5.000023, 5.000071, 
    5.000197, 5.000516, 5.001256, 5.002826, 5.005837, 5.011214, 5.020035, 
    5.033278, 5.051542, 5.073155, 5.094623, 5.109491, 5.114835, 5.109491, 
    5.094623, 5.073154, 5.05154, 5.033274, 5.020027, 5.011199, 5.005819, 
    5.002808, 5.001259, 5.000525, 5.000204, 5.000074, 5.000025, 5.000008, 
    5.000002, 5, 5, 5, 5, 5, 5, 5, 5,
  // height(3,9, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000008, 5.000024, 5.000072, 5.000215, 
    5.000583, 5.001472, 5.003447, 5.007477, 5.01482, 5.027332, 5.046957, 
    5.07516, 5.112832, 5.155911, 5.197577, 5.225729, 5.235758, 5.225728, 
    5.197576, 5.155908, 5.112823, 5.075142, 5.046923, 5.027278, 5.014745, 
    5.00741, 5.003462, 5.001504, 5.000608, 5.000228, 5.00008, 5.000026, 
    5.000009, 5.000002, 5, 5, 5, 5, 5, 5, 5,
  // height(3,10, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000007, 5.000022, 5.000071, 5.000216, 
    5.00061, 5.001602, 5.003899, 5.008797, 5.018371, 5.034782, 5.061243, 
    5.100461, 5.15364, 5.221577, 5.295402, 5.36382, 5.408352, 5.423996, 
    5.408351, 5.363815, 5.29539, 5.221547, 5.153577, 5.100338, 5.061041, 
    5.034512, 5.018124, 5.008841, 5.004006, 5.001688, 5.000662, 5.000242, 
    5.000082, 5.000026, 5.000008, 5.000002, 5, 5, 5, 5, 5, 5,
  // height(3,11, 0-49)
    5, 5, 5, 5, 5, 5, 5.000001, 5.000006, 5.000021, 5.000064, 5.000203, 
    5.000594, 5.001617, 5.004089, 5.009582, 5.020787, 5.04175, 5.075024, 
    5.125049, 5.193873, 5.280046, 5.383638, 5.488432, 5.579867, 5.636599, 
    5.656176, 5.636593, 5.57985, 5.488389, 5.383534, 5.279824, 5.193449, 
    5.124352, 5.074101, 5.040899, 5.020916, 5.009921, 5.004369, 5.001788, 
    5.000681, 5.000242, 5.00008, 5.000025, 5.000008, 5.000002, 5, 5, 5, 5, 5,
  // height(3,12, 0-49)
    5, 5, 5, 5, 5, 5, 5.000005, 5.000017, 5.000055, 5.000177, 5.000535, 
    5.001513, 5.003968, 5.009657, 5.021753, 5.045288, 5.087358, 5.14761, 
    5.230261, 5.333305, 5.449304, 5.57871, 5.698251, 5.795069, 5.852182, 
    5.871558, 5.852166, 5.795019, 5.698119, 5.578391, 5.448622, 5.331985, 
    5.228084, 5.144711, 5.084641, 5.045663, 5.022761, 5.010503, 5.004496, 
    5.001788, 5.000662, 5.000228, 5.000074, 5.000023, 5.000007, 5.000001, 5, 
    5, 5, 5,
  // height(3,13, 0-49)
    5, 5, 5, 5, 5, 5.000002, 5.000013, 5.000043, 5.000142, 5.000446, 
    5.001304, 5.003549, 5.008974, 5.021013, 5.045398, 5.090425, 5.167326, 
    5.262846, 5.378967, 5.506453, 5.631666, 5.760675, 5.867614, 5.947062, 
    5.992007, 6.007091, 5.991964, 5.946927, 5.867256, 5.75981, 5.629799, 
    5.502812, 5.372893, 5.25464, 5.159427, 5.091476, 5.048205, 5.023404, 
    5.010503, 5.004369, 5.001688, 5.000608, 5.000204, 5.000064, 5.00002, 
    5.000005, 5, 5, 5, 5,
  // height(3,14, 0-49)
    5, 5, 5, 5, 5.000001, 5.000009, 5.000031, 5.000105, 5.00034, 5.001029, 
    5.002908, 5.007648, 5.018635, 5.041913, 5.086556, 5.164249, 5.291772, 
    5.421392, 5.55587, 5.681244, 5.783919, 5.882294, 5.952684, 5.99908, 
    6.024866, 6.03354, 6.024758, 5.998743, 5.951796, 5.880162, 5.77933, 
    5.672307, 5.540854, 5.400769, 5.271254, 5.167127, 5.093842, 5.048205, 
    5.022761, 5.009921, 5.004006, 5.001504, 5.000525, 5.000171, 5.000052, 
    5.000016, 5.000004, 5, 5, 5,
  // height(3,15, 0-49)
    5, 5, 5, 5, 5.000005, 5.00002, 5.000069, 5.000233, 5.000735, 5.002163, 
    5.005921, 5.015044, 5.035314, 5.076136, 5.14962, 5.26931, 5.461556, 
    5.608839, 5.731626, 5.821412, 5.873544, 5.920516, 5.942305, 5.950413, 
    5.955587, 5.957473, 5.955333, 5.949632, 5.940266, 5.915689, 5.863268, 
    5.801664, 5.698636, 5.56323, 5.414839, 5.276899, 5.167127, 5.091476, 
    5.045663, 5.020916, 5.00884, 5.003462, 5.001259, 5.000427, 5.000136, 
    5.000041, 5.000012, 5.000003, 5, 5,
  // height(3,16, 0-49)
    5, 5, 5, 5.000002, 5.000011, 5.000041, 5.000143, 5.000468, 5.001436, 
    5.004103, 5.010897, 5.026792, 5.060598, 5.124972, 5.232549, 5.396155, 
    5.662586, 5.799902, 5.878317, 5.906157, 5.892824, 5.879972, 5.850737, 
    5.821409, 5.806584, 5.801819, 5.806024, 5.819709, 5.846377, 5.869823, 
    5.871604, 5.866385, 5.813318, 5.711125, 5.5706, 5.414839, 5.271254, 
    5.159427, 5.084641, 5.040899, 5.018124, 5.00741, 5.002808, 5.000989, 
    5.000327, 5.000101, 5.00003, 5.000008, 5.000001, 5,
  // height(3,17, 0-49)
    5, 5, 5.000001, 5.000005, 5.000021, 5.000075, 5.000259, 5.000828, 
    5.002479, 5.006911, 5.017881, 5.042683, 5.093165, 5.18362, 5.322259, 
    5.521502, 5.866402, 5.969814, 5.983183, 5.936786, 5.854723, 5.780489, 
    5.701207, 5.636169, 5.601222, 5.58957, 5.600065, 5.632699, 5.692458, 
    5.76054, 5.814003, 5.863031, 5.867137, 5.816883, 5.711125, 5.56323, 
    5.400769, 5.25464, 5.144711, 5.0741, 5.034512, 5.014745, 5.005819, 
    5.00213, 5.000726, 5.000232, 5.00007, 5.00002, 5.000005, 5,
  // height(3,18, 0-49)
    5, 5, 5.000002, 5.000009, 5.000031, 5.000117, 5.000395, 5.001246, 
    5.003667, 5.010052, 5.025521, 5.059556, 5.126149, 5.238306, 5.394081, 
    5.615667, 6.035935, 6.101533, 6.04922, 5.929343, 5.78085, 5.644381, 
    5.515065, 5.414158, 5.357251, 5.337825, 5.354997, 5.407474, 5.498516, 
    5.607554, 5.707836, 5.802571, 5.86004, 5.867137, 5.813318, 5.698636, 
    5.540854, 5.372893, 5.228083, 5.124352, 5.061041, 5.027278, 5.011199, 
    5.004254, 5.001501, 5.000495, 5.000153, 5.000045, 5.000013, 5.000002,
  // height(3,19, 0-49)
    5, 5, 5.000002, 5.000011, 5.000038, 5.00014, 5.000471, 5.001475, 
    5.004326, 5.011827, 5.029943, 5.069492, 5.145236, 5.266404, 5.417098, 
    5.657688, 6.133231, 6.183744, 6.085767, 5.90326, 5.691944, 5.490312, 
    5.308599, 5.169163, 5.086947, 5.058302, 5.082806, 5.156998, 5.279012, 
    5.426208, 5.569045, 5.70021, 5.80257, 5.863031, 5.866385, 5.801664, 
    5.672307, 5.502812, 5.331985, 5.193449, 5.100338, 5.046923, 5.020027, 
    5.007874, 5.00287, 5.000974, 5.000309, 5.000092, 5.000025, 5.000007,
  // height(3,20, 0-49)
    5, 5, 5.000001, 5.000006, 5.000022, 5.000076, 5.000246, 5.000745, 
    5.002099, 5.005454, 5.012992, 5.028082, 5.054316, 5.092286, 5.134862, 0, 
    6.537839, 6.444597, 6.224334, 5.931908, 5.627497, 5.341224, 5.09673, 
    4.91181, 4.799217, 4.759322, 4.791854, 4.890079, 5.043821, 5.226887, 
    5.408791, 5.569041, 5.707834, 5.814003, 5.871604, 5.863268, 5.779329, 
    5.629799, 5.448622, 5.279824, 5.153577, 5.075142, 5.033274, 5.013503, 
    5.005065, 5.001767, 5.000576, 5.000175, 5.000051, 5.000014,
  // height(3,21, 0-49)
    5, 5, 5, 5.000002, 5.000011, 5.000037, 5.000119, 5.000364, 5.001029, 
    5.002694, 5.006472, 5.01416, 5.027897, 5.048741, 5.073972, 0, 6.715348, 
    6.582877, 6.306049, 5.934135, 5.539999, 5.157746, 4.834559, 4.587932, 
    4.433352, 4.378251, 4.422956, 4.55676, 4.757838, 4.992012, 5.226871, 
    5.426194, 5.607547, 5.760535, 5.869822, 5.915688, 5.880161, 5.75981, 
    5.578391, 5.383534, 5.221547, 5.112823, 5.05154, 5.021459, 5.008235, 
    5.002935, 5.000975, 5.000303, 5.000089, 5.000024,
  // height(3,22, 0-49)
    5, 5, 5, 5, 5.000004, 5.000016, 5.000052, 5.00016, 5.000462, 5.001224, 
    5.002986, 5.006641, 5.013321, 5.023751, 5.036767, 0, 6.819324, 6.665093, 
    6.350619, 5.917248, 5.445622, 4.973551, 4.571023, 4.255342, 4.050066, 
    3.976002, 4.036703, 4.214768, 4.470624, 4.757758, 5.043741, 5.278961, 
    5.498487, 5.692443, 5.846371, 5.940264, 5.951795, 5.867255, 5.69812, 
    5.488389, 5.29539, 5.155908, 5.073154, 5.0311, 5.012152, 5.004404, 
    5.001488, 5.000471, 5.000139, 5.000038,
  // height(3,23, 0-49)
    5, 5, 5, 5, 5.000001, 5.000007, 5.000022, 5.00007, 5.000204, 5.000552, 
    5.001373, 5.003109, 5.006342, 5.011469, 5.017878, 0, 6.881858, 6.715767, 
    6.377157, 5.89924, 5.365091, 4.814788, 4.335211, 3.944315, 3.680533, 
    3.584269, 3.664799, 3.895799, 4.214448, 4.556406, 4.88979, 5.156824, 
    5.407378, 5.63265, 5.819686, 5.949622, 5.99874, 5.946925, 5.795018, 
    5.57985, 5.363815, 5.197576, 5.094623, 5.040833, 5.016148, 5.005916, 
    5.002019, 5.000645, 5.000192, 5.000054,
  // height(3,24, 0-49)
    5, 5, 5, 5, 5, 5.000004, 5.000014, 5.000044, 5.000131, 5.000354, 
    5.000885, 5.002009, 5.004103, 5.00741, 5.011444, 0, 6.913795, 6.743283, 
    6.393038, 5.88919, 5.313772, 4.708361, 4.169513, 3.717096, 3.405324, 
    3.291309, 3.388295, 3.663615, 4.035308, 4.421719, 4.790909, 5.082253, 
    5.354696, 5.599913, 5.805953, 5.955301, 6.024744, 5.991959, 5.852164, 
    5.636593, 5.40835, 5.225728, 5.109491, 5.047673, 5.018981, 5.006993, 
    5.0024, 5.000771, 5.00023, 5.000065,
  // height(3,25, 0-49)
    5, 5, 5, 5, 5.000001, 5.000007, 5.000023, 5.000068, 5.000196, 5.000519, 
    5.001256, 5.00277, 5.005505, 5.009689, 5.014659, 0, 6.917509, 6.746934, 
    6.394336, 5.883124, 5.294426, 4.670211, 4.109842, 3.634244, 3.304592, 
    3.184185, 3.287201, 3.579186, 3.97121, 4.374317, 4.756428, 5.056643, 
    5.336924, 5.589113, 5.801601, 5.957374, 6.033497, 6.007074, 5.871552, 
    5.656174, 5.423996, 5.235758, 5.114835, 5.050141, 5.020005, 5.007383, 
    5.002537, 5.000815, 5.000245, 5.000069,
  // height(3,26, 0-49)
    5, 5, 5, 5, 5.000005, 5.000018, 5.000054, 5.000162, 5.000451, 5.001157, 
    5.00272, 5.005827, 5.011258, 5.019319, 5.028754, 0, 6.889607, 6.723534, 
    6.378369, 5.879577, 5.308405, 4.705863, 4.168527, 3.716762, 3.405225, 
    3.291283, 3.388287, 3.663613, 4.035307, 4.421719, 4.790908, 5.082252, 
    5.354695, 5.599913, 5.805953, 5.955301, 6.024744, 5.991959, 5.852164, 
    5.636593, 5.40835, 5.225728, 5.109491, 5.047673, 5.018981, 5.006993, 
    5.0024, 5.000771, 5.00023, 5.000065,
  // height(3,27, 0-49)
    5, 5, 5, 5.000003, 5.000013, 5.000042, 5.000131, 5.000385, 5.001048, 
    5.002628, 5.006048, 5.012661, 5.02387, 5.039977, 5.058367, 0, 6.826754, 
    6.670672, 6.343395, 5.876875, 5.352436, 4.808751, 4.332749, 3.943442, 
    3.680258, 3.58419, 3.664778, 3.895793, 4.214446, 4.556406, 4.889789, 
    5.156823, 5.407378, 5.63265, 5.819686, 5.949621, 5.99874, 5.946925, 
    5.795018, 5.57985, 5.363815, 5.197576, 5.094623, 5.040833, 5.016148, 
    5.005916, 5.002019, 5.000645, 5.000192, 5.000054,
  // height(3,28, 0-49)
    5, 5, 5.000001, 5.000009, 5.000028, 5.000093, 5.000291, 5.000842, 
    5.002254, 5.005562, 5.012565, 5.025754, 5.047345, 5.076943, 5.108829, 0, 
    6.720564, 6.584433, 6.289873, 5.876649, 5.422355, 4.96215, 4.566208, 
    4.253551, 4.049467, 3.975818, 4.036649, 4.214753, 4.470621, 4.757757, 
    5.04374, 5.27896, 5.498487, 5.692443, 5.846371, 5.940264, 5.951794, 
    5.867256, 5.69812, 5.488389, 5.29539, 5.155908, 5.073154, 5.0311, 
    5.012152, 5.004404, 5.001488, 5.000471, 5.000139, 5.000038,
  // height(3,29, 0-49)
    5, 5, 5.000004, 5.000016, 5.000057, 5.000186, 5.000579, 5.001659, 
    5.004405, 5.010764, 5.024003, 5.048273, 5.086257, 5.134563, 5.180684, 0, 
    6.556565, 6.454806, 6.209808, 5.869759, 5.502885, 5.139183, 4.826483, 
    4.584808, 4.432256, 4.377896, 4.422847, 4.556728, 4.757828, 4.99201, 
    5.226871, 5.426193, 5.607547, 5.760535, 5.869822, 5.915688, 5.880161, 
    5.75981, 5.578391, 5.383534, 5.221547, 5.112823, 5.05154, 5.021459, 
    5.008235, 5.002935, 5.000975, 5.000303, 5.000089, 5.000024,
  // height(3,30, 0-49)
    5, 5.000002, 5.000008, 5.000027, 5.0001, 5.000338, 5.001072, 5.003178, 
    5.008781, 5.022519, 5.053143, 5.113769, 5.216212, 5.355342, 5.494076, 
    5.709598, 6.125762, 6.156536, 6.034242, 5.81732, 5.566053, 5.311934, 
    5.084235, 4.906974, 4.7975, 4.758753, 4.791675, 4.890025, 5.043805, 
    5.226883, 5.40879, 5.569041, 5.707834, 5.814003, 5.871604, 5.863268, 
    5.779329, 5.629799, 5.448622, 5.279824, 5.153577, 5.075142, 5.033274, 
    5.013503, 5.005065, 5.001767, 5.000576, 5.000175, 5.000051, 5.000014,
  // height(3,31, 0-49)
    5, 5.000001, 5.000006, 5.000023, 5.000086, 5.000294, 5.000936, 5.002785, 
    5.007725, 5.019886, 5.047167, 5.101953, 5.197631, 5.337241, 5.499212, 
    5.707389, 6.101362, 6.130861, 6.032712, 5.862597, 5.666519, 5.477023, 
    5.3025, 5.166655, 5.086007, 5.057975, 5.082697, 5.156963, 5.279002, 
    5.426205, 5.569045, 5.70021, 5.80257, 5.863031, 5.866385, 5.801664, 
    5.672307, 5.502812, 5.331985, 5.193449, 5.100338, 5.046923, 5.020027, 
    5.007874, 5.00287, 5.000974, 5.000309, 5.000092, 5.000025, 5.000007,
  // height(3,32, 0-49)
    5, 5, 5.000003, 5.000016, 5.000057, 5.000198, 5.000641, 5.001941, 
    5.005484, 5.014384, 5.034873, 5.077482, 5.155878, 5.27987, 5.442998, 
    5.649105, 5.993998, 6.054826, 6.009722, 5.902009, 5.764829, 5.636314, 
    5.511456, 5.412694, 5.356704, 5.337633, 5.354934, 5.407454, 5.49851, 
    5.607553, 5.707836, 5.802571, 5.86004, 5.867137, 5.813318, 5.698636, 
    5.540854, 5.372893, 5.228083, 5.124352, 5.061041, 5.027278, 5.011199, 
    5.004254, 5.001501, 5.000495, 5.000153, 5.000045, 5.000013, 5.000002,
  // height(3,33, 0-49)
    5, 5, 5.000001, 5.000009, 5.000031, 5.000113, 5.000374, 5.00116, 
    5.003356, 5.009038, 5.022561, 5.051877, 5.108922, 5.206487, 5.349631, 
    5.540675, 5.829793, 5.934906, 5.95664, 5.919773, 5.845279, 5.775891, 
    5.699202, 5.635369, 5.600927, 5.589468, 5.600031, 5.632689, 5.692454, 
    5.760539, 5.814003, 5.863031, 5.867137, 5.816883, 5.711125, 5.563231, 
    5.400769, 5.25464, 5.144711, 5.0741, 5.034512, 5.014745, 5.005819, 
    5.00213, 5.000726, 5.000232, 5.00007, 5.00002, 5.000005, 5,
  // height(3,34, 0-49)
    5, 5, 5, 5.000003, 5.000016, 5.000058, 5.000192, 5.000611, 5.001822, 
    5.00506, 5.013054, 5.031149, 5.068315, 5.13659, 5.246739, 5.405913, 
    5.637955, 5.777564, 5.862308, 5.896429, 5.887648, 5.877523, 5.849693, 
    5.821001, 5.806437, 5.801769, 5.806009, 5.819705, 5.846376, 5.869823, 
    5.871605, 5.866385, 5.813318, 5.711125, 5.5706, 5.414839, 5.271254, 
    5.159427, 5.084641, 5.040899, 5.018124, 5.00741, 5.002808, 5.000989, 
    5.000327, 5.000101, 5.00003, 5.000008, 5.000001, 5,
  // height(3,35, 0-49)
    5, 5, 5, 5.000001, 5.000007, 5.000026, 5.000089, 5.00029, 5.000893, 
    5.002561, 5.006839, 5.016948, 5.038792, 5.081545, 5.156356, 5.273779, 
    5.448004, 5.596495, 5.722991, 5.816328, 5.870923, 5.919303, 5.941797, 
    5.950219, 5.955517, 5.957448, 5.955325, 5.949628, 5.940266, 5.915689, 
    5.863268, 5.801664, 5.698636, 5.56323, 5.414839, 5.276899, 5.167127, 
    5.091476, 5.045663, 5.020916, 5.00884, 5.003462, 5.001259, 5.000427, 
    5.000136, 5.000041, 5.000012, 5.000003, 5, 5,
  // height(3,36, 0-49)
    5, 5, 5, 5, 5.000002, 5.000011, 5.000038, 5.000125, 5.000399, 5.001182, 
    5.00327, 5.008418, 5.020082, 5.044224, 5.089479, 5.166116, 5.285483, 
    5.41548, 5.55173, 5.678836, 5.782701, 5.881738, 5.952456, 5.998994, 
    6.024836, 6.033529, 6.024755, 5.998743, 5.951795, 5.880162, 5.77933, 
    5.672307, 5.540854, 5.400769, 5.271254, 5.167127, 5.093842, 5.048205, 
    5.022761, 5.009921, 5.004006, 5.001504, 5.000525, 5.000171, 5.000052, 
    5.000016, 5.000004, 5, 5, 5,
  // height(3,37, 0-49)
    5, 5, 5, 5, 5, 5.000004, 5.000015, 5.000051, 5.000163, 5.000501, 
    5.001435, 5.003837, 5.00953, 5.021924, 5.046564, 5.091146, 5.164802, 
    5.260377, 5.377213, 5.50543, 5.631152, 5.760442, 5.867519, 5.947026, 
    5.991995, 6.007086, 5.991962, 5.946927, 5.867255, 5.75981, 5.629799, 
    5.502812, 5.372893, 5.25464, 5.159427, 5.091476, 5.048205, 5.023404, 
    5.010503, 5.004369, 5.001688, 5.000608, 5.000204, 5.000064, 5.00002, 
    5.000005, 5, 5, 5, 5,
  // height(3,38, 0-49)
    5, 5, 5, 5, 5, 5, 5.000005, 5.00002, 5.000062, 5.000195, 5.00058, 
    5.001613, 5.004166, 5.009988, 5.022183, 5.045549, 5.086459, 5.146701, 
    5.229607, 5.33292, 5.449109, 5.578621, 5.698215, 5.795055, 5.852177, 
    5.871556, 5.852166, 5.79502, 5.69812, 5.578392, 5.448622, 5.331985, 
    5.228083, 5.144711, 5.084641, 5.045663, 5.022761, 5.010503, 5.004496, 
    5.001788, 5.000662, 5.000228, 5.000074, 5.000023, 5.000007, 5.000001, 5, 
    5, 5, 5,
  // height(3,39, 0-49)
    5, 5, 5, 5, 5, 5, 5.000001, 5.000007, 5.000022, 5.000071, 5.000218, 
    5.000627, 5.001684, 5.004201, 5.00973, 5.020876, 5.04146, 5.074723, 
    5.124831, 5.193744, 5.27998, 5.383608, 5.48842, 5.579863, 5.636596, 
    5.656175, 5.636593, 5.57985, 5.488389, 5.383535, 5.279824, 5.193449, 
    5.124352, 5.0741, 5.040899, 5.020916, 5.009921, 5.004369, 5.001788, 
    5.000681, 5.000242, 5.00008, 5.000025, 5.000008, 5.000002, 5, 5, 5, 5, 5,
  // height(3,40, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000008, 5.000024, 5.000075, 5.000226, 
    5.00063, 5.001637, 5.003948, 5.008826, 5.018284, 5.034691, 5.061178, 
    5.100423, 5.153621, 5.221567, 5.295398, 5.363819, 5.408352, 5.423996, 
    5.408351, 5.363815, 5.29539, 5.221547, 5.153577, 5.100338, 5.061041, 
    5.034512, 5.018124, 5.00884, 5.004006, 5.001688, 5.000662, 5.000242, 
    5.000082, 5.000026, 5.000008, 5.000002, 5, 5, 5, 5, 5, 5,
  // height(3,41, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000008, 5.000024, 5.000076, 5.00022, 
    5.000594, 5.001486, 5.003456, 5.007452, 5.014793, 5.027314, 5.046945, 
    5.075154, 5.112829, 5.15591, 5.197577, 5.225729, 5.235758, 5.225728, 
    5.197576, 5.155908, 5.112823, 5.075142, 5.046923, 5.027278, 5.014745, 
    5.00741, 5.003462, 5.001504, 5.000608, 5.000228, 5.00008, 5.000026, 
    5.000009, 5.000002, 5, 5, 5, 5, 5, 5, 5,
  // height(3,42, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000008, 5.000024, 5.000072, 
    5.0002, 5.000521, 5.001258, 5.002819, 5.00583, 5.011209, 5.020034, 
    5.033277, 5.051541, 5.073155, 5.094623, 5.109491, 5.114835, 5.109491, 
    5.094623, 5.073154, 5.05154, 5.033274, 5.020027, 5.011199, 5.005819, 
    5.002808, 5.001259, 5.000525, 5.000204, 5.000074, 5.000025, 5.000008, 
    5.000002, 5, 5, 5, 5, 5, 5, 5, 5,
  // height(3,43, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000008, 5.000023, 5.000063, 
    5.00017, 5.000428, 5.000993, 5.002134, 5.004256, 5.007876, 5.013503, 
    5.021459, 5.0311, 5.040833, 5.047673, 5.050141, 5.047673, 5.040833, 
    5.0311, 5.021459, 5.013503, 5.007874, 5.004254, 5.00213, 5.000989, 
    5.000427, 5.000171, 5.000064, 5.000023, 5.000008, 5.000002, 5, 5, 5, 5, 
    5, 5, 5, 5, 5,
  // height(3,44, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000007, 5.00002, 5.000052, 
    5.000136, 5.000328, 5.000727, 5.001502, 5.002871, 5.005065, 5.008235, 
    5.012152, 5.016148, 5.018981, 5.020005, 5.018981, 5.016148, 5.012152, 
    5.008235, 5.005065, 5.00287, 5.001501, 5.000726, 5.000327, 5.000136, 
    5.000052, 5.00002, 5.000007, 5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // height(3,45, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000005, 5.000016, 
    5.000041, 5.000101, 5.000232, 5.000495, 5.000975, 5.001767, 5.002935, 
    5.004404, 5.005916, 5.006993, 5.007383, 5.006993, 5.005916, 5.004404, 
    5.002935, 5.001767, 5.000974, 5.000495, 5.000232, 5.000101, 5.000041, 
    5.000016, 5.000005, 5.000001, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // height(3,46, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000004, 5.000012, 5.00003, 
    5.00007, 5.000153, 5.000309, 5.000576, 5.000975, 5.001488, 5.002019, 
    5.0024, 5.002537, 5.0024, 5.002019, 5.001488, 5.000975, 5.000576, 
    5.000309, 5.000153, 5.00007, 5.00003, 5.000012, 5.000004, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5,
  // height(3,47, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000003, 5.000008, 5.00002, 
    5.000045, 5.000092, 5.000175, 5.000303, 5.000471, 5.000645, 5.000771, 
    5.000815, 5.000771, 5.000645, 5.000471, 5.000303, 5.000175, 5.000092, 
    5.000045, 5.00002, 5.000008, 5.000003, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5,
  // height(3,48, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000005, 
    5.000013, 5.000025, 5.000051, 5.000089, 5.000139, 5.000192, 5.000231, 
    5.000245, 5.000231, 5.000192, 5.000139, 5.000089, 5.000051, 5.000025, 
    5.000013, 5.000005, 5.000001, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // height(3,49, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000006, 
    5.000012, 5.000023, 5.000038, 5.000055, 5.000067, 5.000071, 5.000067, 
    5.000055, 5.000038, 5.000023, 5.000012, 5.000006, 5.000002, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // height(4,0, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000006, 5.000013, 
    5.000028, 5.000057, 5.000112, 5.000206, 5.000354, 5.000569, 5.00085, 
    5.001171, 5.001479, 5.001697, 5.001776, 5.001697, 5.001479, 5.001171, 
    5.00085, 5.000569, 5.000354, 5.000206, 5.000112, 5.000057, 5.000028, 
    5.000013, 5.000006, 5.000001, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // height(4,1, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000003, 5.000008, 5.000018, 5.000039, 
    5.000082, 5.000166, 5.000319, 5.000575, 5.000974, 5.001544, 5.002285, 
    5.003127, 5.003933, 5.004504, 5.00471, 5.004504, 5.003933, 5.003127, 
    5.002285, 5.001544, 5.000974, 5.000575, 5.000319, 5.000166, 5.000082, 
    5.000038, 5.000018, 5.000008, 5.000003, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // height(4,2, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000004, 5.00001, 5.000022, 5.00005, 
    5.000111, 5.000235, 5.000467, 5.000876, 5.001545, 5.002564, 5.003994, 
    5.005826, 5.00789, 5.009855, 5.011244, 5.011746, 5.011244, 5.009855, 
    5.00789, 5.005825, 5.003993, 5.002563, 5.001543, 5.000874, 5.000466, 
    5.000235, 5.000111, 5.00005, 5.000022, 5.00001, 5.000004, 5, 5, 5, 5, 5, 
    5, 5, 5, 5,
  // height(4,3, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000005, 5.000011, 5.000026, 5.000062, 
    5.000142, 5.000312, 5.000645, 5.001252, 5.002286, 5.003933, 5.006382, 
    5.00975, 5.014007, 5.018755, 5.023253, 5.026416, 5.027557, 5.026416, 
    5.023252, 5.018755, 5.014006, 5.009748, 5.006378, 5.003928, 5.002279, 
    5.001247, 5.000645, 5.000314, 5.000144, 5.000063, 5.000027, 5.000011, 
    5.000005, 5.000001, 5, 5, 5, 5, 5, 5, 5,
  // height(4,4, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000005, 5.000012, 5.00003, 5.000073, 
    5.000174, 5.000391, 5.000835, 5.001678, 5.003172, 5.005635, 5.009448, 
    5.014966, 5.022386, 5.031617, 5.041789, 5.051358, 5.058033, 5.060435, 
    5.058033, 5.051356, 5.041786, 5.031611, 5.022377, 5.014951, 5.009429, 
    5.005613, 5.003155, 5.001675, 5.00084, 5.000397, 5.000178, 5.000076, 
    5.000031, 5.000013, 5.000005, 5.000001, 5, 5, 5, 5, 5, 5,
  // height(4,5, 0-49)
    5, 5, 5, 5, 5, 5, 5.000002, 5.000006, 5.000013, 5.000031, 5.000082, 
    5.0002, 5.000464, 5.00102, 5.002115, 5.004128, 5.00759, 5.013093, 
    5.021336, 5.032907, 5.048047, 5.066521, 5.086531, 5.105149, 5.117974, 
    5.122565, 5.117973, 5.105145, 5.086521, 5.066501, 5.048014, 5.032856, 
    5.021269, 5.01302, 5.007533, 5.004119, 5.002128, 5.001039, 5.00048, 
    5.00021, 5.000087, 5.000034, 5.000014, 5.000006, 5.000002, 5, 5, 5, 5, 5,
  // height(4,6, 0-49)
    5, 5, 5, 5, 5, 5.000001, 5.000006, 5.000013, 5.000033, 5.000086, 
    5.000218, 5.00052, 5.001176, 5.002513, 5.005054, 5.009583, 5.017104, 
    5.028571, 5.04509, 5.06742, 5.095617, 5.129127, 5.164507, 5.196824, 
    5.218638, 5.226384, 5.218632, 5.196807, 5.164472, 5.12906, 5.095507, 
    5.067253, 5.04487, 5.028332, 5.016919, 5.009551, 5.005095, 5.002568, 
    5.001224, 5.00055, 5.000236, 5.000094, 5.000036, 5.000015, 5.000007, 
    5.000002, 5, 5, 5, 5,
  // height(4,7, 0-49)
    5, 5, 5, 5, 5, 5.000005, 5.000013, 5.000032, 5.000086, 5.000224, 
    5.000552, 5.001284, 5.002817, 5.005834, 5.011383, 5.020915, 5.036179, 
    5.058282, 5.0886, 5.12762, 5.174555, 5.228317, 5.28298, 5.331494, 
    5.363276, 5.374424, 5.363256, 5.331442, 5.282871, 5.228115, 5.174216, 
    5.12711, 5.08793, 5.057558, 5.035612, 5.020813, 5.011489, 5.00599, 
    5.002948, 5.001372, 5.000603, 5.00025, 5.000099, 5.000037, 5.000015, 
    5.000006, 5.000001, 5, 5, 5,
  // height(4,8, 0-49)
    5, 5, 5, 5, 5.000004, 5.000011, 5.00003, 5.000083, 5.000219, 5.000553, 
    5.001321, 5.002983, 5.00635, 5.012745, 5.024074, 5.042771, 5.071508, 
    5.110453, 5.160557, 5.220954, 5.288945, 5.363122, 5.434719, 5.495795, 
    5.534249, 5.547521, 5.534192, 5.49565, 5.434417, 5.36256, 5.288007, 
    5.219527, 5.158675, 5.108407, 5.069887, 5.04248, 5.024346, 5.013159, 
    5.006711, 5.003231, 5.001469, 5.000631, 5.000257, 5.000099, 5.000036, 
    5.000014, 5.000005, 5.000001, 5, 5,
  // height(4,9, 0-49)
    5, 5, 5, 5.000003, 5.00001, 5.000027, 5.000073, 5.000201, 5.000522, 
    5.001283, 5.002978, 5.006522, 5.013456, 5.026117, 5.047627, 5.081541, 
    5.131313, 5.193063, 5.26604, 5.346703, 5.429886, 5.515448, 5.592755, 
    5.65555, 5.693194, 5.705945, 5.693052, 5.655185, 5.592003, 5.51405, 
    5.427536, 5.343099, 5.261235, 5.187773, 5.12704, 5.0808, 5.048308, 
    5.027168, 5.014386, 5.00718, 5.00338, 5.001504, 5.000631, 5.00025, 
    5.000094, 5.000034, 5.000013, 5.000005, 5, 5,
  // height(4,10, 0-49)
    5, 5, 5.000001, 5.000008, 5.000023, 5.000062, 5.000174, 5.000464, 
    5.001174, 5.002803, 5.006311, 5.01339, 5.026711, 5.050013, 5.087704, 
    5.143996, 5.222599, 5.309128, 5.400571, 5.490787, 5.573659, 5.653591, 
    5.720015, 5.770827, 5.799431, 5.808886, 5.799106, 5.770001, 5.718316, 
    5.65044, 5.568353, 5.482604, 5.389545, 5.296785, 5.212377, 5.142366, 
    5.089346, 5.052536, 5.028989, 5.015037, 5.007341, 5.00338, 5.001469, 
    5.000603, 5.000236, 5.000087, 5.000031, 5.000011, 5.000004, 5,
  // height(4,11, 0-49)
    5, 5.000001, 5.000006, 5.000018, 5.000051, 5.000142, 5.000389, 5.00101, 
    5.002481, 5.005745, 5.012537, 5.025723, 5.049498, 5.089058, 5.149407, 
    5.233919, 5.346392, 5.451672, 5.547588, 5.628493, 5.690985, 5.747229, 
    5.788034, 5.816257, 5.830287, 5.834641, 5.829595, 5.814518, 5.784492, 
    5.740716, 5.680092, 5.611754, 5.524933, 5.425946, 5.324495, 5.230956, 
    5.153233, 5.094786, 5.05476, 5.029618, 5.015037, 5.00718, 5.003231, 
    5.001372, 5.00055, 5.00021, 5.000076, 5.000027, 5.00001, 5.000003,
  // height(4,12, 0-49)
    5, 5.000003, 5.000013, 5.000038, 5.000109, 5.000305, 5.000814, 5.002055, 
    5.004901, 5.011015, 5.023273, 5.046094, 5.08526, 5.146695, 5.233996, 
    5.347453, 5.493467, 5.603019, 5.683767, 5.735504, 5.761001, 5.781113, 
    5.78789, 5.788424, 5.785759, 5.784305, 5.784378, 5.784986, 5.780982, 
    5.768596, 5.740397, 5.704315, 5.641876, 5.555245, 5.451858, 5.343374, 
    5.242486, 5.158862, 5.096653, 5.05476, 5.028989, 5.014386, 5.006711, 
    5.002948, 5.001224, 5.00048, 5.000178, 5.000063, 5.000022, 5.000008,
  // height(4,13, 0-49)
    5.000001, 5.000009, 5.000026, 5.000077, 5.000224, 5.000611, 5.001587, 
    5.003901, 5.009038, 5.019696, 5.040237, 5.07673, 5.135884, 5.222372, 
    5.33526, 5.470407, 5.644621, 5.740721, 5.789155, 5.798397, 5.778439, 
    5.757261, 5.727443, 5.699325, 5.679906, 5.672492, 5.677281, 5.692876, 
    5.71471, 5.734662, 5.742108, 5.744841, 5.718772, 5.661288, 5.574646, 
    5.467301, 5.352917, 5.246391, 5.158862, 5.094786, 5.052536, 5.027167, 
    5.013159, 5.00599, 5.002568, 5.001039, 5.000397, 5.000144, 5.00005, 
    5.000018,
  // height(4,14, 0-49)
    5.000004, 5.000016, 5.000051, 5.00015, 5.000423, 5.001134, 5.002876, 
    5.006879, 5.015491, 5.032723, 5.064547, 5.118182, 5.199555, 5.309104, 
    5.438466, 5.581018, 5.776528, 5.845946, 5.853991, 5.817026, 5.75099, 
    5.688416, 5.622475, 5.56643, 5.530651, 5.517122, 5.525881, 5.554883, 
    5.600159, 5.649828, 5.690797, 5.731436, 5.745387, 5.726641, 5.672071, 
    5.58408, 5.472425, 5.352917, 5.242486, 5.153233, 5.089346, 5.048308, 
    5.024346, 5.011489, 5.005095, 5.002128, 5.00084, 5.000314, 5.000111, 
    5.000039,
  // height(4,15, 0-49)
    5.000009, 5.00003, 5.000093, 5.000268, 5.000741, 5.001943, 5.004808, 
    5.011213, 5.02456, 5.050291, 5.095673, 5.167803, 5.269303, 5.393564, 
    5.523967, 5.657652, 5.868953, 5.907986, 5.878179, 5.799743, 5.692262, 
    5.590435, 5.489555, 5.406311, 5.354075, 5.333925, 5.345757, 5.386508, 
    5.452232, 5.527853, 5.598085, 5.67159, 5.722934, 5.744675, 5.730055, 
    5.67552, 5.58408, 5.467301, 5.343374, 5.230956, 5.142365, 5.080799, 
    5.04248, 5.020813, 5.009551, 5.004119, 5.001675, 5.000645, 5.000236, 
    5.000084,
  // height(4,16, 0-49)
    5.000016, 5.000051, 5.000154, 5.000436, 5.001185, 5.003041, 5.007361, 
    5.016769, 5.035784, 5.071095, 5.130445, 5.218989, 5.333667, 5.459665, 
    5.573878, 5.686548, 5.908281, 5.92311, 5.866307, 5.756901, 5.615705, 
    5.477578, 5.342819, 5.232497, 5.162915, 5.135132, 5.148944, 5.199866, 
    5.28306, 5.380913, 5.476108, 5.57633, 5.659531, 5.718256, 5.744269, 
    5.730054, 5.672071, 5.574646, 5.451857, 5.324495, 5.212377, 5.12704, 
    5.069887, 5.035612, 5.016918, 5.007533, 5.003155, 5.001247, 5.000467, 
    5.000169,
  // height(4,17, 0-49)
    5.000024, 5.000076, 5.000226, 5.000637, 5.0017, 5.004287, 5.01019, 
    5.022752, 5.047452, 5.091729, 5.162721, 5.26203, 5.379788, 5.493896, 
    5.577772, 5.66574, 5.886785, 5.890759, 5.822771, 5.696401, 5.531397, 
    5.360797, 5.193435, 5.055688, 4.967145, 4.93014, 4.944488, 5.003893, 
    5.101617, 5.218238, 5.334838, 5.456188, 5.56532, 5.655404, 5.718253, 
    5.744672, 5.726639, 5.661288, 5.555245, 5.425946, 5.296785, 5.187774, 
    5.108407, 5.057558, 5.028332, 5.01302, 5.005613, 5.00228, 5.000876, 
    5.000325,
  // height(4,18, 0-49)
    5.000031, 5.000098, 5.00029, 5.000809, 5.002132, 5.005311, 5.012467, 
    5.027443, 5.05629, 5.106589, 5.184099, 5.286392, 5.397364, 5.489583, 
    5.535452, 5.605662, 5.800894, 5.810308, 5.749249, 5.622153, 5.445377, 
    5.247847, 5.050285, 4.884759, 4.775092, 4.726635, 4.739514, 4.805339, 
    4.914531, 5.046517, 5.181646, 5.319603, 5.449533, 5.565309, 5.659521, 
    5.722928, 5.745382, 5.718771, 5.641876, 5.524933, 5.389545, 5.261234, 
    5.158674, 5.08793, 5.04487, 5.021269, 5.009429, 5.003929, 5.001545, 
    5.000584,
  // height(4,19, 0-49)
    5.000033, 5.000104, 5.000303, 5.000842, 5.002212, 5.00549, 5.012845, 
    5.02818, 5.057574, 5.108389, 5.185361, 5.283393, 5.381967, 5.449668, 
    5.45941, 5.528225, 5.651516, 5.679839, 5.644249, 5.534561, 5.360603, 
    5.14432, 4.920958, 4.727758, 4.594412, 4.531527, 4.540184, 4.609795, 
    4.727152, 4.870959, 5.022038, 5.172999, 5.319552, 5.45614, 5.576295, 
    5.67157, 5.731426, 5.744835, 5.704313, 5.611754, 5.482604, 5.343098, 
    5.219526, 5.12711, 5.067253, 5.032856, 5.014951, 5.00638, 5.002567, 
    5.000986,
  // height(4,20, 0-49)
    5.000022, 5.000071, 5.000206, 5.000566, 5.001461, 5.003547, 5.008075, 
    5.017149, 5.033758, 5.061057, 5.100434, 5.148736, 5.196876, 5.232886, 
    5.249486, 0, 5.72522, 5.722096, 5.663104, 5.536474, 5.342846, 5.092929, 
    4.832631, 4.601823, 4.436234, 4.352537, 4.352442, 4.422397, 4.544476, 
    4.696456, 4.860911, 5.021814, 5.181428, 5.334681, 5.476007, 5.598027, 
    5.690766, 5.742093, 5.74039, 5.680089, 5.568351, 5.427535, 5.288007, 
    5.174216, 5.095507, 5.048014, 5.022378, 5.00975, 5.003997, 5.001556,
  // height(4,21, 0-49)
    5.000014, 5.000044, 5.000126, 5.000348, 5.000903, 5.002204, 5.005051, 
    5.010816, 5.021541, 5.039646, 5.06693, 5.102845, 5.142964, 5.179457, 
    5.204838, 0, 5.693264, 5.683771, 5.624491, 5.49779, 5.296422, 5.020554, 
    4.725423, 4.45422, 4.252345, 4.146114, 4.139155, 4.214416, 4.347202, 
    4.512626, 4.695527, 4.870046, 5.045835, 5.217789, 5.380641, 5.527698, 
    5.649745, 5.734621, 5.768576, 5.740706, 5.650436, 5.514049, 5.36256, 
    5.228116, 5.12906, 5.066501, 5.031611, 5.014006, 5.005826, 5.002292,
  // height(4,22, 0-49)
    5.000008, 5.000024, 5.000072, 5.000199, 5.000521, 5.00129, 5.002997, 
    5.006517, 5.013214, 5.024857, 5.043125, 5.068581, 5.099402, 5.130821, 
    5.156437, 0, 5.645344, 5.631002, 5.571152, 5.445369, 5.241158, 4.948497, 
    4.63036, 4.328893, 4.096667, 3.969621, 3.954431, 4.03174, 4.170502, 
    4.343932, 4.540859, 4.72441, 4.91267, 5.100444, 5.282361, 5.451836, 
    5.599946, 5.7146, 5.780928, 5.784469, 5.718306, 5.591999, 5.434416, 
    5.28287, 5.164471, 5.086521, 5.041785, 5.018754, 5.007888, 5.003124,
  // height(4,23, 0-49)
    5.000003, 5.000014, 5.000041, 5.000118, 5.000312, 5.000783, 5.001848, 
    5.004087, 5.008446, 5.016229, 5.028857, 5.047226, 5.070715, 5.096325, 
    5.118713, 0, 5.596464, 5.578844, 5.518146, 5.392861, 5.187092, 4.88203, 
    4.546795, 4.220427, 3.96124, 3.815448, 3.794108, 3.875613, 4.021391, 
    4.202407, 4.412063, 4.602664, 4.800696, 5.001018, 5.198163, 5.385542, 
    5.554357, 5.692601, 5.784849, 5.814455, 5.769972, 5.655174, 5.495645, 
    5.33144, 5.196806, 5.105144, 5.051356, 5.023251, 5.009851, 5.003916,
  // height(4,24, 0-49)
    5.000002, 5.000011, 5.000033, 5.000093, 5.000248, 5.000626, 5.001483, 
    5.003294, 5.006839, 5.01322, 5.023686, 5.039129, 5.059257, 5.081702, 
    5.101663, 0, 5.556334, 5.537187, 5.476232, 5.351586, 5.145324, 4.83245, 
    4.485684, 4.140932, 3.860631, 3.700632, 3.676901, 3.765053, 3.9187, 
    4.106887, 4.327, 4.52336, 4.728728, 4.937836, 5.14499, 5.343493, 
    5.524635, 5.676622, 5.784046, 5.829436, 5.799034, 5.693022, 5.534179, 
    5.363252, 5.21863, 5.117971, 5.058032, 5.026413, 5.011236, 5.004478,
  // height(4,25, 0-49)
    5.000005, 5.000016, 5.000045, 5.000125, 5.000327, 5.000806, 5.00187, 
    5.004066, 5.00826, 5.015623, 5.027387, 5.044277, 5.06568, 5.088906, 
    5.109101, 0, 5.530094, 5.511153, 5.450953, 5.327627, 5.122614, 4.808633, 
    4.459426, 4.109352, 3.822037, 3.657288, 3.633398, 3.724782, 3.881723, 
    4.07268, 4.296721, 4.495244, 4.70334, 4.915673, 5.126443, 5.328887, 
    5.514308, 5.670983, 5.783531, 5.834264, 5.808712, 5.705871, 5.54749, 
    5.374413, 5.226382, 5.122564, 5.060434, 5.027554, 5.011736, 5.004682,
  // height(4,26, 0-49)
    5.00001, 5.00003, 5.000083, 5.000225, 5.000573, 5.001377, 5.003111, 
    5.006579, 5.012978, 5.023774, 5.040254, 5.062696, 5.089457, 5.116624, 
    5.138906, 0, 5.520136, 5.503262, 5.445169, 5.324215, 5.122498, 4.814704, 
    4.473166, 4.133136, 3.856438, 3.698707, 3.676142, 3.764788, 3.918613, 
    4.10686, 4.326991, 4.523357, 4.728727, 4.937836, 5.144989, 5.343493, 
    5.524634, 5.676622, 5.784046, 5.829436, 5.799034, 5.693022, 5.534179, 
    5.363252, 5.21863, 5.117971, 5.058032, 5.026413, 5.011236, 5.004478,
  // height(4,27, 0-49)
    5.000019, 5.000056, 5.000157, 5.000415, 5.001042, 5.002456, 5.005435, 
    5.011232, 5.021597, 5.038417, 5.062864, 5.094123, 5.128512, 5.160077, 
    5.183197, 0, 5.526995, 5.513671, 5.458173, 5.339542, 5.142099, 4.846486, 
    4.52138, 4.204391, 3.952483, 3.811342, 3.79244, 3.875007, 4.021184, 
    4.202338, 4.412041, 4.602656, 4.800694, 5.001017, 5.198163, 5.385541, 
    5.554357, 5.692601, 5.784849, 5.814455, 5.769972, 5.655174, 5.495645, 
    5.33144, 5.196806, 5.105144, 5.051356, 5.023251, 5.009851, 5.003916,
  // height(4,28, 0-49)
    5.000035, 5.0001, 5.000277, 5.000724, 5.001793, 5.004173, 5.009095, 
    5.018476, 5.034788, 5.060286, 5.095444, 5.137174, 5.178433, 5.210751, 
    5.229156, 0, 5.549765, 5.540964, 5.487337, 5.369511, 5.17579, 4.895623, 
    4.591888, 4.304254, 4.082989, 3.963053, 3.951664, 4.030686, 4.170128, 
    4.343802, 4.540814, 4.724395, 4.912664, 5.100442, 5.28236, 5.451836, 
    5.599946, 5.7146, 5.780928, 5.784469, 5.718305, 5.591999, 5.434416, 
    5.28287, 5.164471, 5.086521, 5.041785, 5.018754, 5.007888, 5.003124,
  // height(4,29, 0-49)
    5.000054, 5.000159, 5.000442, 5.001153, 5.00284, 5.006568, 5.014205, 
    5.028555, 5.05294, 5.08968, 5.137436, 5.189026, 5.232651, 5.257787, 
    5.262488, 0, 5.584862, 5.579939, 5.525392, 5.405305, 5.214372, 4.952533, 
    4.675216, 4.421723, 4.234072, 4.137152, 4.135252, 4.212865, 4.346626, 
    4.51242, 4.695455, 4.870021, 5.045825, 5.217786, 5.380639, 5.527698, 
    5.649745, 5.734621, 5.768576, 5.740706, 5.650436, 5.514049, 5.36256, 
    5.228116, 5.12906, 5.066501, 5.031611, 5.014006, 5.005826, 5.002292,
  // height(4,30, 0-49)
    5.000076, 5.000227, 5.000637, 5.001688, 5.004233, 5.010009, 5.022226, 
    5.046075, 5.08837, 5.154881, 5.244466, 5.342824, 5.423133, 5.457164, 
    5.429102, 5.460217, 5.513269, 5.527208, 5.492916, 5.390181, 5.221525, 
    4.998848, 4.766492, 4.560466, 4.413423, 4.341393, 4.347546, 4.42042, 
    4.543725, 4.696185, 4.860814, 5.02178, 5.181416, 5.334677, 5.476006, 
    5.598026, 5.690766, 5.742093, 5.74039, 5.680089, 5.568351, 5.427535, 
    5.288007, 5.174216, 5.095507, 5.048014, 5.022378, 5.00975, 5.003997, 
    5.001556,
  // height(4,31, 0-49)
    5.000073, 5.000221, 5.000621, 5.001653, 5.00416, 5.009876, 5.02202, 
    5.045835, 5.088351, 5.155962, 5.249051, 5.356033, 5.453192, 5.513427, 
    5.51753, 5.549628, 5.688647, 5.683352, 5.618227, 5.4899, 5.309708, 
    5.098572, 4.885837, 4.704521, 4.580997, 4.524658, 4.537004, 4.608436, 
    4.726605, 4.870749, 5.021959, 5.17297, 5.319542, 5.456137, 5.576294, 
    5.671569, 5.731426, 5.744835, 5.704313, 5.611754, 5.482604, 5.343098, 
    5.219526, 5.12711, 5.067253, 5.032856, 5.014951, 5.00638, 5.002567, 
    5.000986,
  // height(4,32, 0-49)
    5.000058, 5.000175, 5.000499, 5.001343, 5.003422, 5.008226, 5.018595, 
    5.039321, 5.077241, 5.13961, 5.229686, 5.340741, 5.453701, 5.542929, 
    5.586711, 5.634364, 5.810377, 5.794869, 5.715106, 5.578702, 5.402011, 
    5.211908, 5.024439, 4.868459, 4.765963, 4.722025, 4.737376, 4.804413, 
    4.91415, 5.046367, 5.181589, 5.319583, 5.449525, 5.565306, 5.65952, 
    5.722928, 5.745382, 5.718771, 5.641876, 5.524932, 5.389545, 5.261234, 
    5.158674, 5.08793, 5.04487, 5.021269, 5.009429, 5.003929, 5.001545, 
    5.000584,
  // height(4,33, 0-49)
    5.00004, 5.000121, 5.000348, 5.000955, 5.002475, 5.006059, 5.013967, 
    5.030193, 5.060858, 5.113483, 5.193935, 5.30105, 5.422253, 5.535433, 
    5.617548, 5.69124, 5.875936, 5.864213, 5.786301, 5.657351, 5.496267, 
    5.333714, 5.17509, 5.044634, 4.961142, 4.927159, 4.943112, 5.003295, 
    5.101369, 5.218139, 5.334802, 5.456174, 5.565315, 5.655402, 5.718253, 
    5.744672, 5.726639, 5.661288, 5.555245, 5.425946, 5.296785, 5.187774, 
    5.108407, 5.057558, 5.028332, 5.01302, 5.005613, 5.00228, 5.000876, 
    5.000325,
  // height(4,34, 0-49)
    5.000024, 5.000075, 5.000218, 5.000609, 5.001614, 5.004035, 5.009521, 
    5.021117, 5.043819, 5.084566, 5.150602, 5.245469, 5.363938, 5.490148, 
    5.602442, 5.704795, 5.886364, 5.892461, 5.832005, 5.724312, 5.588806, 
    5.458125, 5.330325, 5.225271, 5.159105, 5.133275, 5.148096, 5.1995, 
    5.282907, 5.380851, 5.476084, 5.576321, 5.659528, 5.718254, 5.744268, 
    5.730054, 5.672071, 5.574646, 5.451857, 5.324495, 5.212377, 5.12704, 
    5.069887, 5.035612, 5.016918, 5.007533, 5.003155, 5.001247, 5.000467, 
    5.000169,
  // height(4,35, 0-49)
    5.000014, 5.000041, 5.000124, 5.000355, 5.000961, 5.002462, 5.00596, 
    5.013583, 5.029061, 5.058093, 5.107836, 5.184575, 5.289448, 5.414499, 
    5.54309, 5.668658, 5.844255, 5.878744, 5.849082, 5.774486, 5.672875, 
    5.577171, 5.48142, 5.401774, 5.351748, 5.332812, 5.345255, 5.386293, 
    5.452143, 5.527818, 5.598071, 5.671585, 5.722932, 5.744674, 5.730054, 
    5.67552, 5.58408, 5.467301, 5.343374, 5.230956, 5.142365, 5.080799, 
    5.04248, 5.020813, 5.009551, 5.004119, 5.001675, 5.000645, 5.000236, 
    5.000084,
  // height(4,36, 0-49)
    5.000007, 5.000022, 5.000065, 5.00019, 5.000528, 5.001387, 5.003449, 
    5.008088, 5.01785, 5.036942, 5.071377, 5.128031, 5.211954, 5.322424, 
    5.450345, 5.586574, 5.754741, 5.821698, 5.831575, 5.79887, 5.73787, 
    5.679853, 5.617424, 5.563701, 5.529284, 5.51648, 5.525597, 5.554762, 
    5.600111, 5.649807, 5.69079, 5.731433, 5.745385, 5.72664, 5.672071, 
    5.58408, 5.472425, 5.352917, 5.242486, 5.153233, 5.089346, 5.048308, 
    5.024346, 5.011489, 5.005095, 5.002128, 5.00084, 5.000314, 5.000111, 
    5.000039,
  // height(4,37, 0-49)
    5.000002, 5.000011, 5.000032, 5.000094, 5.00027, 5.000727, 5.001855, 
    5.004479, 5.010196, 5.021828, 5.043808, 5.082083, 5.142909, 5.230166, 
    5.342067, 5.472644, 5.628459, 5.722989, 5.773468, 5.786318, 5.77012, 
    5.752038, 5.724462, 5.697757, 5.679138, 5.672138, 5.677126, 5.692811, 
    5.714684, 5.734652, 5.742105, 5.744839, 5.718772, 5.661288, 5.574646, 
    5.467301, 5.352917, 5.246391, 5.158862, 5.094786, 5.052536, 5.027167, 
    5.013159, 5.00599, 5.002568, 5.001039, 5.000397, 5.000144, 5.00005, 
    5.000018,
  // height(4,38, 0-49)
    5, 5.000005, 5.000015, 5.000044, 5.000129, 5.000355, 5.000931, 5.002315, 
    5.005435, 5.012023, 5.025013, 5.048794, 5.088931, 5.150884, 5.237588, 
    5.348084, 5.483159, 5.591568, 5.673834, 5.728097, 5.756079, 5.778114, 
    5.786222, 5.787565, 5.785347, 5.784119, 5.784297, 5.784952, 5.780969, 
    5.768591, 5.740396, 5.704315, 5.641877, 5.555245, 5.451857, 5.343374, 
    5.242486, 5.158862, 5.096653, 5.05476, 5.028989, 5.014386, 5.006711, 
    5.002948, 5.001224, 5.00048, 5.000178, 5.000063, 5.000022, 5.000008,
  // height(4,39, 0-49)
    5, 5.000001, 5.000007, 5.00002, 5.000057, 5.000163, 5.000438, 5.00112, 
    5.002711, 5.006193, 5.013331, 5.026992, 5.051274, 5.091135, 5.151162, 
    5.233976, 5.340683, 5.445152, 5.541938, 5.624341, 5.688284, 5.745618, 
    5.787155, 5.815814, 5.830077, 5.834549, 5.829556, 5.814503, 5.784487, 
    5.740712, 5.680091, 5.611754, 5.524933, 5.425946, 5.324495, 5.230956, 
    5.153233, 5.094786, 5.05476, 5.029618, 5.015037, 5.00718, 5.003231, 
    5.001372, 5.00055, 5.00021, 5.000076, 5.000027, 5.00001, 5.000003,
  // height(4,40, 0-49)
    5, 5, 5.000002, 5.000009, 5.000025, 5.00007, 5.000193, 5.000509, 
    5.001269, 5.002991, 5.006652, 5.013947, 5.027512, 5.050968, 5.088504, 
    5.143935, 5.219826, 5.305856, 5.397701, 5.488678, 5.572298, 5.652788, 
    5.719582, 5.770612, 5.799332, 5.808841, 5.799087, 5.769994, 5.718313, 
    5.650439, 5.568352, 5.482605, 5.389545, 5.296785, 5.212377, 5.142365, 
    5.089346, 5.052536, 5.028989, 5.015037, 5.007341, 5.00338, 5.001469, 
    5.000603, 5.000236, 5.000087, 5.000031, 5.000011, 5.000004, 5,
  // height(4,41, 0-49)
    5, 5, 5, 5.000003, 5.000011, 5.000029, 5.000081, 5.000217, 5.000558, 
    5.001357, 5.003117, 5.006752, 5.013795, 5.026531, 5.047973, 5.081492, 
    5.130116, 5.191607, 5.264742, 5.345742, 5.429265, 5.515083, 5.592558, 
    5.655453, 5.693151, 5.705927, 5.693044, 5.655183, 5.592001, 5.51405, 
    5.427535, 5.343099, 5.261235, 5.187774, 5.12704, 5.080799, 5.048308, 
    5.027167, 5.014386, 5.00718, 5.00338, 5.001504, 5.000631, 5.00025, 
    5.000094, 5.000034, 5.000013, 5.000005, 5, 5,
  // height(4,42, 0-49)
    5, 5, 5, 5, 5.000005, 5.000012, 5.000032, 5.000088, 5.000232, 5.00058, 
    5.001373, 5.003073, 5.006487, 5.012912, 5.024214, 5.042749, 5.071041, 
    5.10987, 5.16003, 5.220561, 5.28869, 5.362971, 5.434639, 5.495757, 
    5.534231, 5.547513, 5.534188, 5.495649, 5.434417, 5.36256, 5.288007, 
    5.219526, 5.158674, 5.108407, 5.069887, 5.04248, 5.024346, 5.013159, 
    5.006711, 5.003231, 5.001469, 5.000631, 5.000257, 5.000099, 5.000036, 
    5.000014, 5.000005, 5.000001, 5, 5,
  // height(4,43, 0-49)
    5, 5, 5, 5, 5.000001, 5.000005, 5.000013, 5.000034, 5.000092, 5.000234, 
    5.000571, 5.001317, 5.002868, 5.005898, 5.011437, 5.020907, 5.036011, 
    5.058069, 5.088407, 5.127475, 5.17446, 5.228262, 5.28295, 5.331479, 
    5.36327, 5.374421, 5.363255, 5.331441, 5.28287, 5.228115, 5.174216, 
    5.12711, 5.08793, 5.057558, 5.035612, 5.020813, 5.011489, 5.00599, 
    5.002948, 5.001372, 5.000603, 5.00025, 5.000099, 5.000037, 5.000015, 
    5.000006, 5.000001, 5, 5, 5,
  // height(4,44, 0-49)
    5, 5, 5, 5, 5, 5.000001, 5.000006, 5.000014, 5.000034, 5.00009, 5.000225, 
    5.000533, 5.001195, 5.002535, 5.005076, 5.009581, 5.017048, 5.028498, 
    5.045024, 5.067372, 5.095585, 5.129107, 5.164498, 5.196819, 5.218636, 
    5.226383, 5.218631, 5.196807, 5.164472, 5.12906, 5.095506, 5.067253, 
    5.044869, 5.028332, 5.016918, 5.009551, 5.005095, 5.002568, 5.001224, 
    5.00055, 5.000236, 5.000094, 5.000036, 5.000015, 5.000007, 5.000002, 5, 
    5, 5, 5,
  // height(4,45, 0-49)
    5, 5, 5, 5, 5, 5, 5.000002, 5.000006, 5.000013, 5.000032, 5.000083, 
    5.000204, 5.000471, 5.001028, 5.002122, 5.004128, 5.007573, 5.013069, 
    5.021315, 5.032892, 5.048037, 5.066514, 5.086528, 5.105148, 5.117975, 
    5.122566, 5.117973, 5.105145, 5.086521, 5.0665, 5.048013, 5.032856, 
    5.021268, 5.013019, 5.007533, 5.004119, 5.002128, 5.001039, 5.00048, 
    5.00021, 5.000087, 5.000034, 5.000014, 5.000006, 5.000002, 5, 5, 5, 5, 5,
  // height(4,46, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000005, 5.000012, 5.00003, 5.000074, 
    5.000175, 5.000395, 5.000838, 5.001678, 5.003167, 5.005628, 5.009441, 
    5.01496, 5.022381, 5.031613, 5.041788, 5.051359, 5.058036, 5.060439, 
    5.058036, 5.051358, 5.041786, 5.03161, 5.022376, 5.014949, 5.009427, 
    5.005613, 5.003155, 5.001675, 5.00084, 5.000397, 5.000178, 5.000076, 
    5.000031, 5.000013, 5.000005, 5.000001, 5, 5, 5, 5, 5, 5,
  // height(4,47, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000005, 5.000011, 5.000026, 5.000062, 
    5.000143, 5.000313, 5.000644, 5.001248, 5.002281, 5.003928, 5.006376, 
    5.009744, 5.014003, 5.018755, 5.023259, 5.026426, 5.027568, 5.026426, 
    5.023259, 5.018755, 5.014002, 5.009743, 5.006373, 5.003924, 5.002277, 
    5.001245, 5.000643, 5.000314, 5.000143, 5.000063, 5.000027, 5.000011, 
    5.000005, 5.000001, 5, 5, 5, 5, 5, 5, 5,
  // height(4,48, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000004, 5.00001, 5.000022, 5.000049, 
    5.000109, 5.000232, 5.000462, 5.000867, 5.001534, 5.002549, 5.003979, 
    5.005815, 5.007891, 5.009873, 5.011274, 5.01178, 5.011274, 5.009873, 
    5.007891, 5.005815, 5.003978, 5.002548, 5.001532, 5.000866, 5.000462, 
    5.000232, 5.000109, 5.000049, 5.000022, 5.00001, 5.000004, 5, 5, 5, 5, 5, 
    5, 5, 5, 5,
  // height(4,49, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000005, 5.000012, 5.00003, 
    5.000065, 5.000139, 5.000275, 5.000512, 5.000896, 5.001465, 5.002233, 
    5.00314, 5.004033, 5.004668, 5.004897, 5.004668, 5.004033, 5.00314, 
    5.002233, 5.001465, 5.000896, 5.000512, 5.000275, 5.000139, 5.000065, 
    5.00003, 5.000012, 5.000005, 5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // height(5,0, 0-49)
    5, 5, 5, 5, 5, 5, 5.000002, 5.000006, 5.000013, 5.000028, 5.000061, 
    5.00013, 5.000265, 5.000516, 5.00096, 5.001699, 5.002862, 5.004584, 
    5.006996, 5.010178, 5.014109, 5.018611, 5.023259, 5.027408, 5.030265, 
    5.031285, 5.030264, 5.027405, 5.023253, 5.018603, 5.014096, 5.010162, 
    5.006977, 5.004565, 5.002849, 5.001694, 5.000961, 5.00052, 5.000268, 
    5.000132, 5.000062, 5.000028, 5.000013, 5.000006, 5.000002, 5, 5, 5, 5, 5,
  // height(5,1, 0-49)
    5, 5, 5, 5, 5, 5.000004, 5.000008, 5.000015, 5.000031, 5.000068, 
    5.000149, 5.000312, 5.000626, 5.0012, 5.002189, 5.003802, 5.006291, 
    5.0099, 5.01486, 5.021302, 5.029162, 5.038113, 5.047316, 5.055529, 
    5.06116, 5.063167, 5.061155, 5.05552, 5.047298, 5.038086, 5.029122, 
    5.021251, 5.0148, 5.00984, 5.006246, 5.003785, 5.002189, 5.001209, 
    5.000637, 5.00032, 5.000154, 5.000071, 5.000032, 5.000015, 5.000008, 
    5.000004, 5, 5, 5, 5,
  // height(5,2, 0-49)
    5, 5, 5, 5, 5.000005, 5.000009, 5.000016, 5.000033, 5.000074, 5.000168, 
    5.000363, 5.000746, 5.001466, 5.00274, 5.004883, 5.00829, 5.013408, 
    5.020618, 5.030261, 5.042474, 5.057049, 5.073393, 5.08998, 5.104668, 
    5.114639, 5.118178, 5.114626, 5.10464, 5.089929, 5.07331, 5.056931, 
    5.042319, 5.030082, 5.020443, 5.013276, 5.008237, 5.00488, 5.002761, 
    5.001492, 5.000769, 5.000379, 5.000178, 5.000082, 5.000035, 5.000017, 
    5.000009, 5.000005, 5.000001, 5, 5,
  // height(5,3, 0-49)
    5, 5, 5, 5.000004, 5.000009, 5.000016, 5.000034, 5.000081, 5.000184, 
    5.000405, 5.000853, 5.001713, 5.00328, 5.005985, 5.010404, 5.017234, 
    5.027194, 5.040734, 5.058229, 5.079662, 5.104465, 5.131642, 5.158663, 
    5.182254, 5.198014, 5.203566, 5.197978, 5.182171, 5.158515, 5.131409, 
    5.104133, 5.079228, 5.057729, 5.040246, 5.026826, 5.017087, 5.010396, 
    5.006039, 5.00335, 5.001772, 5.000896, 5.000432, 5.000201, 5.000089, 
    5.000038, 5.000018, 5.00001, 5.000006, 5.000001, 5,
  // height(5,4, 0-49)
    5, 5, 5.000002, 5.000008, 5.000016, 5.000034, 5.000082, 5.000193, 
    5.000432, 5.000931, 5.001913, 5.003746, 5.006992, 5.012434, 5.021055, 
    5.033954, 5.052146, 5.075799, 5.105033, 5.139303, 5.177319, 5.217662, 
    5.25659, 5.289864, 5.311574, 5.319134, 5.311477, 5.289647, 5.256206, 
    5.217056, 5.176451, 5.13817, 5.103726, 5.074522, 5.051179, 5.033571, 
    5.021023, 5.012565, 5.007167, 5.003901, 5.002026, 5.001004, 5.000476, 
    5.000216, 5.000093, 5.00004, 5.000018, 5.00001, 5.000005, 5,
  // height(5,5, 0-49)
    5, 5.000001, 5.000006, 5.000015, 5.000033, 5.000081, 5.000193, 5.000442, 
    5.000971, 5.002039, 5.004083, 5.00779, 5.014157, 5.024488, 5.040304, 
    5.063102, 5.094024, 5.131987, 5.176251, 5.225178, 5.276432, 5.328592, 
    5.376917, 5.417064, 5.442416, 5.451099, 5.442188, 5.416547, 5.376002, 
    5.32715, 5.274362, 5.222458, 5.173093, 5.128881, 5.09165, 5.062176, 
    5.040218, 5.024799, 5.014578, 5.008171, 5.004367, 5.002228, 5.001084, 
    5.000504, 5.000224, 5.000095, 5.00004, 5.000018, 5.000009, 5.000004,
  // height(5,6, 0-49)
    5.000001, 5.000005, 5.000013, 5.000031, 5.000074, 5.000183, 5.00043, 
    5.000967, 5.002075, 5.004246, 5.008282, 5.015374, 5.02715, 5.045572, 
    5.072659, 5.110019, 5.15846, 5.213607, 5.273174, 5.334088, 5.393208, 
    5.450352, 5.500582, 5.540859, 5.565177, 5.573293, 5.564681, 5.539737, 
    5.498604, 5.447233, 5.388718, 5.328151, 5.266213, 5.206674, 5.153087, 
    5.107989, 5.072482, 5.046282, 5.028121, 5.016266, 5.008961, 5.004705, 
    5.002356, 5.001125, 5.000514, 5.000224, 5.000093, 5.000038, 5.000018, 
    5.000008,
  // height(5,7, 0-49)
    5.000004, 5.00001, 5.000028, 5.000067, 5.000166, 5.0004, 5.000918, 
    5.002015, 5.004214, 5.008401, 5.015932, 5.02872, 5.04916, 5.079797, 
    5.122718, 5.178854, 5.248075, 5.319426, 5.389174, 5.453479, 5.509659, 
    5.560696, 5.602446, 5.634424, 5.65239, 5.658066, 5.651396, 5.632189, 
    5.598525, 5.554535, 5.500804, 5.441733, 5.375283, 5.305392, 5.237004, 
    5.174875, 5.122472, 5.081369, 5.051301, 5.030718, 5.017484, 5.009469, 
    5.004883, 5.002399, 5.001125, 5.000504, 5.000216, 5.000089, 5.000036, 
    5.000016,
  // height(5,8, 0-49)
    5.000009, 5.000022, 5.000058, 5.000145, 5.000354, 5.000831, 5.001863, 
    5.003988, 5.008126, 5.015749, 5.028997, 5.050632, 5.083705, 5.130813, 
    5.193053, 5.269456, 5.35902, 5.440007, 5.509358, 5.56441, 5.604834, 
    5.638444, 5.662354, 5.67907, 5.686673, 5.688493, 5.684813, 5.674917, 
    5.655134, 5.627209, 5.588828, 5.543271, 5.484299, 5.414421, 5.338465, 
    5.262632, 5.193025, 5.134175, 5.088205, 5.054886, 5.03237, 5.018123, 
    5.009644, 5.004883, 5.002356, 5.001084, 5.000476, 5.000201, 5.000082, 
    5.000034,
  // height(5,9, 0-49)
    5.000019, 5.000048, 5.00012, 5.000298, 5.000716, 5.001643, 5.003593, 
    5.007489, 5.014842, 5.027926, 5.049793, 5.083932, 5.133445, 5.199761, 
    5.281408, 5.374544, 5.47942, 5.558947, 5.615193, 5.648915, 5.663444, 
    5.671911, 5.672351, 5.669973, 5.665254, 5.662431, 5.661954, 5.662679, 
    5.659845, 5.652761, 5.636622, 5.613993, 5.574114, 5.516903, 5.445178, 
    5.364569, 5.282547, 5.20661, 5.142382, 5.092508, 5.056751, 5.032938, 
    5.018123, 5.009469, 5.004705, 5.002228, 5.001004, 5.000433, 5.00018, 
    5.000075,
  // height(5,10, 0-49)
    5.000036, 5.000093, 5.000239, 5.000585, 5.001373, 5.003076, 5.006561, 
    5.013308, 5.02562, 5.046711, 5.08042, 5.130344, 5.198357, 5.283011, 
    5.378876, 5.479668, 5.591911, 5.658225, 5.691349, 5.696425, 5.68037, 
    5.66087, 5.636159, 5.613672, 5.596256, 5.58842, 5.590661, 5.601462, 
    5.615591, 5.630049, 5.638243, 5.642887, 5.629557, 5.59555, 5.540604, 
    5.467718, 5.383308, 5.296116, 5.215004, 5.146606, 5.093976, 5.056751, 
    5.03237, 5.017484, 5.008961, 5.004367, 5.002027, 5.000896, 5.000381, 
    5.000162,
  // height(5,11, 0-49)
    5.000071, 5.000181, 5.000453, 5.001088, 5.002494, 5.005449, 5.011323, 
    5.022336, 5.041712, 5.073508, 5.121789, 5.189017, 5.274099, 5.371275, 
    5.471056, 5.567159, 5.679311, 5.724144, 5.729917, 5.705225, 5.659316, 
    5.612999, 5.564149, 5.522204, 5.492456, 5.479336, 5.483345, 5.502607, 
    5.531834, 5.56584, 5.596796, 5.628322, 5.64375, 5.638568, 5.609673, 
    5.556548, 5.482425, 5.39456, 5.302978, 5.217842, 5.146606, 5.092508, 
    5.054886, 5.030718, 5.016266, 5.008171, 5.003901, 5.001774, 5.000774, 
    5.000335,
  // height(5,12, 0-49)
    5.000131, 5.00033, 5.000812, 5.001908, 5.004274, 5.00911, 5.018438, 
    5.035336, 5.0639, 5.108568, 5.172517, 5.255433, 5.351807, 5.45142, 
    5.54234, 5.622025, 5.729712, 5.750149, 5.730207, 5.67971, 5.608513, 
    5.538956, 5.468381, 5.40834, 5.366759, 5.347938, 5.352461, 5.37809, 
    5.419709, 5.470071, 5.520361, 5.575464, 5.617815, 5.642097, 5.643387, 
    5.618141, 5.565696, 5.48967, 5.398307, 5.302978, 5.215004, 5.142382, 
    5.088205, 5.051301, 5.028121, 5.014579, 5.007169, 5.003353, 5.001502, 
    5.000663,
  // height(5,13, 0-49)
    5.000229, 5.000569, 5.001369, 5.00315, 5.006894, 5.014339, 5.02826, 
    5.052577, 5.091915, 5.1502, 5.228284, 5.321659, 5.420121, 5.510469, 
    5.580884, 5.636158, 5.738116, 5.735927, 5.695858, 5.626519, 5.536742, 
    5.448798, 5.359662, 5.283228, 5.230228, 5.205044, 5.208557, 5.238231, 
    5.289241, 5.352497, 5.418259, 5.492509, 5.55786, 5.608896, 5.639956, 
    5.645646, 5.622089, 5.568675, 5.48967, 5.39456, 5.296116, 5.20661, 
    5.134175, 5.081369, 5.046282, 5.0248, 5.012568, 5.006046, 5.00278, 
    5.001256,
  // height(5,14, 0-49)
    5.000374, 5.000917, 5.002163, 5.004873, 5.010436, 5.021191, 5.040668, 
    5.073408, 5.123923, 5.194474, 5.282308, 5.378265, 5.468612, 5.539557, 
    5.581494, 5.609149, 5.704862, 5.684734, 5.631863, 5.551764, 5.45104, 
    5.350298, 5.246478, 5.15581, 5.091814, 5.059381, 5.060057, 5.091223, 
    5.148467, 5.22124, 5.298869, 5.387869, 5.471773, 5.545377, 5.60301, 
    5.638582, 5.646293, 5.622088, 5.565695, 5.482424, 5.383307, 5.282547, 
    5.193025, 5.122472, 5.072483, 5.040219, 5.021027, 5.010407, 5.004912, 
    5.002266,
  // height(5,15, 0-49)
    5.000567, 5.001374, 5.003187, 5.00704, 5.014763, 5.029299, 5.054786, 
    5.09597, 5.156433, 5.235746, 5.326997, 5.417121, 5.49086, 5.535902, 
    5.545708, 5.546775, 5.632914, 5.60088, 5.542744, 5.459904, 5.356049, 
    5.248635, 5.134977, 5.033073, 4.95883, 4.918158, 4.913803, 4.943549, 
    5.003622, 5.082602, 5.168946, 5.268797, 5.367137, 5.458964, 5.538911, 
    5.600954, 5.638575, 5.645641, 5.618137, 5.556546, 5.467716, 5.364568, 
    5.262632, 5.174875, 5.10799, 5.062179, 5.033578, 5.017106, 5.008286, 
    5.003901,
  // height(5,16, 0-49)
    5.000793, 5.001904, 5.004345, 5.009432, 5.01941, 5.037717, 5.06884, 
    5.117216, 5.184804, 5.268004, 5.356136, 5.433732, 5.48586, 5.502688, 
    5.480472, 5.459173, 5.525829, 5.488203, 5.431913, 5.353796, 5.254422, 
    5.146871, 5.029435, 4.92056, 4.837578, 4.787774, 4.775797, 4.80067, 
    4.859735, 4.941498, 5.033751, 5.14112, 5.250391, 5.356567, 5.454606, 
    5.538887, 5.602984, 5.639937, 5.643376, 5.609665, 5.5406, 5.445177, 
    5.338465, 5.237003, 5.153089, 5.091654, 5.05119, 5.026856, 5.013346, 
    5.006411,
  // height(5,17, 0-49)
    5.001009, 5.002405, 5.005424, 5.01161, 5.023516, 5.044888, 5.080247, 
    5.133332, 5.204224, 5.28643, 5.36658, 5.428285, 5.457914, 5.448078, 
    5.397178, 5.359798, 5.38727, 5.349489, 5.301646, 5.235264, 5.147697, 
    5.046798, 4.932895, 4.822896, 4.733915, 4.674499, 4.651908, 4.667727, 
    4.721311, 4.802092, 4.897588, 5.009571, 5.126815, 5.244068, 5.35647, 
    5.458864, 5.5453, 5.608845, 5.642067, 5.638551, 5.595541, 5.5169, 
    5.414419, 5.305392, 5.206675, 5.128885, 5.074537, 5.040285, 5.020535, 
    5.010053,
  // height(5,18, 0-49)
    5.001149, 5.002726, 5.006095, 5.012916, 5.025878, 5.048788, 5.085967, 
    5.140407, 5.210714, 5.288495, 5.358942, 5.405567, 5.415976, 5.384698, 
    5.312162, 5.264491, 5.221843, 5.186554, 5.153127, 5.1055, 5.037116, 
    4.949855, 4.847899, 4.744311, 4.653742, 4.585035, 4.548517, 4.550172, 
    4.592954, 4.668444, 4.76445, 4.87837, 5.000965, 5.126472, 5.250022, 
    5.366846, 5.471569, 5.55773, 5.617738, 5.643708, 5.629535, 5.574101, 
    5.484294, 5.375281, 5.266214, 5.1731, 5.103745, 5.057774, 5.03019, 
    5.015046,
  // height(5,19, 0-49)
    5.001132, 5.00268, 5.005971, 5.012604, 5.025155, 5.04725, 5.082956, 
    5.134978, 5.201641, 5.274235, 5.337543, 5.374701, 5.373543, 5.330182, 
    5.248117, 5.187968, 5.03577, 5.00039, 4.986063, 4.964749, 4.923753, 
    4.857672, 4.777114, 4.68915, 4.603427, 4.527005, 4.473067, 4.454343, 
    4.479911, 4.545097, 4.638662, 4.751842, 4.87722, 5.008308, 5.14009, 
    5.268059, 5.38738, 5.492204, 5.575282, 5.62822, 5.642832, 5.613966, 
    5.543258, 5.441728, 5.32815, 5.222465, 5.138189, 5.079276, 5.042429, 
    5.021496,
  // height(5,20, 0-49)
    5.000885, 5.002056, 5.004517, 5.009397, 5.018436, 5.033949, 5.05833, 
    5.092862, 5.13604, 5.182454, 5.22361, 5.251111, 5.26051, 5.253445, 
    5.236856, 0, 4.882641, 4.890296, 4.897371, 4.893323, 4.87047, 4.819962, 
    4.758723, 4.686413, 4.605082, 4.517176, 4.437809, 4.388928, 4.388727, 
    4.437592, 4.525457, 4.634996, 4.760348, 4.894176, 5.031245, 5.167237, 
    5.297763, 5.417573, 5.519956, 5.596563, 5.638118, 5.636558, 5.588799, 
    5.500793, 5.388714, 5.274365, 5.176466, 5.104169, 5.057017, 5.029309,
  // height(5,21, 0-49)
    5.000641, 5.001482, 5.003266, 5.006831, 5.013499, 5.025104, 5.043731, 
    5.070997, 5.106867, 5.148563, 5.190476, 5.225755, 5.249031, 5.258772, 
    5.257997, 0, 4.74108, 4.76133, 4.784954, 4.801523, 4.801844, 4.771854, 
    4.732392, 4.676557, 4.600542, 4.503641, 4.402691, 4.328095, 4.306149, 
    4.341571, 4.42612, 4.532413, 4.657756, 4.794104, 4.93592, 5.078889, 
    5.218863, 5.351027, 5.469194, 5.565336, 5.629769, 5.652613, 5.627135, 
    5.554501, 5.447219, 5.327146, 5.217059, 5.131421, 5.073335, 5.038131,
  // height(5,22, 0-49)
    5.000444, 5.00103, 5.002293, 5.004852, 5.009718, 5.018359, 5.0326, 
    5.054197, 5.084013, 5.121048, 5.161894, 5.201262, 5.233709, 5.255754, 
    5.267343, 0, 4.627163, 4.653697, 4.689208, 4.723159, 4.745467, 4.737381, 
    4.725026, 4.694858, 4.635277, 4.538174, 4.417841, 4.312981, 4.261384, 
    4.275565, 4.351222, 4.44836, 4.569024, 4.704297, 4.848145, 4.995989, 
    5.143591, 5.286217, 5.41789, 5.530775, 5.614996, 5.659525, 5.65497, 
    5.598444, 5.498568, 5.375984, 5.256189, 5.158487, 5.089858, 5.047126,
  // height(5,23, 0-49)
    5.000326, 5.000756, 5.0017, 5.003643, 5.007394, 5.014186, 5.025643, 
    5.043532, 5.069174, 5.102598, 5.141809, 5.182737, 5.220225, 5.249777, 
    5.26927, 0, 4.542715, 4.572813, 4.616893, 4.664588, 4.705509, 4.716725, 
    4.729808, 4.725214, 4.68426, 4.591591, 4.457345, 4.326142, 4.246144, 
    4.238336, 4.303779, 4.389193, 4.502711, 4.634574, 4.778222, 4.928749, 
    5.081713, 5.232281, 5.374473, 5.500473, 5.600245, 5.662012, 5.674566, 
    5.632014, 5.539653, 5.416502, 5.289604, 5.182093, 5.104459, 5.055098,
  // height(5,24, 0-49)
    5.000295, 5.00068, 5.00153, 5.00328, 5.006674, 5.012842, 5.023315, 
    5.039814, 5.063758, 5.095514, 5.133634, 5.174624, 5.213623, 5.245886, 
    5.268474, 0, 4.488168, 4.520331, 4.569875, 4.626774, 4.680708, 4.705749, 
    4.737486, 4.751808, 4.725004, 4.637198, 4.495549, 4.347715, 4.248083, 
    4.223984, 4.28151, 4.357102, 4.464386, 4.592849, 4.73542, 4.886861, 
    5.042512, 5.19742, 5.345583, 5.479222, 5.588269, 5.660618, 5.684098, 
    5.651032, 5.564503, 5.442098, 5.311407, 5.19786, 5.114362, 5.060548,
  // height(5,25, 0-49)
    5.000359, 5.000815, 5.001808, 5.003817, 5.007643, 5.014476, 5.025854, 
    5.043424, 5.068394, 5.100799, 5.138853, 5.178908, 5.216267, 5.246636, 
    5.267615, 0, 4.464517, 4.497284, 4.548565, 4.608568, 4.667108, 4.6971, 
    4.73595, 4.757792, 4.737058, 4.652288, 4.509429, 4.356791, 4.250607, 
    4.22062, 4.27515, 4.34684, 4.451613, 4.57867, 4.72073, 4.872409, 
    5.028946, 5.185324, 5.335518, 5.471749, 5.583937, 5.659878, 5.6871, 
    5.657343, 5.572935, 5.450924, 5.319024, 5.203423, 5.117879, 5.062491,
  // height(5,26, 0-49)
    5.000526, 5.001181, 5.002566, 5.005302, 5.010374, 5.01916, 5.033297, 
    5.054275, 5.082738, 5.117734, 5.156352, 5.194211, 5.226768, 5.250868, 
    5.265858, 0, 4.47485, 4.506453, 4.555189, 4.611245, 4.664432, 4.688535, 
    4.720223, 4.735377, 4.710451, 4.625587, 4.487513, 4.343034, 4.245784, 
    4.222999, 4.281123, 4.356955, 4.46433, 4.592826, 4.735413, 4.886859, 
    5.042512, 5.19742, 5.345583, 5.479222, 5.588269, 5.660618, 5.684098, 
    5.651031, 5.564503, 5.442098, 5.311407, 5.19786, 5.114362, 5.060548,
  // height(5,27, 0-49)
    5.000805, 5.001794, 5.003833, 5.007775, 5.014898, 5.026875, 5.045452, 
    5.071789, 5.105519, 5.144054, 5.182762, 5.21631, 5.240609, 5.254356, 
    5.259472, 0, 4.523546, 4.551486, 4.592946, 4.637959, 4.676403, 4.684864, 
    4.697034, 4.693454, 4.655822, 4.568797, 4.441556, 4.316923, 4.241585, 
    4.236356, 4.302987, 4.388885, 4.502593, 4.634529, 4.778204, 4.928742, 
    5.081711, 5.232281, 5.374472, 5.500473, 5.600244, 5.662012, 5.674566, 
    5.632014, 5.539653, 5.416502, 5.289604, 5.182093, 5.104459, 5.055098,
  // height(5,28, 0-49)
    5.001189, 5.002643, 5.005589, 5.011191, 5.021119, 5.037401, 5.061837, 
    5.094956, 5.134828, 5.176611, 5.213614, 5.239749, 5.252041, 5.251792, 
    5.243953, 0, 4.61626, 4.63638, 4.665257, 4.692745, 4.709127, 4.695071, 
    4.679724, 4.649843, 4.594497, 4.505446, 4.395233, 4.299756, 4.254767, 
    4.27263, 4.350018, 4.447882, 4.568835, 4.704223, 4.848115, 4.995977, 
    5.143586, 5.286216, 5.417889, 5.530774, 5.614996, 5.659525, 5.65497, 
    5.598445, 5.498568, 5.375984, 5.256189, 5.158487, 5.089858, 5.047126,
  // height(5,29, 0-49)
    5.001638, 5.003657, 5.007708, 5.01534, 5.02871, 5.05025, 5.081713, 
    5.122604, 5.168763, 5.212454, 5.244812, 5.259601, 5.255975, 5.238696, 
    5.215979, 0, 4.757369, 4.761571, 4.770969, 4.774717, 4.763777, 4.723468, 
    4.678093, 4.621346, 4.550265, 4.463518, 4.37518, 4.311992, 4.297986, 
    4.337866, 4.424553, 4.531772, 4.657499, 4.794, 4.935878, 5.078872, 
    5.218856, 5.351024, 5.469192, 5.565335, 5.629769, 5.652613, 5.627135, 
    5.554501, 5.447219, 5.327146, 5.217059, 5.131421, 5.073335, 5.038131,
  // height(5,30, 0-49)
    5.002085, 5.004748, 5.010147, 5.020489, 5.03899, 5.069524, 5.115261, 
    5.176115, 5.24598, 5.31214, 5.358694, 5.372374, 5.346906, 5.283526, 
    5.188242, 5.105539, 4.913468, 4.864236, 4.846265, 4.829531, 4.79874, 
    4.743309, 4.680916, 4.612876, 4.541994, 4.469274, 4.40619, 4.370837, 
    4.379624, 4.433442, 4.523681, 4.634262, 4.760047, 4.894053, 5.031196, 
    5.167217, 5.297757, 5.417571, 5.519956, 5.596563, 5.638118, 5.636558, 
    5.588799, 5.500793, 5.388714, 5.274365, 5.176466, 5.104169, 5.057017, 
    5.029309,
  // height(5,31, 0-49)
    5.002143, 5.004889, 5.010488, 5.021266, 5.040632, 5.072723, 5.12099, 
    5.185519, 5.260214, 5.332315, 5.385979, 5.407974, 5.391459, 5.335916, 
    5.244624, 5.177097, 5.096328, 5.048657, 5.011378, 4.966193, 4.904812, 
    4.824902, 4.735695, 4.645541, 4.563855, 4.495916, 4.451912, 4.441776, 
    4.473276, 4.541901, 4.637214, 4.751214, 4.876952, 5.008195, 5.140043, 
    5.268041, 5.387373, 5.492201, 5.575282, 5.62822, 5.642832, 5.613966, 
    5.543258, 5.441728, 5.328151, 5.222465, 5.138189, 5.079276, 5.042429, 
    5.021496,
  // height(5,32, 0-49)
    5.001922, 5.004405, 5.009535, 5.019537, 5.037773, 5.068523, 5.115789, 
    5.180799, 5.258986, 5.338832, 5.40467, 5.442245, 5.443079, 5.405014, 
    5.329818, 5.271312, 5.264867, 5.214771, 5.161846, 5.095674, 5.012313, 
    4.915738, 4.80939, 4.706865, 4.621886, 4.561248, 4.53286, 4.540988, 
    4.588072, 4.666042, 4.76333, 4.877868, 5.000745, 5.126377, 5.249983, 
    5.366829, 5.471562, 5.557727, 5.617737, 5.643708, 5.629536, 5.574101, 
    5.484294, 5.375281, 5.266214, 5.1731, 5.103745, 5.057774, 5.03019, 
    5.015046,
  // height(5,33, 0-49)
    5.00155, 5.003578, 5.007845, 5.01632, 5.032094, 5.059364, 5.102615, 
    5.16453, 5.242973, 5.328912, 5.40777, 5.464293, 5.487687, 5.473557, 
    5.422353, 5.376557, 5.412996, 5.361646, 5.298301, 5.217968, 5.119894, 
    5.013451, 4.898541, 4.791826, 4.709034, 4.656785, 4.640617, 4.661203, 
    4.717844, 4.800365, 4.89677, 5.009197, 5.126649, 5.243997, 5.35644, 
    5.458851, 5.545294, 5.608843, 5.642066, 5.638551, 5.595541, 5.5169, 
    5.414419, 5.305392, 5.206675, 5.128885, 5.074537, 5.040285, 5.020535, 
    5.010053,
  // height(5,34, 0-49)
    5.001143, 5.002663, 5.005934, 5.012573, 5.025232, 5.04776, 5.084791, 
    5.14025, 5.21467, 5.302464, 5.391526, 5.466604, 5.514605, 5.528172, 
    5.505728, 5.478414, 5.53635, 5.487955, 5.419987, 5.331903, 5.225847, 
    5.115927, 5, 4.895658, 4.818719, 4.774924, 4.767848, 4.796153, 4.857343, 
    4.940302, 5.033179, 5.140856, 5.250273, 5.356515, 5.454584, 5.538877, 
    5.60298, 5.639935, 5.643376, 5.609665, 5.5406, 5.445177, 5.338465, 
    5.237003, 5.153089, 5.091654, 5.05119, 5.026856, 5.013346, 5.006411,
  // height(5,35, 0-49)
    5.000779, 5.001836, 5.004165, 5.009008, 5.018488, 5.035882, 5.065555, 
    5.112102, 5.1783, 5.262308, 5.355819, 5.445318, 5.51646, 5.558745, 
    5.567586, 5.563785, 5.631766, 5.591699, 5.525231, 5.435889, 5.328604, 
    5.221323, 5.110783, 5.013813, 4.944966, 4.909076, 4.90834, 4.940494, 
    5.002017, 5.0818, 5.168562, 5.26862, 5.367057, 5.45893, 5.538898, 
    5.600948, 5.638573, 5.645639, 5.618137, 5.556546, 5.467717, 5.364568, 
    5.262632, 5.174875, 5.10799, 5.062179, 5.033578, 5.017106, 5.008286, 
    5.003901,
  // height(5,36, 0-49)
    5.000493, 5.00118, 5.002732, 5.006036, 5.012685, 5.025267, 5.047535, 
    5.084073, 5.139023, 5.213765, 5.304395, 5.400975, 5.489923, 5.558537, 
    5.598734, 5.621789, 5.695973, 5.669862, 5.611474, 5.527821, 5.42626, 
    5.327377, 5.227425, 5.141449, 5.081936, 5.053137, 5.056394, 5.089209, 
    5.147419, 5.22072, 5.298621, 5.387753, 5.471721, 5.545353, 5.603, 
    5.638578, 5.646291, 5.622087, 5.565695, 5.482424, 5.383308, 5.282547, 
    5.193025, 5.122472, 5.072483, 5.040219, 5.021027, 5.010407, 5.004912, 
    5.002266,
  // height(5,37, 0-49)
    5.000292, 5.00071, 5.00168, 5.003798, 5.008177, 5.016725, 5.032395, 
    5.059221, 5.101714, 5.163327, 5.244109, 5.338745, 5.436703, 5.525202, 
    5.5934, 5.644053, 5.725108, 5.718331, 5.675017, 5.604451, 5.51567, 
    5.430519, 5.345299, 5.272915, 5.223416, 5.200871, 5.206166, 5.236938, 
    5.288577, 5.352169, 5.418102, 5.492436, 5.557827, 5.608882, 5.639949, 
    5.645644, 5.622088, 5.568674, 5.489669, 5.39456, 5.296116, 5.20661, 
    5.134175, 5.081369, 5.046282, 5.0248, 5.012568, 5.006046, 5.00278, 
    5.001256,
  // height(5,38, 0-49)
    5.000163, 5.000402, 5.000972, 5.002252, 5.004967, 5.01043, 5.02079, 
    5.039236, 5.069869, 5.116913, 5.18307, 5.267374, 5.363808, 5.462077, 
    5.550688, 5.62586, 5.715589, 5.73241, 5.710911, 5.660795, 5.591628, 
    5.525109, 5.458025, 5.401213, 5.362216, 5.345235, 5.350946, 5.377285, 
    5.419301, 5.469871, 5.520268, 5.57542, 5.617796, 5.642089, 5.643384, 
    5.61814, 5.565695, 5.489669, 5.398307, 5.302978, 5.215004, 5.142382, 
    5.088205, 5.051301, 5.028121, 5.014579, 5.007169, 5.003353, 5.001502, 
    5.000663,
  // height(5,39, 0-49)
    5.000086, 5.000216, 5.000532, 5.00126, 5.002849, 5.006141, 5.012588, 
    5.024494, 5.045127, 5.078468, 5.128332, 5.196746, 5.282134, 5.37842, 
    5.476128, 5.568144, 5.666311, 5.708275, 5.713571, 5.690119, 5.646567, 
    5.603043, 5.557014, 5.517471, 5.489532, 5.477641, 5.482416, 5.502121, 
    5.53159, 5.565724, 5.596741, 5.628298, 5.64374, 5.638564, 5.60967, 
    5.556547, 5.482424, 5.39456, 5.302978, 5.217841, 5.146606, 5.092508, 
    5.054886, 5.030718, 5.016266, 5.008171, 5.003901, 5.001774, 5.000774, 
    5.000335,
  // height(5,40, 0-49)
    5.000043, 5.00011, 5.000275, 5.000667, 5.001546, 5.00342, 5.007205, 
    5.014437, 5.02746, 5.049472, 5.084197, 5.134979, 5.203325, 5.287435, 
    5.381662, 5.479102, 5.581413, 5.64549, 5.67866, 5.685199, 5.671315, 
    5.65408, 5.631466, 5.610655, 5.594442, 5.587394, 5.59011, 5.601179, 
    5.615451, 5.629982, 5.638213, 5.642873, 5.629552, 5.595548, 5.540603, 
    5.467717, 5.383308, 5.296116, 5.215004, 5.146606, 5.093976, 5.056751, 
    5.03237, 5.017484, 5.008961, 5.004367, 5.002027, 5.000896, 5.000381, 
    5.000162,
  // height(5,41, 0-49)
    5.000021, 5.000053, 5.000136, 5.000334, 5.000796, 5.001806, 5.003906, 
    5.008049, 5.015777, 5.029372, 5.051832, 5.086515, 5.136288, 5.202295, 
    5.282791, 5.373473, 5.471925, 5.54978, 5.606205, 5.641187, 5.657415, 
    5.667536, 5.669413, 5.668134, 5.664176, 5.661833, 5.66164, 5.662522, 
    5.65977, 5.652724, 5.636606, 5.613986, 5.57411, 5.516902, 5.445177, 
    5.364569, 5.282547, 5.20661, 5.142382, 5.092508, 5.056751, 5.032938, 
    5.018123, 5.009469, 5.004705, 5.002228, 5.001004, 5.000433, 5.00018, 
    5.000075,
  // height(5,42, 0-49)
    5.00001, 5.000026, 5.000064, 5.00016, 5.000389, 5.000905, 5.002008, 
    5.004252, 5.008577, 5.016464, 5.030032, 5.051978, 5.08522, 5.132163, 
    5.193682, 5.268489, 5.354282, 5.43411, 5.503586, 5.559516, 5.601096, 
    5.635793, 5.660614, 5.678005, 5.686062, 5.688162, 5.684644, 5.674834, 
    5.655095, 5.62719, 5.588821, 5.543266, 5.484297, 5.41442, 5.338465, 
    5.262631, 5.193025, 5.134175, 5.088205, 5.054886, 5.03237, 5.018123, 
    5.009644, 5.004883, 5.002356, 5.001084, 5.000476, 5.000201, 5.000082, 
    5.000034,
  // height(5,43, 0-49)
    5.000005, 5.000013, 5.00003, 5.000073, 5.000181, 5.000431, 5.000981, 
    5.002132, 5.00442, 5.008735, 5.016428, 5.029381, 5.049916, 5.080473, 
    5.122991, 5.178202, 5.245416, 5.316042, 5.385835, 5.450653, 5.507519, 
    5.559199, 5.60148, 5.633844, 5.652066, 5.657897, 5.651314, 5.632151, 
    5.598507, 5.554525, 5.500799, 5.441729, 5.37528, 5.30539, 5.237002, 
    5.174874, 5.122472, 5.081368, 5.051301, 5.030718, 5.017484, 5.009469, 
    5.004883, 5.002399, 5.001125, 5.000504, 5.000216, 5.000089, 5.000036, 
    5.000016,
  // height(5,44, 0-49)
    5.000001, 5.000006, 5.000015, 5.000033, 5.000081, 5.000196, 5.000456, 
    5.001016, 5.002163, 5.004395, 5.008506, 5.01568, 5.027507, 5.045893, 
    5.072774, 5.109653, 5.157123, 5.211867, 5.271431, 5.332604, 5.392085, 
    5.449572, 5.500086, 5.540573, 5.56503, 5.573226, 5.564657, 5.539729, 
    5.498598, 5.447226, 5.38871, 5.328142, 5.266205, 5.206667, 5.153083, 
    5.107986, 5.07248, 5.046281, 5.028121, 5.016266, 5.008961, 5.004705, 
    5.002356, 5.001125, 5.000514, 5.000224, 5.000093, 5.000038, 5.000018, 
    5.000008,
  // height(5,45, 0-49)
    5, 5.000002, 5.000007, 5.000016, 5.000035, 5.000085, 5.000203, 5.000461, 
    5.001007, 5.002101, 5.004179, 5.007924, 5.014315, 5.024631, 5.040349, 
    5.062917, 5.093406, 5.131166, 5.175416, 5.224458, 5.275883, 5.328215, 
    5.376691, 5.416956, 5.442389, 5.451115, 5.442218, 5.416569, 5.376009, 
    5.327141, 5.274342, 5.222435, 5.173072, 5.128863, 5.091638, 5.062168, 
    5.040212, 5.024796, 5.014577, 5.00817, 5.004367, 5.002228, 5.001084, 
    5.000504, 5.000224, 5.000095, 5.00004, 5.000018, 5.000009, 5.000004,
  // height(5,46, 0-49)
    5, 5, 5.000003, 5.000008, 5.000017, 5.000037, 5.000086, 5.0002, 5.000446, 
    5.000955, 5.001951, 5.0038, 5.007055, 5.012488, 5.021063, 5.033856, 
    5.051858, 5.075415, 5.104631, 5.138946, 5.177042, 5.217485, 5.256517, 
    5.289888, 5.311668, 5.319259, 5.311596, 5.289727, 5.256232, 5.217037, 
    5.176403, 5.138111, 5.10367, 5.074477, 5.051146, 5.033548, 5.021009, 
    5.012557, 5.007162, 5.003898, 5.002025, 5.001004, 5.000476, 5.000216, 
    5.000093, 5.00004, 5.000018, 5.00001, 5.000005, 5,
  // height(5,47, 0-49)
    5, 5, 5, 5.000004, 5.00001, 5.000017, 5.000035, 5.000082, 5.000188, 
    5.000413, 5.000865, 5.001729, 5.003295, 5.005988, 5.010376, 5.017145, 
    5.027009, 5.040486, 5.057955, 5.079401, 5.10426, 5.131539, 5.158699, 
    5.182441, 5.198313, 5.203908, 5.198285, 5.182379, 5.15859, 5.131369, 
    5.104017, 5.079085, 5.057591, 5.040131, 5.026741, 5.017027, 5.010357, 
    5.006016, 5.003337, 5.001766, 5.000893, 5.000431, 5.000199, 5.000088, 
    5.000038, 5.000018, 5.00001, 5.000006, 5.000001, 5,
  // height(5,48, 0-49)
    5, 5, 5, 5, 5.000005, 5.000009, 5.000016, 5.000033, 5.000074, 5.000168, 
    5.00036, 5.000737, 5.001443, 5.002692, 5.004791, 5.008132, 5.013163, 
    5.020295, 5.029888, 5.0421, 5.056754, 5.073282, 5.09015, 5.105158, 
    5.115366, 5.118993, 5.115357, 5.105136, 5.090113, 5.073223, 5.056668, 
    5.041988, 5.029758, 5.020169, 5.013067, 5.00809, 5.004785, 5.002703, 
    5.001458, 5.00075, 5.000369, 5.000174, 5.000078, 5.000034, 5.000016, 
    5.000009, 5.000005, 5.000001, 5, 5,
  // height(5,49, 0-49)
    5, 5, 5, 5, 5, 5.000002, 5.000004, 5.00001, 5.000021, 5.000049, 5.00011, 
    5.000237, 5.000488, 5.000957, 5.001791, 5.003193, 5.005428, 5.008776, 
    5.013537, 5.019944, 5.02806, 5.037715, 5.048037, 5.057581, 5.064183, 
    5.06655, 5.064181, 5.057576, 5.048025, 5.037696, 5.028031, 5.019907, 
    5.013492, 5.008731, 5.005393, 5.003181, 5.001791, 5.000962, 5.000493, 
    5.000242, 5.000113, 5.000051, 5.000022, 5.00001, 5.000005, 5.000002, 5, 
    5, 5, 5,
  // height(6,0, 0-49)
    5.000001, 5.000006, 5.00001, 5.000018, 5.000034, 5.000072, 5.000154, 
    5.000316, 5.000631, 5.001208, 5.002222, 5.003925, 5.006657, 5.010836, 
    5.01693, 5.025394, 5.036568, 5.050474, 5.066961, 5.08557, 5.105506, 
    5.125745, 5.144631, 5.160282, 5.170508, 5.174044, 5.170405, 5.160065, 
    5.144283, 5.12525, 5.104868, 5.084815, 5.066161, 5.049734, 5.036002, 
    5.025083, 5.016811, 5.010836, 5.006715, 5.003999, 5.002289, 5.00126, 
    5.000666, 5.00034, 5.000166, 5.000079, 5.000038, 5.000019, 5.000011, 
    5.000007,
  // height(6,1, 0-49)
    5.000005, 5.00001, 5.000018, 5.000033, 5.00007, 5.000151, 5.00032, 
    5.000653, 5.001278, 5.002406, 5.004348, 5.007544, 5.012561, 5.020073, 
    5.030783, 5.045307, 5.064008, 5.086517, 5.11232, 5.140503, 5.169809, 
    5.198979, 5.225753, 5.247741, 5.261885, 5.266718, 5.261647, 5.247239, 
    5.224946, 5.197832, 5.168324, 5.13874, 5.110439, 5.084771, 5.062673, 
    5.044592, 5.030516, 5.020079, 5.012699, 5.007718, 5.004508, 5.002532, 
    5.001365, 5.000708, 5.000353, 5.00017, 5.00008, 5.000038, 5.000021, 
    5.000012,
  // height(6,2, 0-49)
    5.000009, 5.000016, 5.000031, 5.000069, 5.000152, 5.000327, 5.000679, 
    5.001356, 5.002598, 5.004784, 5.008452, 5.014331, 5.023312, 5.036367, 
    5.054408, 5.078065, 5.107471, 5.141197, 5.177971, 5.216177, 5.254053, 
    5.290477, 5.322897, 5.349, 5.365357, 5.37082, 5.364851, 5.347931, 
    5.321181, 5.288037, 5.250886, 5.212396, 5.173913, 5.137403, 5.104555, 
    5.076529, 5.053838, 5.036386, 5.023619, 5.014725, 5.008818, 5.005071, 
    5.002802, 5.001487, 5.000758, 5.000372, 5.000178, 5.000082, 5.000039, 
    5.000021,
  // height(6,3, 0-49)
    5.000015, 5.000031, 5.000066, 5.000148, 5.000325, 5.000685, 5.001394, 
    5.002722, 5.005103, 5.009176, 5.015826, 5.026171, 5.041471, 5.06295, 
    5.091514, 5.127439, 5.170224, 5.216258, 5.26322, 5.308789, 5.351055, 
    5.389846, 5.422889, 5.44876, 5.464318, 5.469281, 5.463325, 5.446671, 
    5.41954, 5.385091, 5.344875, 5.301375, 5.2552, 5.208684, 5.164347, 
    5.124405, 5.090402, 5.063021, 5.042137, 5.027025, 5.016627, 5.009819, 
    5.005565, 5.003028, 5.001583, 5.000794, 5.000385, 5.00018, 5.000083, 
    5.00004,
  // height(6,4, 0-49)
    5.000029, 5.000062, 5.00014, 5.00031, 5.000668, 5.001381, 5.002748, 
    5.005244, 5.009598, 5.016839, 5.0283, 5.045533, 5.070081, 5.103135, 
    5.145094, 5.195261, 5.252154, 5.308517, 5.361249, 5.407907, 5.447248, 
    5.481152, 5.508186, 5.528504, 5.5398, 5.542978, 5.537997, 5.524723, 
    5.502158, 5.472632, 5.436204, 5.394633, 5.346801, 5.294731, 5.241333, 
    5.189841, 5.143176, 5.103406, 5.07149, 5.047315, 5.029989, 5.018214, 
    5.010605, 5.005923, 5.003174, 5.001634, 5.000808, 5.000386, 5.00018, 
    5.000086,
  // height(6,5, 0-49)
    5.000058, 5.000128, 5.000286, 5.000626, 5.001318, 5.002669, 5.005185, 
    5.009661, 5.017243, 5.029462, 5.048134, 5.075124, 5.1119, 5.158987, 
    5.215483, 5.279093, 5.347617, 5.408614, 5.459496, 5.498811, 5.526948, 
    5.548717, 5.563705, 5.573915, 5.578139, 5.578449, 5.57507, 5.567517, 
    5.553593, 5.534558, 5.508757, 5.477044, 5.435779, 5.385819, 5.329535, 
    5.270462, 5.212655, 5.159855, 5.114769, 5.078687, 5.051541, 5.032279, 
    5.019346, 5.011106, 5.006111, 5.003226, 5.001635, 5.000797, 5.000378, 
    5.000181,
  // height(6,6, 0-49)
    5.000115, 5.000255, 5.000564, 5.001209, 5.002492, 5.00493, 5.009352, 
    5.016989, 5.029522, 5.049008, 5.077607, 5.11707, 5.168053, 5.229499, 
    5.298431, 5.370821, 5.445284, 5.502716, 5.543248, 5.567499, 5.578008, 
    5.582731, 5.581964, 5.579405, 5.574989, 5.571723, 5.570034, 5.569163, 
    5.56598, 5.56068, 5.55012, 5.534544, 5.507586, 5.468422, 5.417926, 
    5.358761, 5.295095, 5.231841, 5.173631, 5.123855, 5.084163, 5.05453, 
    5.033725, 5.019936, 5.011277, 5.006112, 5.003177, 5.001587, 5.000769, 
    5.000376,
  // height(6,7, 0-49)
    5.000226, 5.000491, 5.001064, 5.002233, 5.004501, 5.008698, 5.016093, 
    5.028466, 5.048059, 5.0773, 5.118228, 5.171681, 5.236503, 5.309232, 
    5.384604, 5.457738, 5.530963, 5.576744, 5.600434, 5.605077, 5.595113, 
    5.581197, 5.563703, 5.547695, 5.534246, 5.527015, 5.526596, 5.532055, 
    5.539679, 5.548707, 5.554925, 5.558561, 5.5509, 5.529508, 5.493343, 
    5.443217, 5.382048, 5.31462, 5.246725, 5.183888, 5.130181, 5.087585, 
    5.056075, 5.034219, 5.019936, 5.011107, 5.005926, 5.003036, 5.001507, 
    5.000752,
  // height(6,8, 0-49)
    5.000422, 5.000904, 5.001921, 5.003942, 5.007765, 5.014642, 5.026388, 
    5.045363, 5.074217, 5.115291, 5.169679, 5.236262, 5.311226, 5.388562, 
    5.461514, 5.526134, 5.591987, 5.620574, 5.624623, 5.609064, 5.579417, 
    5.548193, 5.515173, 5.486481, 5.46438, 5.452968, 5.453032, 5.463569, 
    5.480635, 5.502585, 5.524538, 5.547294, 5.560452, 5.560471, 5.544627, 
    5.511597, 5.462111, 5.399347, 5.328711, 5.256863, 5.190205, 5.133425, 
    5.088749, 5.056075, 5.033725, 5.019349, 5.010611, 5.00558, 5.002838, 
    5.001445,
  // height(6,9, 0-49)
    5.000753, 5.001589, 5.003309, 5.006641, 5.012774, 5.023482, 5.041159, 
    5.068617, 5.108491, 5.162234, 5.228955, 5.304729, 5.382974, 5.456024, 
    5.5172, 5.565434, 5.620588, 5.629872, 5.615059, 5.581898, 5.535974, 
    5.490709, 5.444725, 5.404984, 5.375036, 5.359287, 5.358814, 5.372686, 
    5.397056, 5.429439, 5.464555, 5.504181, 5.536883, 5.558599, 5.565522, 
    5.554592, 5.52423, 5.475126, 5.410761, 5.337203, 5.261992, 5.192336, 
    5.133425, 5.087586, 5.054531, 5.032286, 5.018225, 5.009846, 5.005136, 
    5.00267,
  // height(6,10, 0-49)
    5.001282, 5.002665, 5.005434, 5.010663, 5.020015, 5.035825, 5.060974, 
    5.098361, 5.149876, 5.215099, 5.290311, 5.368649, 5.441668, 5.501667, 
    5.54359, 5.570598, 5.614685, 5.605386, 5.574833, 5.52846, 5.471034, 
    5.416002, 5.360381, 5.31177, 5.275041, 5.254829, 5.25267, 5.267902, 
    5.297109, 5.337039, 5.382149, 5.435371, 5.484737, 5.526087, 5.55515, 
    5.567821, 5.560739, 5.532126, 5.482728, 5.416425, 5.34004, 5.261992, 
    5.190205, 5.130182, 5.084167, 5.051551, 5.03001, 5.016677, 5.008926, 
    5.004739,
  // height(6,11, 0-49)
    5.002078, 5.004252, 5.008497, 5.016294, 5.029826, 5.051929, 5.085682, 
    5.133456, 5.195515, 5.268737, 5.346379, 5.41946, 5.479264, 5.519618, 
    5.53792, 5.542086, 5.576544, 5.550974, 5.508726, 5.454051, 5.390294, 
    5.330138, 5.268671, 5.213834, 5.171679, 5.146977, 5.141926, 5.156423, 
    5.187869, 5.232409, 5.284306, 5.34762, 5.410196, 5.467977, 5.516637, 
    5.551656, 5.568658, 5.564036, 5.535913, 5.485223, 5.416424, 5.337204, 
    5.256864, 5.183889, 5.12386, 5.078702, 5.04735, 5.027104, 5.014899, 
    5.008082,
  // height(6,12, 0-49)
    5.003199, 5.006451, 5.012627, 5.023664, 5.042225, 5.071439, 5.11411, 
    5.171338, 5.240982, 5.31694, 5.390095, 5.450813, 5.491652, 5.508848, 
    5.502183, 5.484329, 5.5107, 5.471681, 5.42171, 5.363332, 5.298191, 
    5.237552, 5.174379, 5.116498, 5.070714, 5.04173, 5.032598, 5.044168, 
    5.075143, 5.121388, 5.177038, 5.247113, 5.3195, 5.390254, 5.455167, 
    5.509714, 5.549153, 5.568865, 5.565066, 5.535909, 5.482724, 5.41076, 
    5.328711, 5.246729, 5.17364, 5.114793, 5.071546, 5.042262, 5.023884, 
    5.013244,
  // height(6,13, 0-49)
    5.004665, 5.00928, 5.017808, 5.032618, 5.056721, 5.093204, 5.144015, 
    5.208309, 5.2812, 5.354035, 5.416568, 5.459991, 5.479059, 5.472442, 
    5.441646, 5.404009, 5.422162, 5.372473, 5.318215, 5.260051, 5.197939, 
    5.141232, 5.080792, 5.023685, 4.976696, 4.944057, 4.92978, 4.936145, 
    4.963764, 5.008761, 5.065294, 5.139062, 5.21817, 5.298661, 5.376439, 
    5.447134, 5.506054, 5.548239, 5.568853, 5.564024, 5.532117, 5.475121, 
    5.399345, 5.314625, 5.231855, 5.159892, 5.10349, 5.063205, 5.036771, 
    5.020852,
  // height(6,14, 0-49)
    5.006432, 5.012634, 5.023786, 5.042606, 5.072232, 5.115298, 5.172375, 
    5.240322, 5.311727, 5.376356, 5.424157, 5.448103, 5.445302, 5.416306, 
    5.363493, 5.308928, 5.315402, 5.257618, 5.201933, 5.147207, 5.091923, 
    5.043219, 4.99018, 4.938323, 4.893336, 4.858306, 4.838092, 4.836915, 
    4.85803, 4.898629, 4.953203, 5.027792, 5.110849, 5.19822, 5.285783, 
    5.369319, 5.444354, 5.506011, 5.549108, 5.568622, 5.560715, 5.524216, 
    5.462107, 5.382053, 5.295115, 5.212708, 5.143295, 5.09066, 5.054367, 
    5.031552,
  // height(6,15, 0-49)
    5.008353, 5.01623, 5.03002, 5.052654, 5.087132, 5.135281, 5.196004, 
    5.263953, 5.329874, 5.383046, 5.414553, 5.419429, 5.396732, 5.348141, 
    5.276179, 5.207609, 5.194048, 5.130501, 5.075865, 5.027326, 4.982164, 
    4.945155, 4.904314, 4.862773, 4.823861, 4.788546, 4.762092, 4.751051, 
    4.762189, 4.794866, 4.844478, 4.917047, 5.001487, 5.09321, 5.187871, 
    5.281279, 5.369182, 5.446979, 5.509586, 5.551565, 5.567762, 5.554559, 
    5.511582, 5.443219, 5.358788, 5.270534, 5.190001, 5.124745, 5.077209, 
    5.045891,
  // height(6,16, 0-49)
    5.010181, 5.019599, 5.035693, 5.061436, 5.099479, 5.150658, 5.212265, 
    5.277219, 5.335279, 5.376088, 5.392232, 5.380555, 5.341426, 5.277007, 
    5.189547, 5.10928, 5.061175, 4.993652, 4.942364, 4.902635, 4.870674, 
    4.848741, 4.82494, 4.799216, 4.771264, 4.738774, 4.706534, 4.683522, 
    4.680879, 4.701571, 4.742841, 4.810379, 4.893664, 4.987398, 5.086774, 
    5.187449, 5.285298, 5.376024, 5.45486, 5.516427, 5.555016, 5.565443, 
    5.544588, 5.493336, 5.417953, 5.329622, 5.241532, 5.164762, 5.10537, 
    5.064186,
  // height(6,17, 0-49)
    5.011572, 5.022128, 5.039799, 5.067472, 5.107347, 5.159363, 5.219592, 
    5.279918, 5.329862, 5.35982, 5.363729, 5.339694, 5.288814, 5.213394, 
    5.115401, 5.023416, 4.91982, 4.848852, 4.803052, 4.775018, 4.75953, 
    4.755941, 4.754036, 4.749845, 4.738373, 4.712875, 4.676379, 4.639837, 
    4.619423, 4.623429, 4.652407, 4.711521, 4.790933, 4.884343, 4.986193, 
    5.091783, 5.19697, 5.297701, 5.389572, 5.46752, 5.525795, 5.558423, 
    5.560376, 5.529471, 5.46844, 5.385913, 5.294955, 5.209147, 5.138294, 
    5.086379,
  // height(6,18, 0-49)
    5.012167, 5.023161, 5.04132, 5.069361, 5.109135, 5.160046, 5.217618, 
    5.273468, 5.317338, 5.340284, 5.337028, 5.306277, 5.249497, 5.169226, 
    5.067511, 4.957667, 4.773083, 4.697157, 4.658534, 4.645606, 4.650552, 
    4.668773, 4.693651, 4.71667, 4.727506, 4.714119, 4.676271, 4.625728, 
    4.583766, 4.56583, 4.577911, 4.624625, 4.69708, 4.787639, 4.889681, 
    4.997922, 5.108042, 5.21612, 5.318082, 5.409255, 5.484136, 5.536518, 
    5.560242, 5.550798, 5.507571, 5.435857, 5.34702, 5.255654, 5.174771, 
    5.111942,
  // height(6,19, 0-49)
    5.011673, 5.022164, 5.039426, 5.06602, 5.103715, 5.152024, 5.206848, 
    5.260324, 5.302584, 5.324714, 5.321186, 5.290559, 5.234613, 5.15659, 
    5.058802, 4.913702, 4.622737, 4.538507, 4.507798, 4.513911, 4.544353, 
    4.588445, 4.64507, 4.700685, 4.73955, 4.744065, 4.709301, 4.645968, 
    4.579593, 4.53436, 4.524497, 4.554203, 4.616135, 4.700994, 4.800754, 
    4.909312, 5.022017, 5.134962, 5.244314, 5.345772, 5.434191, 5.503454, 
    5.546865, 5.558331, 5.534452, 5.477069, 5.394795, 5.301735, 5.213065, 
    5.139863,
  // height(6,20, 0-49)
    5.009789, 5.018234, 5.032057, 5.053111, 5.08257, 5.119898, 5.161999, 
    5.20331, 5.237241, 5.258398, 5.264359, 5.256173, 5.237612, 5.213781, 
    5.189564, 0, 4.351584, 4.34895, 4.370693, 4.414233, 4.476791, 4.54938, 
    4.639208, 4.728305, 4.795688, 4.818511, 4.786697, 4.708689, 4.613272, 
    4.53438, 4.497091, 4.504663, 4.552106, 4.628093, 4.722847, 4.829231, 
    4.942132, 5.057541, 5.171772, 5.280826, 5.379914, 5.463161, 5.523698, 
    5.554443, 5.54987, 5.508664, 5.436234, 5.345024, 5.251167, 5.168735,
  // height(6,21, 0-49)
    5.008009, 5.014865, 5.026288, 5.044007, 5.069425, 5.102808, 5.142482, 
    5.184568, 5.223716, 5.254673, 5.273949, 5.280734, 5.276828, 5.265878, 
    5.252289, 0, 4.170659, 4.190443, 4.237646, 4.309671, 4.403232, 4.505134, 
    4.625941, 4.743216, 4.833209, 4.872109, 4.84777, 4.765993, 4.654385, 
    4.551601, 4.492404, 4.478347, 4.510312, 4.576025, 4.664337, 4.767112, 
    4.878688, 4.994842, 5.111915, 5.226116, 5.33296, 5.426864, 5.501005, 
    5.547768, 5.560138, 5.534248, 5.47243, 5.384887, 5.287694, 5.197131,
  // height(6,22, 0-49)
    5.006531, 5.012131, 5.021671, 5.036806, 5.059116, 5.089477, 5.127281, 
    5.16994, 5.2131, 5.25171, 5.281518, 5.300305, 5.308352, 5.308174, 
    5.303796, 0, 4.030805, 4.065196, 4.131796, 4.227709, 4.348972, 4.477757, 
    4.627515, 4.771355, 4.883232, 4.939029, 4.924598, 4.842271, 4.716929, 
    4.590865, 4.509266, 4.470721, 4.484496, 4.53761, 4.617585, 4.715239, 
    4.824254, 4.940064, 5.058887, 5.17696, 5.289956, 5.392478, 5.47778, 
    5.537942, 5.564931, 5.552924, 5.501613, 5.41886, 5.320036, 5.22286,
  // height(6,23, 0-49)
    5.005608, 5.010423, 5.018781, 5.032283, 5.052613, 5.081013, 5.117546, 
    5.160475, 5.206153, 5.249742, 5.28655, 5.313443, 5.329684, 5.337036, 
    5.339309, 0, 3.936208, 3.979444, 4.05963, 4.173486, 4.31631, 4.465572, 
    4.636799, 4.799335, 4.926097, 4.994142, 4.988685, 4.909207, 4.776904, 
    4.635037, 4.536873, 4.476786, 4.473642, 4.514404, 4.585753, 4.677729, 
    4.783483, 4.898127, 5.017705, 5.138398, 5.255899, 5.364881, 5.458617, 
    5.528984, 5.567272, 5.566283, 5.52371, 5.445437, 5.345931, 5.243716,
  // height(6,24, 0-49)
    5.005395, 5.009989, 5.017999, 5.030992, 5.050661, 5.078343, 5.114321, 
    5.157181, 5.203599, 5.248916, 5.288375, 5.318546, 5.338296, 5.349046, 
    5.354481, 0, 3.885182, 3.932935, 4.020948, 4.145664, 4.301788, 4.463101, 
    4.646461, 4.818689, 4.952569, 5.026831, 5.027077, 4.951261, 4.817554, 
    4.668488, 4.561754, 4.487683, 4.472909, 4.504726, 4.569493, 4.656837, 
    4.759587, 4.872656, 4.991975, 5.113683, 5.233487, 5.346098, 5.444815, 
    5.521412, 5.566805, 5.572984, 5.536391, 5.461555, 5.362166, 5.257078,
  // height(6,25, 0-49)
    5.005977, 5.010957, 5.019516, 5.033198, 5.053604, 5.081876, 5.118042, 
    5.160445, 5.205666, 5.249183, 5.286569, 5.314772, 5.332943, 5.342594, 
    5.347287, 0, 3.875384, 3.92374, 4.013379, 4.140702, 4.30019, 4.464015, 
    4.64996, 4.823952, 4.9589, 5.034354, 5.036249, 4.962126, 4.829005, 
    4.67878, 4.570251, 4.491889, 4.473286, 4.501997, 4.564393, 4.650023, 
    4.75163, 4.864066, 4.983222, 5.105221, 5.225766, 5.339579, 5.439962, 
    5.518659, 5.566463, 5.575105, 5.5406, 5.46701, 5.367731, 5.261695,
  // height(6,26, 0-49)
    5.007358, 5.013331, 5.023318, 5.038845, 5.061301, 5.09135, 5.128307, 
    5.169772, 5.211891, 5.250265, 5.281169, 5.302535, 5.31439, 5.318717, 
    5.319005, 0, 3.907399, 3.952108, 4.036621, 4.157588, 4.309739, 4.466147, 
    4.645107, 4.813356, 4.943969, 5.016002, 5.015329, 4.94009, 4.808348, 
    4.662022, 4.557912, 4.485681, 4.471959, 4.5043, 4.569307, 4.656758, 
    4.759554, 4.872642, 4.991968, 5.113681, 5.233484, 5.346098, 5.444815, 
    5.521413, 5.566805, 5.572984, 5.53639, 5.461555, 5.362166, 5.257078,
  // height(6,27, 0-49)
    5.009464, 5.016989, 5.029191, 5.047569, 5.07317, 5.105905, 5.143998, 
    5.18394, 5.221245, 5.251712, 5.272612, 5.283283, 5.285047, 5.280668, 
    5.273688, 0, 3.984281, 4.020194, 4.092436, 4.198112, 4.332588, 4.472099, 
    4.634583, 4.789214, 4.909461, 4.973031, 4.965724, 4.887423, 4.759062, 
    4.622608, 4.529527, 4.472963, 4.471822, 4.513583, 4.585392, 4.677572, 
    4.783415, 4.898097, 5.017692, 5.138393, 5.255897, 5.36488, 5.458617, 
    5.528984, 5.567272, 5.566283, 5.52371, 5.445437, 5.345931, 5.243716,
  // height(6,28, 0-49)
    5.012121, 5.021662, 5.036722, 5.058746, 5.08832, 5.12436, 5.163691, 
    5.201473, 5.232535, 5.253003, 5.261386, 5.258695, 5.247797, 5.232471, 
    5.216447, 0, 4.109945, 4.130611, 4.183319, 4.265604, 4.37358, 4.487952, 
    4.624791, 4.757003, 4.859302, 4.908553, 4.891548, 4.811182, 4.691791, 
    4.573579, 4.499115, 4.465442, 4.481968, 4.536459, 4.617074, 4.715014, 
    4.824155, 4.940021, 5.058867, 5.176952, 5.289953, 5.392476, 5.477779, 
    5.537941, 5.564931, 5.552924, 5.501613, 5.41886, 5.320036, 5.22286,
  // height(6,29, 0-49)
    5.01504, 5.026921, 5.045306, 5.071594, 5.1058, 5.145628, 5.186234, 
    5.221255, 5.244844, 5.253647, 5.247667, 5.229831, 5.204763, 5.177385, 
    5.151611, 0, 4.284205, 4.28185, 4.307784, 4.359859, 4.434813, 4.518023, 
    4.622173, 4.724629, 4.802577, 4.8335, 4.806474, 4.727848, 4.624166, 
    4.531176, 4.480493, 4.472147, 4.507318, 4.574645, 4.663714, 4.766834, 
    4.878564, 4.994786, 5.11189, 5.226105, 5.332955, 5.426862, 5.501004, 
    5.547768, 5.560138, 5.534248, 5.47243, 5.384888, 5.287694, 5.197131,
  // height(6,30, 0-49)
    5.01805, 5.03292, 5.056044, 5.089447, 5.133391, 5.184988, 5.237677, 
    5.28241, 5.310273, 5.315083, 5.294526, 5.249707, 5.183735, 5.100007, 
    5.000019, 4.8457, 4.545903, 4.460265, 4.430046, 4.441324, 4.48198, 
    4.537408, 4.612211, 4.688424, 4.746189, 4.764202, 4.733611, 4.662929, 
    4.579001, 4.51218, 4.48446, 4.498162, 4.54897, 4.626636, 4.722182, 
    4.82893, 4.941996, 5.057481, 5.171744, 5.280814, 5.379909, 5.463158, 
    5.523697, 5.554443, 5.54987, 5.508664, 5.436234, 5.345024, 5.251167, 
    5.168735,
  // height(6,31, 0-49)
    5.019023, 5.03479, 5.059389, 5.094986, 5.141794, 5.196579, 5.252171, 
    5.298905, 5.32757, 5.332101, 5.310494, 5.263934, 5.195178, 5.107091, 
    5.00141, 4.883553, 4.684901, 4.605775, 4.566805, 4.557559, 4.570552, 
    4.598731, 4.639916, 4.681739, 4.709561, 4.707233, 4.671093, 4.611933, 
    4.553517, 4.517052, 4.514324, 4.54877, 4.613411, 4.699682, 4.800136, 
    4.909025, 5.021885, 5.134902, 5.244286, 5.345759, 5.434185, 5.503451, 
    5.546865, 5.558331, 5.534452, 5.477069, 5.394795, 5.301735, 5.213065, 
    5.139863,
  // height(6,32, 0-49)
    5.018395, 5.033809, 5.058214, 5.094069, 5.14203, 5.199332, 5.259036, 
    5.311258, 5.346146, 5.356833, 5.340679, 5.298523, 5.232965, 5.146788, 
    5.041823, 4.942011, 4.822749, 4.747123, 4.69965, 4.673524, 4.664025, 
    4.668962, 4.681037, 4.693107, 4.696065, 4.679071, 4.64244, 4.597218, 
    4.562731, 4.552108, 4.569833, 4.620241, 4.694829, 4.786526, 4.889145, 
    4.997667, 5.107924, 5.216065, 5.318056, 5.409244, 5.484132, 5.536515, 
    5.560241, 5.550798, 5.507571, 5.435857, 5.34702, 5.255654, 5.174771, 
    5.111942,
  // height(6,33, 0-49)
    5.016522, 5.030602, 5.0534, 5.087697, 5.134883, 5.193241, 5.256811, 
    5.316042, 5.360482, 5.382006, 5.376657, 5.344406, 5.287577, 5.209101, 
    5.111249, 5.021931, 4.958303, 4.88466, 4.830286, 4.790932, 4.763344, 
    4.748603, 4.736362, 4.723997, 4.707599, 4.681181, 4.647666, 4.616824, 
    4.603018, 4.612907, 4.64622, 4.708125, 4.789161, 4.883449, 4.985752, 
    5.091572, 5.196871, 5.297654, 5.389551, 5.46751, 5.525791, 5.558421, 
    5.560375, 5.529471, 5.46844, 5.385913, 5.294955, 5.209147, 5.138294, 
    5.086379,
  // height(6,34, 0-49)
    5.013892, 5.025993, 5.046119, 5.077284, 5.121665, 5.178928, 5.244718, 
    5.310551, 5.365828, 5.401097, 5.410602, 5.392849, 5.349452, 5.283387, 
    5.197491, 5.117618, 5.088926, 5.017687, 4.958633, 4.909221, 4.867121, 
    4.835982, 4.804241, 4.772992, 4.742702, 4.71132, 4.683036, 4.66551, 
    4.668421, 4.693704, 4.738229, 4.807829, 4.892317, 4.98671, 5.086431, 
    5.187284, 5.285219, 5.375988, 5.454842, 5.516418, 5.555013, 5.565441, 
    5.544586, 5.493335, 5.417953, 5.329622, 5.241532, 5.164762, 5.10537, 
    5.064186,
  // height(6,35, 0-49)
    5.010988, 5.020812, 5.037631, 5.064511, 5.10425, 5.157928, 5.223202, 
    5.293424, 5.358673, 5.408595, 5.435466, 5.43575, 5.409719, 5.359928, 
    5.289591, 5.220821, 5.212025, 5.144827, 5.083393, 5.026625, 4.973094, 
    4.928782, 4.882309, 4.837645, 4.798489, 4.765621, 4.743443, 4.737309, 
    4.752937, 4.789107, 4.841118, 4.915183, 5.000496, 5.092699, 5.187614, 
    5.281154, 5.369122, 5.446951, 5.509573, 5.55156, 5.56776, 5.554558, 
    5.511581, 5.443218, 5.358788, 5.270534, 5.190001, 5.124745, 5.077209, 
    5.045891,
  // height(6,36, 0-49)
    5.008206, 5.015754, 5.029075, 5.051062, 5.084832, 5.132618, 5.194133, 
    5.265147, 5.33742, 5.400627, 5.445424, 5.465913, 5.46032, 5.430084, 
    5.378282, 5.323157, 5.325123, 5.264044, 5.202501, 5.140908, 5.078958, 
    5.024843, 4.968314, 4.915356, 4.871645, 4.839771, 4.823688, 4.826664, 
    4.851294, 4.894493, 4.950805, 5.026462, 5.110141, 5.197854, 5.285599, 
    5.369229, 5.444311, 5.505991, 5.549098, 5.568619, 5.560713, 5.524215, 
    5.462106, 5.382053, 5.295115, 5.212708, 5.143295, 5.09066, 5.054367, 
    5.031552,
  // height(6,37, 0-49)
    5.005801, 5.011303, 5.021308, 5.038361, 5.065549, 5.105801, 5.160549, 
    5.228139, 5.302862, 5.375661, 5.436546, 5.477478, 5.494156, 5.486094, 
    5.455472, 5.416793, 5.425346, 5.372597, 5.313364, 5.249673, 5.182581, 
    5.122284, 5.060222, 5.003567, 4.958797, 4.929513, 4.918928, 4.928662, 
    4.958955, 5.005849, 5.063618, 5.138137, 5.217677, 5.298407, 5.37631, 
    5.447072, 5.506024, 5.548225, 5.568847, 5.564021, 5.532116, 5.475121, 
    5.399345, 5.314625, 5.231855, 5.159892, 5.10349, 5.063205, 5.036771, 
    5.020852,
  // height(6,38, 0-49)
    5.003891, 5.007699, 5.014834, 5.027377, 5.048105, 5.080132, 5.126007, 
    5.186297, 5.258187, 5.335034, 5.407619, 5.466704, 5.505548, 5.521119, 
    5.513827, 5.494351, 5.508985, 5.466975, 5.412887, 5.350326, 5.281836, 
    5.219258, 5.155951, 5.099565, 5.056434, 5.03064, 5.024622, 5.038822, 
    5.071777, 5.119378, 5.175891, 5.246482, 5.319166, 5.390081, 5.455081, 
    5.509673, 5.549134, 5.568857, 5.565062, 5.535907, 5.482723, 5.41076, 
    5.32871, 5.246728, 5.17364, 5.114793, 5.071546, 5.042262, 5.023884, 
    5.013244,
  // height(6,39, 0-49)
    5.002481, 5.004988, 5.009824, 5.01858, 5.03355, 5.057617, 5.093771, 
    5.144087, 5.20835, 5.282921, 5.360754, 5.432937, 5.491165, 5.529831, 
    5.546874, 5.548873, 5.571401, 5.542856, 5.497346, 5.439801, 5.37418, 
    5.313456, 5.252906, 5.200124, 5.160659, 5.138759, 5.136208, 5.152687, 
    5.185562, 5.231051, 5.283538, 5.347201, 5.409976, 5.467864, 5.516581, 
    5.55163, 5.568645, 5.56403, 5.53591, 5.485222, 5.416424, 5.337203, 
    5.256864, 5.183889, 5.12386, 5.078702, 5.04735, 5.027104, 5.014899, 
    5.008082,
  // height(6,40, 0-49)
    5.001506, 5.003077, 5.006195, 5.012006, 5.022259, 5.039356, 5.066173, 
    5.105471, 5.158852, 5.225492, 5.301316, 5.379313, 5.451182, 5.50957, 
    5.549834, 5.574276, 5.607434, 5.595249, 5.56227, 5.514218, 5.45616, 
    5.401567, 5.34748, 5.301089, 5.266817, 5.248916, 5.24868, 5.265357, 
    5.295565, 5.336142, 5.381646, 5.435097, 5.484591, 5.526011, 5.555113, 
    5.567804, 5.56073, 5.532122, 5.482724, 5.416423, 5.340039, 5.261992, 
    5.190205, 5.130182, 5.084167, 5.051551, 5.03001, 5.016677, 5.008926, 
    5.004739,
  // height(6,41, 0-49)
    5.000872, 5.001811, 5.003726, 5.007394, 5.014062, 5.025565, 5.044321, 
    5.073099, 5.114377, 5.169344, 5.236801, 5.312582, 5.390053, 5.461687, 
    5.521057, 5.566554, 5.612437, 5.619046, 5.602568, 5.568698, 5.523036, 
    5.478834, 5.434624, 5.396982, 5.369114, 5.355171, 5.356116, 5.371006, 
    5.396053, 5.428863, 5.464231, 5.504002, 5.536785, 5.558545, 5.565493, 
    5.554577, 5.524221, 5.475122, 5.410758, 5.337202, 5.261991, 5.192336, 
    5.133424, 5.087586, 5.054531, 5.032286, 5.018225, 5.009846, 5.005136, 
    5.00267,
  // height(6,42, 0-49)
    5.000481, 5.001017, 5.00214, 5.004345, 5.008471, 5.015812, 5.028213, 
    5.048029, 5.077842, 5.119837, 5.174886, 5.241633, 5.316115, 5.392297, 
    5.463521, 5.525497, 5.583997, 5.61024, 5.613234, 5.597641, 5.568791, 
    5.538901, 5.507612, 5.480733, 5.460288, 5.450224, 5.451291, 5.462511, 
    5.480014, 5.502224, 5.524326, 5.547166, 5.560371, 5.560421, 5.544595, 
    5.511576, 5.462096, 5.399337, 5.328705, 5.25686, 5.190202, 5.133424, 
    5.088748, 5.056075, 5.033725, 5.019349, 5.010611, 5.00558, 5.002838, 
    5.001445,
  // height(6,43, 0-49)
    5.000254, 5.000546, 5.001174, 5.002439, 5.00487, 5.009325, 5.017095, 
    5.029969, 5.050164, 5.080025, 5.121449, 5.175093, 5.239628, 5.311485, 
    5.385376, 5.456191, 5.523962, 5.567801, 5.590858, 5.595832, 5.586867, 
    5.574288, 5.558316, 5.543778, 5.53159, 5.525327, 5.525582, 5.531467, 
    5.539334, 5.548489, 5.55477, 5.558441, 5.550801, 5.52943, 5.493284, 
    5.443173, 5.382017, 5.3146, 5.246713, 5.18388, 5.130176, 5.087583, 
    5.056074, 5.034219, 5.019936, 5.011107, 5.005926, 5.003036, 5.001507, 
    5.000752,
  // height(6,44, 0-49)
    5.000128, 5.000281, 5.000617, 5.00131, 5.002675, 5.005249, 5.009875, 
    5.017793, 5.030678, 5.050543, 5.079468, 5.119081, 5.169894, 5.230724, 
    5.298507, 5.369052, 5.439737, 5.495649, 5.53579, 5.560483, 5.571956, 
    5.577868, 5.578365, 5.576972, 5.573505, 5.570918, 5.569647, 5.568985, 
    5.565864, 5.560555, 5.549966, 5.534374, 5.507415, 5.468267, 5.417797, 
    5.358663, 5.295023, 5.231793, 5.1736, 5.123836, 5.084153, 5.054524, 
    5.033722, 5.019935, 5.011277, 5.006111, 5.003177, 5.001587, 5.000769, 
    5.000376,
  // height(6,45, 0-49)
    5.000063, 5.000138, 5.000311, 5.000674, 5.001407, 5.002824, 5.005446, 
    5.010069, 5.017841, 5.03027, 5.049132, 5.07621, 5.112875, 5.159539, 
    5.21521, 5.277477, 5.343553, 5.403429, 5.454043, 5.493758, 5.522719, 
    5.545506, 5.561567, 5.57276, 5.57775, 5.578548, 5.575379, 5.567812, 
    5.55373, 5.5345, 5.508538, 5.476731, 5.435433, 5.385492, 5.329256, 
    5.270243, 5.212493, 5.159744, 5.114697, 5.078644, 5.051517, 5.032265, 
    5.019338, 5.011102, 5.00611, 5.003224, 5.001634, 5.000797, 5.000378, 
    5.000181,
  // height(6,46, 0-49)
    5.000031, 5.000067, 5.00015, 5.000331, 5.000709, 5.001454, 5.002869, 
    5.005435, 5.009881, 5.017223, 5.02877, 5.046025, 5.070468, 5.103213, 
    5.144585, 5.193819, 5.249195, 5.304764, 5.3573, 5.404286, 5.444343, 
    5.479204, 5.507306, 5.528643, 5.540705, 5.544287, 5.539324, 5.525741, 
    5.502674, 5.472641, 5.435821, 5.39402, 5.3461, 5.29405, 5.24074, 
    5.189366, 5.142821, 5.103158, 5.071325, 5.047211, 5.029928, 5.018178, 
    5.010585, 5.005913, 5.00317, 5.001631, 5.000807, 5.000385, 5.000178, 
    5.000086,
  // height(6,47, 0-49)
    5.000016, 5.000032, 5.000071, 5.000156, 5.000339, 5.000712, 5.00144, 
    5.002793, 5.0052, 5.009297, 5.015947, 5.026236, 5.041384, 5.062566, 
    5.090646, 5.125872, 5.167685, 5.213145, 5.259974, 5.305874, 5.348906, 
    5.388846, 5.423281, 5.450551, 5.467137, 5.472547, 5.466381, 5.448959, 
    5.420728, 5.385215, 5.34418, 5.300195, 5.253817, 5.207319, 5.163136, 
    5.123419, 5.089652, 5.062486, 5.041776, 5.026793, 5.016487, 5.009737, 
    5.005519, 5.003005, 5.001571, 5.000789, 5.000381, 5.000178, 5.000082, 
    5.00004,
  // height(6,48, 0-49)
    5.00001, 5.000016, 5.000032, 5.00007, 5.000153, 5.000327, 5.000675, 
    5.00134, 5.002559, 5.004692, 5.008262, 5.013968, 5.022671, 5.035318, 
    5.052807, 5.075786, 5.104437, 5.137691, 5.174414, 5.213105, 5.252073, 
    5.290257, 5.324902, 5.35331, 5.371335, 5.377446, 5.370953, 5.352503, 
    5.323604, 5.288409, 5.249669, 5.210224, 5.171314, 5.134784, 5.102191, 
    5.074564, 5.052313, 5.035273, 5.022853, 5.014224, 5.008505, 5.004887, 
    5.002697, 5.001432, 5.000731, 5.000358, 5.00017, 5.000078, 5.000036, 
    5.000019,
  // height(6,49, 0-49)
    5.000003, 5.000005, 5.00001, 5.000021, 5.000048, 5.000105, 5.000226, 
    5.000469, 5.000938, 5.001801, 5.003329, 5.005904, 5.010058, 5.016455, 
    5.025851, 5.039001, 5.056527, 5.078323, 5.104247, 5.133745, 5.165843, 
    5.199856, 5.232936, 5.261728, 5.280608, 5.287194, 5.280442, 5.261369, 
    5.232347, 5.199001, 5.164706, 5.132356, 5.102732, 5.076899, 5.055445, 
    5.038478, 5.025686, 5.016487, 5.010173, 5.006035, 5.00344, 5.001884, 
    5.000993, 5.000504, 5.000246, 5.000115, 5.000053, 5.000024, 5.000012, 
    5.000007,
  // height(7,0, 0-49)
    5.000065, 5.000127, 5.000259, 5.000518, 5.001007, 5.001891, 5.003428, 
    5.005995, 5.010108, 5.016434, 5.025755, 5.038896, 5.056596, 5.079338, 
    5.107157, 5.139503, 5.175241, 5.211763, 5.247095, 5.279533, 5.307879, 
    5.331899, 5.350907, 5.364714, 5.372608, 5.374767, 5.371186, 5.361848, 
    5.346594, 5.326201, 5.300992, 5.271825, 5.239199, 5.204507, 5.169468, 
    5.135854, 5.105211, 5.078644, 5.05671, 5.039443, 5.026458, 5.017118, 
    5.010684, 5.006434, 5.003739, 5.002098, 5.001138, 5.000597, 5.000308, 
    5.000164,
  // height(7,1, 0-49)
    5.000121, 5.000238, 5.00048, 5.000947, 5.001812, 5.003347, 5.005964, 
    5.010249, 5.016973, 5.027078, 5.041602, 5.061525, 5.087564, 5.119916, 
    5.158052, 5.20067, 5.245986, 5.289452, 5.328742, 5.362245, 5.389309, 
    5.411021, 5.42722, 5.438537, 5.444373, 5.445482, 5.441986, 5.433731, 
    5.419994, 5.40147, 5.377745, 5.349227, 5.315303, 5.277005, 5.236064, 
    5.194644, 5.154975, 5.118989, 5.08803, 5.062733, 5.043062, 5.028478, 
    5.018152, 5.011154, 5.00661, 5.003779, 5.002086, 5.001116, 5.000584, 
    5.000315,
  // height(7,2, 0-49)
    5.000235, 5.000459, 5.00091, 5.001763, 5.003306, 5.005982, 5.010434, 
    5.017533, 5.028368, 5.04416, 5.066104, 5.095097, 5.131435, 5.174539, 
    5.222845, 5.274029, 5.325931, 5.371635, 5.409235, 5.437857, 5.457925, 
    5.47228, 5.481415, 5.48696, 5.488639, 5.487854, 5.484875, 5.479411, 
    5.470135, 5.457471, 5.440103, 5.41785, 5.388554, 5.352391, 5.310528, 
    5.264997, 5.218402, 5.17348, 5.132623, 5.097514, 5.068947, 5.046889, 
    5.030686, 5.019336, 5.011737, 5.006867, 5.003877, 5.00212, 5.001133, 
    5.000619,
  // height(7,3, 0-49)
    5.000447, 5.000865, 5.001686, 5.003202, 5.005878, 5.010405, 5.017734, 
    5.029084, 5.045851, 5.069425, 5.100871, 5.14055, 5.18778, 5.240693, 
    5.296419, 5.351787, 5.405229, 5.447082, 5.476982, 5.495352, 5.503921, 
    5.507381, 5.506683, 5.504385, 5.500591, 5.497306, 5.494962, 5.493176, 
    5.490098, 5.485869, 5.478354, 5.466926, 5.447763, 5.419919, 5.383484, 
    5.339691, 5.290837, 5.239985, 5.190429, 5.145115, 5.106135, 5.074507, 
    5.050228, 5.032541, 5.020276, 5.012163, 5.007035, 5.003933, 5.00215, 
    5.001194,
  // height(7,4, 0-49)
    5.00083, 5.001577, 5.003015, 5.005607, 5.010071, 5.01742, 5.028973, 
    5.046284, 5.070925, 5.104134, 5.146344, 5.196767, 5.253208, 5.312281, 
    5.370041, 5.423226, 5.472451, 5.504696, 5.522296, 5.52714, 5.522073, 
    5.513369, 5.501997, 5.491229, 5.481532, 5.475423, 5.473501, 5.47537, 
    5.478836, 5.483813, 5.487583, 5.489424, 5.484031, 5.469409, 5.444396, 
    5.408932, 5.364272, 5.312967, 5.258545, 5.204911, 5.155597, 5.11315, 
    5.078824, 5.052646, 5.033748, 5.020789, 5.012327, 5.007061, 5.003947, 
    5.002234,
  // height(7,5, 0-49)
    5.00148, 5.002769, 5.005187, 5.009442, 5.016574, 5.027974, 5.045319, 
    5.070355, 5.104497, 5.148292, 5.200894, 5.259817, 5.321171, 5.380404, 
    5.433293, 5.477595, 5.517872, 5.536584, 5.539735, 5.53039, 5.512024, 
    5.492009, 5.470812, 5.452157, 5.436851, 5.427817, 5.425859, 5.430663, 
    5.439898, 5.453335, 5.467922, 5.483245, 5.492867, 5.494058, 5.484577, 
    5.462999, 5.429098, 5.384137, 5.330914, 5.273443, 5.216244, 5.163455, 
    5.118066, 5.081542, 5.053911, 5.034173, 5.020812, 5.012223, 5.006996, 
    5.004036,
  // height(7,6, 0-49)
    5.002537, 5.004672, 5.008571, 5.015256, 5.026145, 5.042995, 5.067703, 
    5.101876, 5.146226, 5.199944, 5.260352, 5.323129, 5.38313, 5.435542, 
    5.476911, 5.507005, 5.535779, 5.539415, 5.528361, 5.50633, 5.476847, 
    5.447856, 5.418829, 5.393694, 5.373574, 5.361693, 5.35911, 5.365716, 
    5.379266, 5.39945, 5.423106, 5.450462, 5.474294, 5.491517, 5.499191, 
    5.494801, 5.476672, 5.444415, 5.399313, 5.344433, 5.284281, 5.224, 
    5.16831, 5.120595, 5.082476, 5.053929, 5.033796, 5.020385, 5.011956, 
    5.007038,
  // height(7,7, 0-49)
    5.004174, 5.007567, 5.013592, 5.023635, 5.039485, 5.063149, 5.09643, 
    5.140269, 5.194015, 5.254954, 5.318458, 5.378851, 5.430717, 5.47008, 
    5.495052, 5.507923, 5.524962, 5.513952, 5.490565, 5.458614, 5.421184, 
    5.386325, 5.352101, 5.322395, 5.298602, 5.284111, 5.280297, 5.287394, 
    5.303493, 5.328266, 5.358603, 5.39561, 5.431551, 5.463284, 5.487547, 
    5.501169, 5.501382, 5.486283, 5.455358, 5.409954, 5.353441, 5.290848, 
    5.227934, 5.169954, 5.120609, 5.081582, 5.052734, 5.032722, 5.019694, 
    5.011834,
  // height(7,8, 0-49)
    5.006591, 5.011756, 5.020663, 5.035065, 5.057024, 5.088521, 5.130782, 
    5.183451, 5.243975, 5.307598, 5.368227, 5.41984, 5.457864, 5.479952, 
    5.486041, 5.480951, 5.487695, 5.463608, 5.430469, 5.391768, 5.349826, 
    5.31244, 5.275925, 5.243874, 5.217835, 5.201171, 5.195599, 5.201853, 
    5.21865, 5.245731, 5.280169, 5.3241, 5.369467, 5.413232, 5.452092, 
    5.482594, 5.501349, 5.505374, 5.492573, 5.462371, 5.416243, 5.357937, 
    5.29305, 5.227945, 5.16834, 5.118135, 5.078969, 5.050519, 5.031245, 
    5.019186,
  // height(7,9, 0-49)
    5.009975, 5.017505, 5.030089, 5.049776, 5.078679, 5.118333, 5.168806, 
    5.227921, 5.291047, 5.351834, 5.403693, 5.44137, 5.461924, 5.464885, 
    5.451752, 5.429615, 5.428216, 5.392973, 5.352669, 5.310205, 5.26699, 
    5.230297, 5.194464, 5.162518, 5.135951, 5.117805, 5.110119, 5.114284, 
    5.12995, 5.157085, 5.193079, 5.241197, 5.293196, 5.346199, 5.396987, 
    5.442087, 5.477869, 5.500757, 5.507577, 5.49611, 5.465787, 5.418324, 
    5.357944, 5.290869, 5.224051, 5.163567, 5.113378, 5.074952, 5.047724, 
    5.029982,
  // height(7,10, 0-49)
    5.01446, 5.02496, 5.041936, 5.067563, 5.103665, 5.150827, 5.207461, 
    5.269351, 5.330144, 5.382782, 5.421267, 5.441902, 5.443639, 5.42762, 
    5.396376, 5.358976, 5.351389, 5.30677, 5.26151, 5.217797, 5.176116, 
    5.143035, 5.110799, 5.081596, 5.056532, 5.03793, 5.028039, 5.029017, 
    5.041786, 5.066779, 5.101882, 5.151564, 5.207518, 5.267011, 5.326935, 
    5.383892, 5.434252, 5.474237, 5.500106, 5.508534, 5.497243, 5.465786, 
    5.416254, 5.353475, 5.284362, 5.216415, 5.155936, 5.106784, 5.070136, 
    5.045145,
  // height(7,11, 0-49)
    5.020058, 5.034059, 5.055914, 5.087668, 5.130448, 5.183438, 5.24315, 
    5.303562, 5.357356, 5.397788, 5.420244, 5.422883, 5.40632, 5.37279, 
    5.325267, 5.274648, 5.261842, 5.209301, 5.160816, 5.117825, 5.079991, 
    5.053068, 5.027225, 5.003541, 4.982328, 4.9647, 4.952865, 4.949788, 
    4.957981, 4.978666, 5.010483, 5.059205, 5.116598, 5.180028, 5.246441, 
    5.312511, 5.374698, 5.429252, 5.472255, 5.499822, 5.50852, 5.4961, 
    5.46238, 5.410001, 5.344549, 5.27369, 5.205394, 5.146018, 5.099126, 
    5.065478,
  // height(7,12, 0-49)
    5.026608, 5.044453, 5.071303, 5.108771, 5.156913, 5.213257, 5.272523, 
    5.327488, 5.37078, 5.396759, 5.402548, 5.387994, 5.354888, 5.305989, 
    5.244225, 5.182299, 5.163545, 5.104256, 5.053853, 5.013101, 4.980991, 
    4.962399, 4.945583, 4.930279, 4.915555, 4.900771, 4.887709, 4.880032, 
    4.882082, 4.896287, 4.922391, 4.967634, 5.024047, 5.089039, 5.159525, 
    5.232173, 5.303509, 5.369896, 5.427476, 5.472199, 5.500046, 5.507537, 
    5.492572, 5.455415, 5.399471, 5.33125, 5.259198, 5.191624, 5.134699, 
    5.091459,
  // height(7,13, 0-49)
    5.033735, 5.05548, 5.086987, 5.129162, 5.180753, 5.237656, 5.293234, 
    5.339825, 5.370763, 5.381915, 5.372065, 5.342326, 5.295123, 5.233254, 
    5.159248, 5.08756, 5.059693, 4.994692, 4.943421, 4.906126, 4.881305, 
    4.872905, 4.867583, 4.863523, 4.858131, 4.848498, 4.835467, 4.823103, 
    4.817653, 4.823181, 4.841021, 4.880143, 4.933115, 4.997382, 5.069714, 
    5.146647, 5.224686, 5.300283, 5.36973, 5.429057, 5.474072, 5.500647, 
    5.505333, 5.486337, 5.44461, 5.384568, 5.313798, 5.241476, 5.176003, 
    5.123024,
  // height(7,14, 0-49)
    5.040861, 5.066214, 5.101596, 5.147029, 5.199935, 5.254867, 5.304424, 
    5.34119, 5.35965, 5.357197, 5.333939, 5.29176, 5.233256, 5.160916, 
    5.076638, 4.99614, 4.952772, 4.88308, 4.831912, 4.799187, 4.783082, 
    4.786512, 4.794985, 4.804932, 4.811784, 4.809976, 4.798848, 4.782353, 
    4.768427, 4.763132, 4.769983, 4.80008, 4.846959, 4.908147, 4.980169, 
    5.059281, 5.141819, 5.224236, 5.302959, 5.374205, 5.433871, 5.477612, 
    5.501223, 5.501401, 5.476885, 5.429611, 5.365265, 5.292587, 5.221282, 
    5.159416,
  // height(7,15, 0-49)
    5.04727, 5.075588, 5.113734, 5.160819, 5.213135, 5.26433, 5.306828, 
    5.333897, 5.341276, 5.327645, 5.294003, 5.242578, 5.175807, 5.095669, 
    5.003297, 4.913842, 4.844732, 4.771318, 4.721283, 4.694343, 4.688432, 
    4.705205, 4.729593, 4.756072, 4.777933, 4.786829, 4.780121, 4.760928, 
    4.738266, 4.720271, 4.713288, 4.731091, 4.768864, 4.824393, 4.893883, 
    4.973128, 5.058129, 5.145205, 5.230836, 5.311429, 5.383089, 5.441543, 
    5.482284, 5.501088, 5.494987, 5.46355, 5.410028, 5.341596, 5.268045, 
    5.19916,
  // height(7,16, 0-49)
    5.052221, 5.082582, 5.122238, 5.169528, 5.219952, 5.266737, 5.302544, 
    5.321485, 5.320392, 5.298859, 5.258375, 5.201202, 5.129457, 5.044556, 
    4.946846, 4.846074, 4.737124, 4.660678, 4.612901, 4.593229, 4.599227, 
    4.630776, 4.672967, 4.718068, 4.757268, 4.779699, 4.780499, 4.761142, 
    4.730637, 4.698801, 4.675304, 4.677201, 4.702387, 4.749299, 4.813816, 
    4.891094, 4.976588, 5.066315, 5.156695, 5.244262, 5.325356, 5.395911, 
    5.45143, 5.487248, 5.499257, 5.485078, 5.445483, 5.385374, 5.313462, 
    5.240213,
  // height(7,17, 0-49)
    5.055084, 5.086399, 5.126359, 5.172816, 5.22089, 5.263784, 5.294598, 
    5.308188, 5.302143, 5.27656, 5.233084, 5.173849, 5.100662, 5.014484, 
    4.914962, 4.796424, 4.630887, 4.5516, 4.507199, 4.496636, 4.516641, 
    4.564325, 4.625845, 4.690973, 4.749099, 4.787496, 4.799221, 4.783396, 
    4.747558, 4.702156, 4.66026, 4.64256, 4.651261, 4.686162, 4.742951, 
    4.81599, 4.899972, 4.990417, 5.083542, 5.175914, 5.264064, 5.344178, 
    5.411934, 5.462564, 5.491307, 5.494365, 5.470315, 5.421548, 5.354854, 
    5.280277,
  // height(7,18, 0-49)
    5.055455, 5.086561, 5.125804, 5.170914, 5.217056, 5.257705, 5.286389, 
    5.298403, 5.291608, 5.26616, 5.223593, 5.165879, 5.094666, 5.010685, 
    4.912883, 4.764289, 4.52522, 4.443193, 4.403152, 4.403866, 4.440429, 
    4.50552, 4.587378, 4.673081, 4.750764, 4.806866, 4.832855, 4.825094, 
    4.788147, 4.731499, 4.671028, 4.630623, 4.61889, 4.638094, 4.684124, 
    4.750472, 4.830854, 4.920098, 5.014065, 5.109241, 5.202271, 5.289577, 
    5.367074, 5.430085, 5.473558, 5.492756, 5.484509, 5.448822, 5.390132, 
    5.31718,
  // height(7,19, 0-49)
    5.053221, 5.082938, 5.120615, 5.164308, 5.209677, 5.250699, 5.281166, 
    5.296271, 5.293453, 5.272348, 5.234126, 5.180676, 5.113756, 5.033909, 
    4.938658, 4.742922, 4.415196, 4.33217, 4.297563, 4.311978, 4.368104, 
    4.45188, 4.554541, 4.660558, 4.75763, 4.832474, 4.875569, 4.880461, 
    4.847667, 4.784114, 4.707324, 4.64267, 4.607326, 4.607371, 4.639596, 
    4.696743, 4.771411, 4.857562, 4.950556, 5.046688, 5.142635, 5.234991, 
    5.319911, 5.392896, 5.448824, 5.4824, 5.489161, 5.467055, 5.418115, 
    5.349228,
  // height(7,20, 0-49)
    5.047519, 5.072911, 5.105344, 5.143125, 5.182673, 5.219129, 5.247638, 
    5.264693, 5.268921, 5.261077, 5.243481, 5.219299, 5.191885, 5.164235, 
    5.138397, 0, 4.114454, 4.114334, 4.146542, 4.211831, 4.306983, 4.4182, 
    4.544752, 4.671088, 4.786033, 4.877743, 4.936459, 4.953573, 4.925799, 
    4.857228, 4.766321, 4.677095, 4.616313, 4.594654, 4.610526, 4.65621, 
    4.723191, 4.804475, 4.894822, 4.990243, 5.087366, 5.182891, 5.273173, 
    5.353907, 5.420018, 5.465905, 5.486187, 5.477157, 5.438637, 5.375458,
  // height(7,21, 0-49)
    5.042906, 5.065928, 5.096264, 5.132921, 5.173195, 5.212954, 5.247571, 
    5.273136, 5.287375, 5.289968, 5.282302, 5.266943, 5.247061, 5.225951, 
    5.206573, 0, 3.960332, 3.978011, 4.033281, 4.12433, 4.2451, 4.375662, 
    4.518851, 4.658369, 4.784651, 4.88853, 4.961393, 4.993842, 4.979385, 
    4.918301, 4.827318, 4.723927, 4.643672, 4.602317, 4.601614, 4.634759, 
    4.692778, 4.76789, 4.85425, 4.947518, 5.044199, 5.141039, 5.234534, 
    5.320562, 5.394155, 5.449563, 5.480793, 5.482881, 5.453789, 5.39637,
  // height(7,22, 0-49)
    5.039219, 5.060489, 5.089365, 5.125412, 5.166588, 5.209273, 5.24895, 
    5.281309, 5.303318, 5.313817, 5.313527, 5.304658, 5.290368, 5.274252, 
    5.259961, 0, 3.835406, 3.868202, 3.942687, 4.05515, 4.197188, 4.343217, 
    4.499814, 4.650155, 4.786009, 4.900363, 4.985329, 5.030774, 5.027747, 
    4.973923, 4.885179, 4.770913, 4.6747, 4.616134, 4.600175, 4.62134, 
    4.670562, 4.739481, 4.821707, 4.912546, 5.008337, 5.105797, 5.201505, 
    5.291459, 5.370781, 5.433647, 5.473652, 5.484908, 5.46392, 5.41185,
  // height(7,23, 0-49)
    5.037024, 5.057234, 5.085255, 5.120999, 5.162849, 5.207517, 5.250546, 
    5.287356, 5.314402, 5.329967, 5.334363, 5.329612, 5.318913, 5.30611, 
    5.295335, 0, 3.75083, 3.794178, 3.882296, 4.009888, 4.166729, 4.322514, 
    4.487185, 4.643687, 4.784962, 4.90581, 4.999001, 5.054017, 5.060269, 
    5.013733, 4.929824, 4.809685, 4.70313, 4.632049, 4.604081, 4.615284, 
    4.656912, 4.720334, 4.798786, 4.887294, 4.982037, 5.079676, 5.176805, 
    5.269478, 5.352865, 5.421083, 5.467453, 5.485446, 5.470525, 5.42257,
  // height(7,24, 0-49)
    5.036716, 5.05663, 5.084397, 5.120026, 5.162042, 5.207297, 5.25141, 
    5.289758, 5.318656, 5.336201, 5.342546, 5.339622, 5.330624, 5.319474, 
    5.310493, 0, 3.710093, 3.758837, 3.854186, 3.98978, 4.154303, 4.314251, 
    4.482039, 4.640524, 4.783451, 4.906882, 5.004126, 5.064573, 5.076762, 
    5.03577, 4.956805, 4.834767, 4.72329, 4.645191, 4.609799, 4.614413, 
    4.65074, 4.710127, 4.785641, 4.872161, 4.96578, 5.063129, 5.160812, 
    5.254916, 5.340633, 5.41205, 5.462324, 5.484553, 5.473571, 5.428463,
  // height(7,25, 0-49)
    5.038471, 5.058876, 5.086976, 5.122606, 5.164133, 5.208367, 5.251034, 
    5.287758, 5.315138, 5.33149, 5.337061, 5.33376, 5.324667, 5.313553, 
    5.304569, 0, 3.712392, 3.76137, 3.857336, 3.993675, 4.158824, 4.318006, 
    4.484923, 4.642324, 4.784227, 4.907133, 5.004549, 5.065886, 5.079467, 
    5.040195, 4.963305, 4.841302, 4.72898, 4.649186, 4.611698, 4.614275, 
    4.648862, 4.706868, 4.781345, 4.867144, 4.960334, 5.057543, 5.155376, 
    5.249931, 5.336409, 5.408885, 5.460465, 5.484119, 5.474478, 5.430358,
  // height(7,26, 0-49)
    5.042217, 5.063863, 5.092844, 5.128556, 5.168951, 5.210625, 5.24946, 
    5.281579, 5.304241, 5.31635, 5.31849, 5.312615, 5.301614, 5.288908, 
    5.278151, 0, 3.755883, 3.80003, 3.890133, 4.020155, 4.179138, 4.333121, 
    4.495686, 4.649438, 4.788105, 4.907743, 5.001677, 5.059398, 5.069646, 
    5.02778, 4.949212, 4.828493, 4.718805, 4.642381, 4.608218, 4.613591, 
    4.650334, 4.709931, 4.785549, 4.872119, 4.96576, 5.06312, 5.160808, 
    5.254914, 5.340632, 5.412049, 5.462324, 5.484553, 5.473571, 5.428463,
  // height(7,27, 0-49)
    5.047648, 5.071205, 5.101556, 5.137453, 5.176219, 5.214128, 5.247229, 
    5.272307, 5.287539, 5.292675, 5.288845, 5.278172, 5.26337, 5.247412, 
    5.233242, 0, 3.837907, 3.872372, 3.950503, 4.067498, 4.213774, 4.358329, 
    4.513062, 4.660518, 4.793601, 4.907108, 4.993864, 5.043576, 5.046104, 
    4.997985, 4.914999, 4.797587, 4.69459, 4.626752, 4.60112, 4.613746, 
    4.65615, 4.719967, 4.798612, 4.887213, 4.981999, 5.079659, 5.176796, 
    5.269475, 5.352864, 5.421082, 5.467452, 5.485446, 5.470524, 5.42257,
  // height(7,28, 0-49)
    5.054279, 5.08032, 5.1125, 5.148775, 5.185695, 5.219107, 5.245215, 
    5.261521, 5.267226, 5.263089, 5.25097, 5.233331, 5.212831, 5.192018, 
    5.172996, 0, 3.95486, 3.975625, 4.036456, 4.134297, 4.261631, 4.392307, 
    4.535101, 4.672795, 4.797129, 4.90109, 4.976916, 5.014869, 5.006731, 
    4.951005, 4.863965, 4.753953, 4.662951, 4.608952, 4.596192, 4.619275, 
    4.669537, 4.738986, 4.821471, 4.912435, 5.008284, 5.105772, 5.201493, 
    5.291453, 5.370779, 5.433645, 5.473652, 5.484908, 5.46392, 5.41185,
  // height(7,29, 0-49)
    5.061519, 5.090569, 5.125088, 5.162135, 5.197347, 5.22602, 5.244443, 
    5.250815, 5.245413, 5.230116, 5.207698, 5.181172, 5.153317, 5.126302, 
    5.101217, 0, 4.100039, 4.105047, 4.144559, 4.218102, 4.320959, 4.433148, 
    4.559563, 4.683653, 4.795854, 4.887011, 4.948723, 4.97219, 4.951942, 
    4.889277, 4.801144, 4.70358, 4.629909, 4.594042, 4.597061, 4.6324, 
    4.6916, 4.767314, 4.853972, 4.947385, 5.044137, 5.141009, 5.23452, 
    5.320555, 5.394152, 5.449561, 5.480793, 5.482881, 5.453789, 5.396369,
  // height(7,30, 0-49)
    5.069942, 5.104444, 5.145037, 5.188226, 5.228665, 5.260446, 5.278681, 
    5.280539, 5.265384, 5.23421, 5.188872, 5.131349, 5.06307, 4.983942, 
    4.890614, 4.694397, 4.378685, 4.306954, 4.281877, 4.30549, 4.370964, 
    4.459809, 4.568273, 4.679267, 4.780853, 4.860884, 4.909776, 4.919673, 
    4.888474, 4.82117, 4.735869, 4.654694, 4.601761, 4.586124, 4.605887, 
    4.653808, 4.721985, 4.803879, 4.89453, 4.990101, 5.087297, 5.182858, 
    5.273158, 5.353899, 5.420014, 5.465903, 5.486187, 5.477157, 5.438637, 
    5.375458,
  // height(7,31, 0-49)
    5.073872, 5.110393, 5.153061, 5.197888, 5.238931, 5.269813, 5.28551, 
    5.283435, 5.26344, 5.227028, 5.17638, 5.113566, 5.040033, 4.956133, 
    4.860312, 4.711382, 4.476999, 4.403505, 4.371749, 4.381316, 4.427418, 
    4.499416, 4.589086, 4.681817, 4.765648, 4.827684, 4.859194, 4.855018, 
    4.817186, 4.75356, 4.681082, 4.623222, 4.59458, 4.599795, 4.6354, 
    4.694525, 4.770272, 4.856986, 4.950268, 5.046546, 5.142564, 5.234956, 
    5.319895, 5.392888, 5.448821, 5.482398, 5.48916, 5.467055, 5.418115, 
    5.349227,
  // height(7,32, 0-49)
    5.074563, 5.111968, 5.156186, 5.203183, 5.24673, 5.279979, 5.297396, 
    5.296023, 5.275575, 5.23764, 5.184599, 5.118748, 5.041742, 4.954269, 
    4.855663, 4.736937, 4.571723, 4.498174, 4.459996, 4.456672, 4.485158, 
    4.540483, 4.610906, 4.684608, 4.750361, 4.79529, 4.81181, 4.797491, 
    4.758013, 4.70317, 4.647774, 4.613843, 4.608014, 4.631615, 4.680494, 
    4.748522, 4.829835, 4.919573, 5.013799, 5.109106, 5.202204, 5.289543, 
    5.367058, 5.430077, 5.473555, 5.492754, 5.484507, 5.448821, 5.390131, 
    5.31718,
  // height(7,33, 0-49)
    5.072055, 5.109157, 5.154137, 5.203316, 5.250513, 5.288494, 5.311002, 
    5.31429, 5.297483, 5.261912, 5.210007, 5.14432, 5.066876, 4.978845, 
    4.880323, 4.778907, 4.66792, 4.594558, 4.550687, 4.536237, 4.549191, 
    4.588276, 4.639575, 4.693966, 4.741624, 4.770691, 4.775239, 4.755387, 
    4.719284, 4.677091, 4.640542, 4.628673, 4.642346, 4.680838, 4.739939, 
    4.814349, 4.8991, 4.989961, 5.083307, 5.175795, 5.264003, 5.344147, 
    5.411918, 5.462556, 5.491303, 5.494362, 5.470314, 5.421547, 5.354854, 
    5.280277,
  // height(7,34, 0-49)
    5.066685, 5.102252, 5.146866, 5.197575, 5.248649, 5.292713, 5.322759, 
    5.333969, 5.324487, 5.295034, 5.247876, 5.185752, 5.11112, 5.025746, 
    4.930516, 4.839296, 4.766814, 4.694075, 4.645786, 4.622183, 4.62171, 
    4.645421, 4.67846, 4.714131, 4.744484, 4.759594, 4.755527, 4.734432, 
    4.705405, 4.677551, 4.65919, 4.666082, 4.695303, 4.745059, 4.811397, 
    4.889759, 4.975869, 5.065935, 5.156497, 5.244161, 5.325305, 5.395886, 
    5.451417, 5.487242, 5.499254, 5.485077, 5.445483, 5.385374, 5.313462, 
    5.240213,
  // height(7,35, 0-49)
    5.059091, 5.091941, 5.134801, 5.18574, 5.23992, 5.290249, 5.329171, 
    5.350695, 5.351656, 5.331776, 5.292833, 5.237574, 5.16882, 5.088939, 
    4.999584, 4.915709, 4.867932, 4.796804, 4.745568, 4.71463, 4.70265, 
    4.712214, 4.728501, 4.746943, 4.761694, 4.765309, 4.755863, 4.73676, 
    4.716686, 4.702873, 4.700494, 4.722412, 4.763369, 4.821098, 4.89199, 
    4.972076, 5.057559, 5.144899, 5.230677, 5.311346, 5.383048, 5.441524, 
    5.482273, 5.501082, 5.494984, 5.463549, 5.410028, 5.341596, 5.268045, 
    5.19916,
  // height(7,36, 0-49)
    5.050116, 5.079262, 5.118917, 5.168323, 5.223925, 5.279467, 5.327296, 
    5.360398, 5.374112, 5.366771, 5.339256, 5.293997, 5.233984, 5.162076, 
    5.080613, 5.003589, 4.970191, 4.901921, 4.849092, 4.81234, 4.790542, 
    4.787408, 4.788884, 4.792263, 4.793777, 4.788606, 4.776517, 4.761394, 
    4.750595, 4.749277, 4.760054, 4.793442, 4.842779, 4.90564, 4.978724, 
    5.058472, 5.141376, 5.223999, 5.302834, 5.37414, 5.433838, 5.477597, 
    5.501214, 5.501397, 5.476884, 5.429609, 5.365265, 5.292587, 5.221282, 
    5.159416,
  // height(7,37, 0-49)
    5.040674, 5.065457, 5.100637, 5.146596, 5.201307, 5.259878, 5.315217, 
    5.359754, 5.387404, 5.394824, 5.381534, 5.34921, 5.300679, 5.239072, 
    5.167283, 5.097776, 5.072126, 5.007897, 4.954634, 4.913358, 4.883272, 
    4.869039, 4.857895, 4.848771, 4.839742, 4.828416, 4.815767, 4.805543, 
    4.803319, 4.812391, 4.833456, 4.87515, 4.92999, 4.995509, 5.06863, 
    5.146039, 5.224351, 5.300103, 5.369635, 5.429007, 5.474048, 5.500636, 
    5.505328, 5.486333, 5.444608, 5.384567, 5.313798, 5.241476, 5.176003, 
    5.123024,
  // height(7,38, 0-49)
    5.031587, 5.051754, 5.081593, 5.122414, 5.173713, 5.232343, 5.292474, 
    5.346719, 5.387997, 5.411265, 5.414304, 5.39752, 5.363111, 5.314147, 
    5.253855, 5.193147, 5.17178, 5.112633, 5.059998, 5.015416, 4.978568, 
    4.954986, 4.933573, 4.914676, 4.897844, 4.882706, 4.870935, 4.86574, 
    4.870833, 4.888049, 4.916724, 4.963934, 5.021742, 5.087658, 5.158724, 
    5.231721, 5.303259, 5.369761, 5.427405, 5.472163, 5.500027, 5.507529, 
    5.492567, 5.455412, 5.39947, 5.33125, 5.259198, 5.191624, 5.134699, 
    5.091459,
  // height(7,39, 0-49)
    5.023478, 5.03917, 5.063326, 5.09785, 5.143517, 5.198998, 5.260269, 
    5.32098, 5.373845, 5.412485, 5.432821, 5.433532, 5.415639, 5.38168, 
    5.334877, 5.284673, 5.266556, 5.213517, 5.162659, 5.11611, 5.074186, 
    5.043216, 5.01401, 4.988095, 4.966056, 4.949053, 4.939028, 4.938462, 
    4.949347, 4.97249, 5.0063, 5.056495, 5.114914, 5.179015, 5.245848, 
    5.312171, 5.374506, 5.429146, 5.472199, 5.499791, 5.508503, 5.496091, 
    5.462376, 5.409999, 5.344549, 5.273689, 5.205394, 5.146018, 5.099126, 
    5.065478,
  // height(7,40, 0-49)
    5.01671, 5.028383, 5.047037, 5.074806, 5.113331, 5.162851, 5.22134, 
    5.284199, 5.344914, 5.396571, 5.433529, 5.452536, 5.452931, 5.436152, 
    5.404949, 5.367265, 5.35313, 5.307418, 5.259766, 5.2129, 5.167883, 
    5.131764, 5.097353, 5.067103, 5.04221, 5.024868, 5.016986, 5.020291, 
    5.035318, 5.062237, 5.098837, 5.149593, 5.206281, 5.266251, 5.326477, 
    5.383618, 5.434089, 5.474142, 5.500051, 5.508503, 5.497226, 5.465776, 
    5.416249, 5.353471, 5.28436, 5.216414, 5.155935, 5.106784, 5.070136, 
    5.045145,
  // height(7,41, 0-49)
    5.011393, 5.019699, 5.033443, 5.054687, 5.08547, 5.127131, 5.179427, 
    5.239829, 5.303455, 5.363914, 5.414792, 5.451157, 5.470404, 5.472347, 
    5.458686, 5.435668, 5.427438, 5.390626, 5.348041, 5.302955, 5.257243, 
    5.218533, 5.181604, 5.149585, 5.123898, 5.107349, 5.101637, 5.107809, 
    5.125257, 5.153823, 5.190883, 5.239744, 5.292246, 5.345578, 5.396583, 
    5.44182, 5.477694, 5.500643, 5.507504, 5.496064, 5.465759, 5.418307, 
    5.357935, 5.290864, 5.224049, 5.163566, 5.113376, 5.074951, 5.047723, 
    5.029982,
  // height(7,42, 0-49)
    5.007448, 5.013103, 5.022773, 5.03824, 5.061559, 5.094617, 5.138445, 
    5.192428, 5.253744, 5.317492, 5.377594, 5.428209, 5.465016, 5.485915, 
    5.491031, 5.484582, 5.484806, 5.458848, 5.423669, 5.382972, 5.339408, 
    5.300989, 5.264325, 5.232959, 5.208259, 5.193301, 5.189502, 5.197357, 
    5.215441, 5.243477, 5.278582, 5.322964, 5.368637, 5.412613, 5.451626, 
    5.482244, 5.501094, 5.50519, 5.492446, 5.462286, 5.416188, 5.357902, 
    5.293029, 5.227933, 5.168333, 5.118133, 5.078968, 5.050518, 5.031245, 
    5.019185,
  // height(7,43, 0-49)
    5.004671, 5.00836, 5.014862, 5.025596, 5.042367, 5.06715, 5.101645, 
    5.146619, 5.201205, 5.262506, 5.325803, 5.385471, 5.436242, 5.474329, 
    5.498009, 5.509168, 5.520347, 5.507353, 5.482279, 5.449014, 5.41083, 
    5.375861, 5.342307, 5.313881, 5.291713, 5.278893, 5.276544, 5.284764, 
    5.301612, 5.326838, 5.35743, 5.394591, 5.430645, 5.462481, 5.486856, 
    5.500595, 5.500926, 5.485937, 5.455106, 5.409778, 5.353324, 5.290773, 
    5.22789, 5.169929, 5.120594, 5.081575, 5.05273, 5.03272, 5.019693, 
    5.011834,
  // height(7,44, 0-49)
    5.002813, 5.005119, 5.009302, 5.016413, 5.027887, 5.045482, 5.071043, 
    5.106079, 5.151144, 5.205262, 5.265625, 5.327862, 5.386883, 5.437991, 
    5.477863, 5.506032, 5.529777, 5.531497, 5.519186, 5.496544, 5.467158, 
    5.438933, 5.411334, 5.388013, 5.36974, 5.359428, 5.357933, 5.365097, 
    5.378753, 5.398783, 5.422194, 5.449341, 5.473051, 5.490255, 5.498004, 
    5.493757, 5.475805, 5.443734, 5.398806, 5.344073, 5.284039, 5.223843, 
    5.168211, 5.120537, 5.082442, 5.053911, 5.033787, 5.020379, 5.011954, 
    5.007036,
  // height(7,45, 0-49)
    5.001627, 5.00301, 5.005588, 5.010087, 5.017568, 5.029425, 5.047313, 
    5.072919, 5.10756, 5.151648, 5.204203, 5.262649, 5.32308, 5.380993, 
    5.432267, 5.474555, 5.510695, 5.527712, 5.530097, 5.520863, 5.503451, 
    5.485116, 5.466168, 5.449955, 5.436787, 5.429237, 5.42793, 5.432586, 
    5.441073, 5.453529, 5.467171, 5.481771, 5.49093, 5.491922, 5.482465, 
    5.461075, 5.427461, 5.382823, 5.329916, 5.272722, 5.215748, 5.163129, 
    5.11786, 5.081418, 5.053839, 5.034134, 5.020792, 5.012212, 5.00699, 
    5.004033,
  // height(7,46, 0-49)
    5.000904, 5.001698, 5.003219, 5.005941, 5.01059, 5.018181, 5.030026, 
    5.047634, 5.072513, 5.105799, 5.147814, 5.197673, 5.25313, 5.310821, 
    5.366889, 5.418075, 5.464053, 5.494967, 5.512374, 5.518117, 5.514961, 
    5.509031, 5.500986, 5.493574, 5.486524, 5.481907, 5.480128, 5.480912, 
    5.48242, 5.485212, 5.486995, 5.487328, 5.480935, 5.465807, 5.440713, 
    5.405491, 5.361278, 5.310514, 5.256648, 5.203514, 5.154617, 5.112494, 
    5.078404, 5.052387, 5.033595, 5.020703, 5.01228, 5.007036, 5.003934, 
    5.002227,
  // height(7,47, 0-49)
    5.000479, 5.000916, 5.001769, 5.003335, 5.006079, 5.010685, 5.018091, 
    5.029477, 5.046185, 5.069523, 5.100471, 5.139313, 5.185328, 5.236683, 
    5.29062, 5.344086, 5.395159, 5.436237, 5.466683, 5.48693, 5.498612, 
    5.506318, 5.510494, 5.51297, 5.512695, 5.511067, 5.508265, 5.504123, 
    5.497348, 5.489172, 5.47811, 5.463986, 5.442956, 5.414068, 5.377319, 
    5.333785, 5.285583, 5.235593, 5.186958, 5.142507, 5.104268, 5.07323, 
    5.049392, 5.032015, 5.019961, 5.011981, 5.006932, 5.003879, 5.00212, 
    5.001179,
  // height(7,48, 0-49)
    5.000237, 5.00046, 5.000906, 5.001745, 5.003255, 5.005858, 5.010167, 
    5.017009, 5.027408, 5.04252, 5.063472, 5.091123, 5.125785, 5.16698, 
    5.213346, 5.262811, 5.313305, 5.359091, 5.398305, 5.430139, 5.45493, 
    5.475578, 5.491802, 5.50423, 5.510761, 5.511994, 5.507837, 5.49834, 
    5.482945, 5.46386, 5.440705, 5.414022, 5.381519, 5.343398, 5.300726, 
    5.255343, 5.209594, 5.165942, 5.126526, 5.092831, 5.06552, 5.044494, 
    5.029083, 5.018308, 5.011105, 5.006493, 5.003665, 5.002002, 5.00107, 
    5.000583,
  // height(7,49, 0-49)
    5.000078, 5.000158, 5.000323, 5.000648, 5.001265, 5.002378, 5.004317, 
    5.007565, 5.012781, 5.020815, 5.032668, 5.049388, 5.071904, 5.100811, 
    5.136148, 5.177304, 5.223419, 5.26947, 5.313471, 5.353898, 5.39002, 
    5.424407, 5.454918, 5.480593, 5.49589, 5.500593, 5.494115, 5.476953, 
    5.449314, 5.416775, 5.380487, 5.34278, 5.30167, 5.258408, 5.214767, 
    5.172745, 5.1342, 5.100561, 5.072627, 5.050539, 5.033884, 5.021892, 
    5.013636, 5.008191, 5.004746, 5.002652, 5.001432, 5.00075, 5.000383, 
    5.000201,
  // height(8,0, 0-49)
    5.001369, 5.00236, 5.004135, 5.007111, 5.011874, 5.019187, 5.02997, 
    5.045208, 5.065813, 5.092411, 5.125103, 5.163265, 5.205472, 5.249606, 
    5.293155, 5.333694, 5.369721, 5.397316, 5.416229, 5.42692, 5.430637, 
    5.429839, 5.425939, 5.420931, 5.415915, 5.412307, 5.410614, 5.410615, 
    5.41119, 5.411488, 5.409767, 5.404738, 5.39423, 5.377171, 5.353137, 
    5.322467, 5.286308, 5.246513, 5.205389, 5.165338, 5.128472, 5.096318, 
    5.069674, 5.048647, 5.032804, 5.021383, 5.013495, 5.008281, 5.005001, 
    5.003084,
  // height(8,1, 0-49)
    5.002229, 5.003803, 5.006566, 5.011106, 5.018226, 5.028921, 5.044301, 
    5.065442, 5.093146, 5.127659, 5.168413, 5.213895, 5.261753, 5.309123, 
    5.353121, 5.391528, 5.424201, 5.445468, 5.456513, 5.458668, 5.453891, 
    5.445782, 5.435674, 5.425931, 5.417472, 5.412071, 5.410341, 5.412109, 
    5.416037, 5.421542, 5.426564, 5.429821, 5.428074, 5.419613, 5.403261, 
    5.378569, 5.345982, 5.306887, 5.263489, 5.218513, 5.174774, 5.134702, 
    5.100015, 5.071559, 5.049369, 5.032875, 5.021171, 5.013241, 5.008139, 
    5.005085,
  // height(8,2, 0-49)
    5.003713, 5.006243, 5.010573, 5.017516, 5.028118, 5.043579, 5.065092, 
    5.093582, 5.12938, 5.171907, 5.219525, 5.269629, 5.319023, 5.3645, 
    5.403409, 5.434417, 5.459604, 5.47129, 5.472511, 5.465329, 5.452096, 
    5.437172, 5.421472, 5.407487, 5.395916, 5.388781, 5.386798, 5.389922, 
    5.39677, 5.407083, 5.418703, 5.430604, 5.438771, 5.441057, 5.435635, 
    5.421216, 5.397282, 5.364281, 5.323711, 5.278013, 5.230247, 5.183597, 
    5.140839, 5.103923, 5.073798, 5.050491, 5.033351, 5.021364, 5.013425, 
    5.008539,
  // height(8,3, 0-49)
    5.006076, 5.010056, 5.016683, 5.027022, 5.042336, 5.063916, 5.092799, 
    5.129389, 5.173098, 5.222139, 5.273632, 5.324032, 5.36979, 5.408006, 
    5.436888, 5.456504, 5.471837, 5.472431, 5.463517, 5.447612, 5.427128, 
    5.40682, 5.386859, 5.369648, 5.355633, 5.346969, 5.344492, 5.348353, 
    5.357283, 5.371386, 5.388593, 5.408371, 5.426187, 5.439701, 5.446662, 
    5.445097, 5.433551, 5.411355, 5.378881, 5.337667, 5.290347, 5.24031, 
    5.191145, 5.146004, 5.107107, 5.075537, 5.051323, 5.033752, 5.021726, 
    5.014085,
  // height(8,4, 0-49)
    5.009637, 5.015692, 5.025481, 5.040294, 5.061502, 5.09025, 5.127049, 
    5.171336, 5.221224, 5.273581, 5.324505, 5.370071, 5.407087, 5.433594, 
    5.449055, 5.455122, 5.460109, 5.449643, 5.431532, 5.408463, 5.382619, 
    5.358882, 5.336395, 5.317299, 5.301744, 5.291907, 5.288743, 5.292657, 
    5.302639, 5.319189, 5.340461, 5.366611, 5.392787, 5.416655, 5.435787, 
    5.447778, 5.450466, 5.442185, 5.42209, 5.39045, 5.348847, 5.300132, 
    5.24806, 5.196651, 5.149448, 5.108942, 5.07633, 5.051642, 5.034104, 
    5.022564,
  // height(8,5, 0-49)
    5.01475, 5.023616, 5.037497, 5.057807, 5.085801, 5.12212, 5.166306, 
    5.216456, 5.269265, 5.320505, 5.365861, 5.401783, 5.426079, 5.438101, 
    5.438597, 5.430701, 5.42629, 5.4058, 5.380095, 5.351824, 5.322756, 
    5.297715, 5.274599, 5.255134, 5.239125, 5.228632, 5.224696, 5.228026, 
    5.237998, 5.255537, 5.279135, 5.309788, 5.342454, 5.374955, 5.404862, 
    5.429592, 5.446565, 5.453413, 5.448264, 5.430104, 5.399138, 5.357038, 
    5.306925, 5.252957, 5.199602, 5.15078, 5.109215, 5.07619, 5.051716, 
    5.034968,
  // height(8,6, 0-49)
    5.021751, 5.034218, 5.053062, 5.079626, 5.114713, 5.158042, 5.207815, 
    5.260664, 5.312117, 5.35747, 5.39277, 5.415498, 5.424806, 5.421356, 
    5.406937, 5.385913, 5.373868, 5.3448, 5.313278, 5.281764, 5.251529, 
    5.227237, 5.205383, 5.187147, 5.171925, 5.161469, 5.156841, 5.159067, 
    5.168033, 5.185125, 5.209272, 5.242446, 5.279513, 5.318528, 5.357177, 
    5.392874, 5.422873, 5.444416, 5.454944, 5.452408, 5.435674, 5.404944, 
    5.362053, 5.310448, 5.254735, 5.199829, 5.15, 5.108155, 5.075609, 5.052327,
  // height(8,7, 0-49)
    5.03087, 5.047679, 5.07213, 5.105202, 5.146861, 5.19554, 5.247961, 
    5.299513, 5.345158, 5.38049, 5.402569, 5.410242, 5.403994, 5.385534, 
    5.357308, 5.324667, 5.306974, 5.270771, 5.235045, 5.202008, 5.172415, 
    5.150715, 5.131906, 5.116521, 5.103456, 5.093926, 5.088892, 5.089666, 
    5.096759, 5.112054, 5.135026, 5.168761, 5.208121, 5.251438, 5.296572, 
    5.341026, 5.38205, 5.416742, 5.442186, 5.45566, 5.454984, 5.438967, 
    5.407883, 5.363819, 5.310629, 5.253408, 5.197519, 5.147527, 5.106443, 
    5.075536,
  // height(8,8, 0-49)
    5.042141, 5.063857, 5.094147, 5.13329, 5.180078, 5.231492, 5.282947, 
    5.329145, 5.365218, 5.387711, 5.395039, 5.387403, 5.366355, 5.334259, 
    5.293848, 5.251297, 5.229727, 5.187588, 5.148976, 5.115803, 5.088339, 
    5.070806, 5.056664, 5.045733, 5.036299, 5.028781, 5.023865, 5.023066, 
    5.027584, 5.039847, 5.060001, 5.092403, 5.132013, 5.177479, 5.226856, 
    5.277767, 5.32753, 5.373251, 5.411896, 5.440407, 5.455941, 5.456232, 
    5.440107, 5.408016, 5.362398, 5.307615, 5.249297, 5.193226, 5.14417, 
    5.105097,
  // height(8,9, 0-49)
    5.055322, 5.08219, 5.118004, 5.162039, 5.21173, 5.262723, 5.309602, 
    5.347069, 5.371074, 5.379469, 5.372033, 5.35006, 5.315778, 5.271844, 
    5.22097, 5.170115, 5.145872, 5.098701, 5.058197, 5.025952, 5.0018, 
    4.989735, 4.981704, 4.976761, 4.972498, 4.968266, 4.964252, 4.962024, 
    4.963476, 4.971612, 4.987387, 5.016612, 5.05449, 5.100041, 5.151529, 
    5.206686, 5.262909, 5.317366, 5.367041, 5.408783, 5.439424, 5.456029, 
    5.456311, 5.439203, 5.405454, 5.357993, 5.301782, 5.243008, 5.187781, 
    5.140861,
  // height(8,10, 0-49)
    5.069841, 5.101693, 5.142138, 5.189268, 5.239218, 5.286673, 5.326009, 
    5.352551, 5.363453, 5.357918, 5.336849, 5.30226, 5.256696, 5.202795, 
    5.143048, 5.085224, 5.058656, 5.007109, 4.965445, 4.934928, 4.915015, 
    4.909478, 4.908812, 4.911294, 4.913756, 4.914239, 4.912184, 4.908985, 
    4.907153, 4.910244, 4.920147, 4.944366, 4.97854, 5.022159, 5.07372, 
    5.131052, 5.191589, 5.252552, 5.310984, 5.363772, 5.407672, 5.439425, 
    5.456047, 5.4553, 5.436343, 5.400368, 5.35093, 5.293661, 5.235225, 
    5.181823,
  // height(8,11, 0-49)
    5.084838, 5.121063, 5.164775, 5.212887, 5.260504, 5.301888, 5.331789, 
    5.346568, 5.34467, 5.326456, 5.293612, 5.248514, 5.193708, 5.13161, 
    5.064352, 5.000533, 4.970798, 4.915408, 4.873148, 4.844985, 4.83006, 
    4.831906, 4.839677, 4.850883, 4.861561, 4.868284, 4.869509, 4.866175, 
    4.861197, 4.858579, 4.861226, 4.878594, 4.907023, 4.946648, 4.996276, 
    5.053806, 5.116663, 5.182054, 5.247064, 5.308654, 5.363636, 5.408683, 
    5.44047, 5.45601, 5.453212, 5.431593, 5.392934, 5.341518, 5.283602, 
    5.226091,
  // height(8,12, 0-49)
    5.099267, 5.138888, 5.184268, 5.231308, 5.274516, 5.308251, 5.328059, 
    5.331479, 5.318122, 5.289199, 5.246833, 5.19346, 5.131418, 5.062748, 
    4.989133, 4.919843, 4.884488, 4.825829, 4.783488, 4.758223, 4.748928, 
    4.758839, 4.775925, 4.796943, 4.817178, 4.831673, 4.837736, 4.835538, 
    4.828052, 4.819459, 4.813668, 4.822335, 4.842855, 4.876289, 4.92189, 
    4.977654, 5.040928, 5.108822, 5.178389, 5.246644, 5.310491, 5.366675, 
    5.411796, 5.442484, 5.455814, 5.449941, 5.424872, 5.383087, 5.32959, 
    5.271071,
  // height(8,13, 0-49)
    5.112081, 5.153917, 5.199409, 5.243758, 5.281303, 5.306915, 5.317125, 
    5.310584, 5.287816, 5.250561, 5.201094, 5.141697, 5.07436, 5.000659, 
    4.921747, 4.846888, 4.801401, 4.740222, 4.698379, 4.676562, 4.673483, 
    4.691962, 4.719002, 4.750622, 4.781459, 4.80514, 4.817774, 4.818466, 
    4.809773, 4.795585, 4.780596, 4.77881, 4.789131, 4.813954, 4.853247, 
    4.905177, 4.966969, 5.035536, 5.107794, 5.180731, 5.25133, 5.316455, 
    5.372781, 5.41683, 5.445218, 5.455135, 5.445074, 5.415627, 5.37001, 
    5.313847,
  // height(8,14, 0-49)
    5.122416, 5.165294, 5.209671, 5.250387, 5.28198, 5.300036, 5.302077, 
    5.287667, 5.25795, 5.214927, 5.160814, 5.097618, 5.026911, 4.949761, 
    4.8667, 4.785186, 4.722669, 4.659978, 4.619365, 4.601606, 4.605288, 
    4.632604, 4.669907, 4.712483, 4.754512, 4.788497, 4.809477, 4.815284, 
    4.807504, 4.789055, 4.764913, 4.75128, 4.749103, 4.762674, 4.793109, 
    4.838937, 4.897255, 4.964674, 5.037851, 5.11364, 5.18903, 5.260995, 
    5.326344, 5.381658, 5.423375, 5.448099, 5.453174, 5.437504, 5.402347, 
    5.351675,
  // height(8,15, 0-49)
    5.129766, 5.172712, 5.215269, 5.252206, 5.278469, 5.290407, 5.286373, 
    5.266594, 5.232567, 5.18635, 5.129982, 5.065152, 4.993019, 4.914148, 
    4.828405, 4.73751, 4.64882, 4.585863, 4.547379, 4.534361, 4.545287, 
    4.581367, 4.628794, 4.682116, 4.735318, 4.780255, 4.811194, 4.824649, 
    4.820728, 4.800571, 4.768612, 4.74255, 4.725894, 4.725502, 4.744281, 
    4.781486, 4.83417, 4.898561, 4.970917, 5.047832, 5.126202, 5.203052, 
    5.275322, 5.339731, 5.392716, 5.430585, 5.449921, 5.448276, 5.425073, 
    5.382407,
  // height(8,16, 0-49)
    5.134052, 5.176439, 5.217067, 5.250836, 5.273164, 5.281045, 5.27343, 
    5.250941, 5.215213, 5.16822, 5.111789, 5.047322, 4.975654, 4.896925, 
    4.81037, 4.704902, 4.579583, 4.517775, 4.48243, 4.474857, 4.49339, 
    4.537728, 4.59462, 4.65787, 4.721575, 4.777524, 4.819635, 4.843246, 
    4.846655, 4.828532, 4.791764, 4.754059, 4.721835, 4.705099, 4.70937, 
    4.735244, 4.779961, 4.839344, 4.909132, 4.985513, 5.065176, 5.145107, 
    5.222342, 5.293738, 5.355831, 5.404837, 5.436883, 5.448555, 5.437765, 
    5.404779,
  // height(8,17, 0-49)
    5.13558, 5.177178, 5.216339, 5.248187, 5.268536, 5.274807, 5.266268, 
    5.243672, 5.208608, 5.162899, 5.108179, 5.045659, 4.975985, 4.899038, 
    4.813493, 4.685416, 4.513347, 4.454445, 4.423234, 4.421718, 4.448077, 
    4.499756, 4.565007, 4.636907, 4.70996, 4.776448, 4.830373, 4.866174, 
    4.880282, 4.868591, 4.831599, 4.784774, 4.737452, 4.702971, 4.690291, 
    4.702183, 4.736541, 4.78889, 4.854359, 4.928604, 5.007979, 5.08934, 
    5.169746, 5.246167, 5.315263, 5.37328, 5.416127, 5.43977, 5.440993, 
    5.418493,
  // height(8,18, 0-49)
    5.134904, 5.175833, 5.214426, 5.246045, 5.266733, 5.274041, 5.267223, 
    5.246889, 5.214422, 5.171445, 5.119457, 5.059613, 4.99252, 4.917845, 
    4.833514, 4.673349, 4.446044, 4.392892, 4.366827, 4.371818, 4.406159, 
    4.46414, 4.53652, 4.615712, 4.696862, 4.773158, 4.838974, 4.888155, 
    4.915483, 4.914273, 4.88238, 4.830496, 4.7705, 4.718554, 4.687547, 
    4.683339, 4.705169, 4.748554, 4.808033, 4.878636, 4.956275, 5.037578, 
    5.119546, 5.199218, 5.273369, 5.338331, 5.389959, 5.423878, 5.43611, 
    5.42413,
  // height(8,19, 0-49)
    5.132595, 5.173156, 5.21232, 5.245671, 5.269256, 5.280378, 5.277858, 
    5.261819, 5.23324, 5.193517, 5.144123, 5.086297, 5.020607, 4.946133, 
    4.858912, 4.659686, 4.369835, 4.327592, 4.308208, 4.320153, 4.362873, 
    4.426592, 4.505294, 4.590879, 4.679287, 4.764817, 4.84228, 4.905135, 
    4.946831, 4.958759, 4.936626, 4.884299, 4.815693, 4.74858, 4.699572, 
    4.678265, 4.686046, 4.71891, 4.770968, 4.836618, 4.91126, 4.991214, 
    5.073359, 5.154741, 5.232225, 5.30225, 5.360712, 5.4031, 5.424982, 
    5.422957,
  // height(8,20, 0-49)
    5.126199, 5.16312, 5.199585, 5.231456, 5.255075, 5.268044, 5.269554, 
    5.260229, 5.241733, 5.216325, 5.186499, 5.154742, 5.123319, 5.093983, 
    5.067405, 0, 4.110707, 4.123703, 4.162252, 4.22343, 4.302578, 4.387699, 
    4.480834, 4.576489, 4.673163, 4.767192, 4.854263, 4.927924, 4.980938, 
    5.003913, 4.991771, 4.940973, 4.867107, 4.788014, 4.72289, 4.684924, 
    4.678152, 4.699588, 4.743227, 4.802933, 4.873587, 4.951164, 5.032368, 
    5.114204, 5.193589, 5.267064, 5.330619, 5.379736, 5.409759, 5.416706,
  // height(8,21, 0-49)
    5.123293, 5.160292, 5.19839, 5.233569, 5.261959, 5.280674, 5.288291, 
    5.284894, 5.271763, 5.25098, 5.225037, 5.196559, 5.168098, 5.141923, 
    5.119676, 0, 4.030297, 4.047019, 4.093606, 4.164876, 4.254046, 4.343937, 
    4.441362, 4.540665, 4.641256, 4.74086, 4.835884, 4.920084, 4.985749, 
    5.023064, 5.026696, 4.98524, 4.915319, 4.832731, 4.757448, 4.705839, 
    4.685367, 4.695097, 4.729599, 4.782505, 4.848262, 4.922476, 5.001632, 
    5.082644, 5.162446, 5.237658, 5.304375, 5.358139, 5.394198, 5.408191,
  // height(8,22, 0-49)
    5.121522, 5.158882, 5.19856, 5.236558, 5.268754, 5.291821, 5.30385, 
    5.304541, 5.29497, 5.277183, 5.253765, 5.227507, 5.201188, 5.177412, 
    5.158434, 0, 3.962537, 3.984438, 4.038232, 4.117738, 4.215069, 4.308348, 
    4.409274, 4.511858, 4.616008, 4.720365, 4.821665, 4.913651, 4.988194, 
    5.035557, 5.051208, 5.016985, 4.95165, 4.868662, 4.787441, 4.726087, 
    4.694775, 4.694649, 4.721154, 4.767963, 4.829233, 4.900268, 4.97734, 
    5.057264, 5.136958, 5.2131, 5.281876, 5.338915, 5.379454, 5.398909,
  // height(8,23, 0-49)
    5.120916, 5.158588, 5.199337, 5.239162, 5.273767, 5.299524, 5.314222, 
    5.31733, 5.309831, 5.293787, 5.271873, 5.247006, 5.222109, 5.199984, 
    5.183231, 0, 3.917093, 3.943388, 4.002137, 4.086914, 4.189435, 4.283938, 
    4.386425, 4.49054, 4.59648, 4.703573, 4.808774, 4.905783, 4.986151, 
    5.040359, 5.064946, 5.036311, 4.975649, 4.894337, 4.810658, 4.743364, 
    4.704498, 4.696982, 4.71723, 4.759143, 4.816749, 4.885137, 4.960407, 
    5.039274, 5.118623, 5.195158, 5.265129, 5.324236, 5.367732, 5.390903,
  // height(8,24, 0-49)
    5.121484, 5.15919, 5.200179, 5.240473, 5.275757, 5.302342, 5.317935, 
    5.321938, 5.315293, 5.30006, 5.278937, 5.254865, 5.230805, 5.209631, 
    5.194072, 0, 3.898081, 3.926662, 3.987599, 4.074533, 4.179204, 4.273223, 
    4.375597, 4.479658, 4.58575, 4.69365, 4.800478, 4.89992, 4.983319, 
    5.04135, 5.071414, 5.046269, 4.989053, 4.909707, 4.825484, 4.755218, 
    4.711973, 4.699844, 4.715989, 4.754571, 4.8096, 4.876063, 4.949962, 
    5.027952, 5.106898, 5.183519, 5.254107, 5.31441, 5.359709, 5.385231,
  // height(8,25, 0-49)
    5.12319, 5.160546, 5.200797, 5.240048, 5.274151, 5.299625, 5.314344, 
    5.317798, 5.31093, 5.295742, 5.274842, 5.251086, 5.227356, 5.206459, 
    5.191058, 0, 3.905595, 3.934001, 3.99451, 4.080811, 4.184822, 4.277218, 
    4.378278, 4.481149, 4.586186, 4.693312, 4.799687, 4.89899, 4.982497, 
    5.040989, 5.072271, 5.047817, 4.991623, 4.913149, 4.829183, 4.758409, 
    4.714091, 4.70067, 4.715574, 4.753094, 4.807269, 4.873075, 4.946495, 
    5.024164, 5.102949, 5.179572, 5.250342, 5.311027, 5.356915, 5.383218,
  // height(8,26, 0-49)
    5.125965, 5.16261, 5.201203, 5.237979, 5.269135, 5.291635, 5.303749, 
    5.305204, 5.296997, 5.28103, 5.259737, 5.235774, 5.211836, 5.190529, 
    5.174261, 0, 3.937386, 3.963501, 4.021425, 4.104737, 4.20558, 4.295581, 
    4.394385, 4.495152, 4.598157, 4.703125, 4.807133, 4.903847, 4.984638, 
    5.040278, 5.0684, 5.04177, 4.983876, 4.904703, 4.821317, 4.752176, 
    4.709991, 4.698662, 4.715331, 4.75422, 4.809419, 4.87597, 4.949917, 
    5.027929, 5.106887, 5.183514, 5.254105, 5.314409, 5.359708, 5.385231,
  // height(8,27, 0-49)
    5.129717, 5.165435, 5.201689, 5.23486, 5.261594, 5.279465, 5.287314, 
    5.285252, 5.274403, 5.256595, 5.234052, 5.209174, 5.184377, 5.16194, 
    5.143804, 0, 3.989284, 4.01185, 4.065571, 4.143941, 4.239443, 4.326462, 
    4.422174, 4.519982, 4.619985, 4.72141, 4.821146, 4.912863, 4.98817, 
    5.037752, 5.058598, 5.027196, 4.965382, 4.884583, 4.802653, 4.737598, 
    4.700779, 4.694783, 4.716008, 4.758492, 4.81641, 4.884964, 4.96032, 
    5.03923, 5.118601, 5.195146, 5.265124, 5.324234, 5.36773, 5.390903,
  // height(8,28, 0-49)
    5.134365, 5.169187, 5.202791, 5.231663, 5.252913, 5.264796, 5.266833, 
    5.25964, 5.244601, 5.223562, 5.198596, 5.171845, 5.145388, 5.121049, 
    5.100052, 0, 4.056873, 4.075941, 4.124346, 4.195992, 4.284093, 4.367258, 
    4.458745, 4.55243, 4.648153, 4.744445, 4.837958, 4.922404, 4.989758, 
    5.030591, 5.041007, 5.003144, 4.936561, 4.854705, 4.776264, 4.7182, 
    4.689766, 4.691714, 4.719532, 4.767098, 4.828782, 4.900036, 4.977222, 
    5.057204, 5.136929, 5.213084, 5.281867, 5.338911, 5.379453, 5.398908,
  // height(8,29, 0-49)
    5.139871, 5.174164, 5.205247, 5.229603, 5.244735, 5.249564, 5.244349, 
    5.230343, 5.209353, 5.183419, 5.154596, 5.124834, 5.095839, 5.068839, 
    5.043989, 0, 4.134919, 4.152247, 4.194923, 4.258248, 4.336938, 4.414831, 
    4.500596, 4.588754, 4.67878, 4.768302, 4.853632, 4.928486, 4.985303, 
    5.014688, 5.012098, 4.966738, 4.896005, 4.815494, 4.744064, 4.696627, 
    4.679617, 4.691761, 4.727758, 4.781523, 4.847747, 4.922211, 5.001495, 
    5.082574, 5.16241, 5.23764, 5.304365, 5.358133, 5.394195, 5.408189,
  // height(8,30, 0-49)
    5.149293, 5.187366, 5.220729, 5.245617, 5.259345, 5.260664, 5.249608, 
    5.227057, 5.194283, 5.152627, 5.103288, 5.047123, 4.984291, 4.913467, 
    4.830404, 4.635087, 4.366791, 4.33845, 4.330659, 4.350416, 4.397135, 
    4.457949, 4.533136, 4.614896, 4.700094, 4.78401, 4.861721, 4.926516, 
    4.971288, 4.987126, 4.969789, 4.916682, 4.843794, 4.76844, 4.708371, 
    4.675247, 4.67223, 4.696182, 4.74135, 4.801925, 4.873054, 4.950885, 
    5.032222, 5.114128, 5.19355, 5.267044, 5.330608, 5.37973, 5.409755, 
    5.416704,
  // height(8,31, 0-49)
    5.154108, 5.192601, 5.225134, 5.247748, 5.25784, 5.254495, 5.238242, 
    5.21049, 5.172945, 5.127208, 5.074561, 5.015869, 4.951433, 4.880641, 
    4.801196, 4.644937, 4.432422, 4.392949, 4.379121, 4.393623, 4.43407, 
    4.491832, 4.56249, 4.638905, 4.717442, 4.792549, 4.859183, 4.911111, 
    4.942367, 4.945229, 4.916481, 4.861229, 4.793419, 4.729975, 4.685867, 
    4.669163, 4.680465, 4.715677, 4.769167, 4.835639, 4.910736, 4.990936, 
    5.073214, 5.154664, 5.232185, 5.30223, 5.360701, 5.403094, 5.424978, 
    5.422956,
  // height(8,32, 0-49)
    5.157407, 5.197023, 5.230282, 5.252917, 5.262111, 5.256892, 5.237898, 
    5.206759, 5.165463, 5.115866, 5.059437, 4.997152, 4.929425, 4.855934, 
    4.775219, 4.651386, 4.489683, 4.443143, 4.423618, 4.431955, 4.465497, 
    4.519353, 4.584921, 4.655719, 4.727498, 4.793783, 4.849238, 4.888139, 
    4.905953, 4.896959, 4.860013, 4.806783, 4.748804, 4.70111, 4.675007, 
    4.67511, 4.700132, 4.745621, 4.806382, 4.877728, 4.955783, 5.037313, 
    5.119405, 5.199143, 5.273329, 5.33831, 5.389947, 5.423872, 5.436106, 
    5.424129,
  // height(8,33, 0-49)
    5.158516, 5.199754, 5.23505, 5.259749, 5.270575, 5.266178, 5.24701, 
    5.214706, 5.171402, 5.119178, 5.05975, 4.994316, 4.923507, 4.847308, 
    4.764863, 4.663693, 4.545833, 4.494422, 4.469296, 4.470886, 4.496832, 
    4.54519, 4.604345, 4.668429, 4.732591, 4.78956, 4.833763, 4.860198, 
    4.866086, 4.848289, 4.808124, 4.76158, 4.717298, 4.687345, 4.679305, 
    4.695044, 4.732172, 4.786329, 4.852901, 4.927793, 5.007535, 5.089099, 
    5.169616, 5.246097, 5.315227, 5.37326, 5.416117, 5.439764, 5.44099, 
    5.418491,
  // height(8,34, 0-49)
    5.156674, 5.199654, 5.237898, 5.26634, 5.281066, 5.280095, 5.263408, 
    5.232435, 5.189331, 5.136365, 5.075525, 5.008317, 4.935713, 4.858127, 
    4.77535, 4.688264, 4.605028, 4.550157, 4.519898, 4.514716, 4.532631, 
    4.573838, 4.625031, 4.68093, 4.736253, 4.78332, 4.816595, 4.832085, 
    4.828914, 4.806611, 4.768563, 4.732501, 4.703937, 4.691649, 4.700083, 
    4.72925, 4.776286, 4.837176, 4.907887, 4.984814, 5.064787, 5.144894, 
    5.222227, 5.293676, 5.355797, 5.404819, 5.436873, 5.448549, 5.437762, 
    5.404777,
  // height(8,35, 0-49)
    5.151281, 5.195655, 5.237204, 5.270538, 5.291034, 5.29586, 5.284276, 
    5.257265, 5.216847, 5.165399, 5.10517, 5.038023, 4.965342, 4.888039, 
    4.806555, 4.727874, 4.66922, 4.612257, 4.577751, 4.566242, 4.576077, 
    4.608909, 4.650864, 4.69726, 4.742668, 4.779547, 4.802795, 4.809654, 
    4.800983, 4.778551, 4.746922, 4.72342, 4.710607, 4.714301, 4.736648, 
    4.776581, 4.831155, 4.89677, 4.969879, 5.047243, 5.125873, 5.202868, 
    5.275223, 5.339676, 5.392687, 5.430571, 5.449914, 5.448271, 5.425071, 
    5.382406,
  // height(8,36, 0-49)
    5.142104, 5.187049, 5.231609, 5.270293, 5.297827, 5.310411, 5.306343, 
    5.285905, 5.250766, 5.203276, 5.145887, 5.080808, 5.009852, 4.934427, 
    4.85556, 4.782229, 4.739129, 4.681488, 4.643786, 4.626654, 4.628716, 
    4.652565, 4.684572, 4.720676, 4.75562, 4.782554, 4.797193, 4.798059, 
    4.787327, 4.768233, 4.745573, 4.734941, 4.736442, 4.753576, 4.786968, 
    4.834998, 4.894826, 4.963222, 5.037002, 5.113153, 5.188756, 5.260842, 
    5.326259, 5.381612, 5.423351, 5.448085, 5.453167, 5.4375, 5.402345, 
    5.351675,
  // height(8,37, 0-49)
    5.129393, 5.173698, 5.220318, 5.263993, 5.299031, 5.320687, 5.326133, 
    5.314678, 5.287379, 5.246348, 5.194114, 5.133163, 5.065706, 4.993609, 
    4.918402, 4.849136, 4.814672, 4.757637, 4.717738, 4.695762, 4.690593, 
    4.705426, 4.727391, 4.753076, 4.777669, 4.795451, 4.803186, 4.800547, 
    4.790458, 4.776838, 4.763995, 4.765265, 4.778885, 4.806695, 4.848376, 
    4.902049, 4.965028, 5.034365, 5.107103, 5.18033, 5.251101, 5.316327, 
    5.372707, 5.41679, 5.445196, 5.455124, 5.445068, 5.415625, 5.370009, 
    5.313847,
  // height(8,38, 0-49)
    5.113876, 5.156118, 5.203286, 5.250753, 5.292802, 5.323964, 5.340252, 
    5.339784, 5.322693, 5.290582, 5.245847, 5.191123, 5.128939, 5.06156, 
    4.990949, 4.92551, 4.895123, 4.839703, 4.798448, 4.772382, 4.760661, 
    4.766866, 4.779205, 4.794943, 4.809895, 4.819722, 4.822293, 4.81818, 
    4.810492, 4.803233, 4.799835, 4.811351, 4.83469, 4.870549, 4.918038, 
    4.975163, 5.039362, 5.107861, 5.17781, 5.2463, 5.31029, 5.36656, 
    5.411729, 5.442446, 5.455794, 5.449931, 5.424867, 5.383084, 5.329588, 
    5.27107,
  // height(8,39, 0-49)
    5.096656, 5.135428, 5.181291, 5.230628, 5.278194, 5.318223, 5.345743, 
    5.35758, 5.352668, 5.331766, 5.29685, 5.250499, 5.195425, 5.134211, 
    5.069193, 5.00797, 4.979156, 4.926097, 4.884192, 4.854754, 4.837235, 
    4.835485, 4.838983, 4.845691, 4.852136, 4.855419, 4.85442, 4.850298, 
    4.845923, 4.844999, 4.849974, 4.869821, 4.900551, 4.94209, 4.99318, 
    5.051761, 5.115341, 5.181213, 5.246534, 5.308325, 5.363435, 5.408561, 
    5.440397, 5.455967, 5.453187, 5.43158, 5.392928, 5.341514, 5.283599, 
    5.22609,
  // height(8,40, 0-49)
    5.079001, 5.113148, 5.155824, 5.20466, 5.255383, 5.302495, 5.340465, 
    5.364939, 5.373489, 5.365705, 5.342792, 5.306976, 5.260952, 5.2075, 
    5.149253, 5.093055, 5.064897, 5.0148, 4.972912, 4.940837, 4.918354, 
    4.909531, 4.905233, 4.904131, 4.903456, 4.901661, 4.898442, 4.895254, 
    4.894445, 4.899253, 4.911187, 4.93741, 4.973363, 5.018431, 5.071098, 
    5.129232, 5.190343, 5.251703, 5.310411, 5.363389, 5.407419, 5.439262, 
    5.455943, 5.455236, 5.436306, 5.400346, 5.350918, 5.293653, 5.235221, 
    5.181822,
  // height(8,41, 0-49)
    5.062121, 5.090923, 5.128824, 5.174737, 5.225716, 5.277128, 5.323496, 
    5.359679, 5.381943, 5.388488, 5.379393, 5.356171, 5.321213, 5.27729, 
    5.227234, 5.177218, 5.149961, 5.103456, 5.062327, 5.028457, 5.001982, 
    4.98717, 4.976339, 4.968845, 4.962564, 4.957095, 4.952728, 4.950969, 
    4.953513, 4.963099, 4.980418, 5.011087, 5.050213, 5.096777, 5.149055, 
    5.204819, 5.261506, 5.316321, 5.366274, 5.40823, 5.439034, 5.455762, 
    5.456133, 5.439089, 5.405383, 5.35795, 5.301758, 5.242993, 5.187772, 
    5.140857,
  // height(8,42, 0-49)
    5.046977, 5.07022, 5.102299, 5.143245, 5.191529, 5.243844, 5.29543, 
    5.341003, 5.375879, 5.396879, 5.402698, 5.393766, 5.371802, 5.339299, 
    5.299088, 5.256725, 5.231469, 5.189376, 5.149957, 5.115338, 5.086065, 
    5.066585, 5.050688, 5.038368, 5.028037, 5.02018, 5.015453, 5.015247, 
    5.020588, 5.033757, 5.054786, 5.087964, 5.128242, 5.174273, 5.224139, 
    5.275482, 5.32564, 5.371724, 5.410694, 5.439491, 5.455265, 5.455751, 
    5.439777, 5.407797, 5.36226, 5.307529, 5.249246, 5.193198, 5.144154, 
    5.105088,
  // height(8,43, 0-49)
    5.034163, 5.052107, 5.077977, 5.1126, 5.155713, 5.205489, 5.25843, 
    5.309834, 5.354713, 5.388844, 5.409515, 5.415804, 5.408386, 5.389111, 
    5.360541, 5.327561, 5.306041, 5.269506, 5.233062, 5.199059, 5.168477, 
    5.145934, 5.126657, 5.111196, 5.098354, 5.089241, 5.084676, 5.085835, 
    5.093141, 5.108504, 5.131452, 5.165137, 5.204473, 5.247838, 5.293118, 
    5.337825, 5.379192, 5.41429, 5.440164, 5.454059, 5.453766, 5.438076, 
    5.407258, 5.363396, 5.310354, 5.253236, 5.197416, 5.147466, 5.106408, 
    5.075515,
  // height(8,44, 0-49)
    5.023893, 5.037152, 5.057038, 5.08481, 5.121122, 5.165492, 5.215907, 
    5.268845, 5.319784, 5.364102, 5.398016, 5.419214, 5.427063, 5.422406, 
    5.407182, 5.385447, 5.369846, 5.3404, 5.308588, 5.276946, 5.246899, 
    5.223215, 5.202463, 5.185639, 5.171791, 5.162381, 5.15825, 5.160318, 
    5.168521, 5.184505, 5.207436, 5.239498, 5.275653, 5.314039, 5.352384, 
    5.388091, 5.418369, 5.440388, 5.451512, 5.449613, 5.433495, 5.403317, 
    5.360887, 5.309646, 5.254205, 5.199492, 5.149795, 5.108033, 5.075538, 
    5.052284,
  // height(8,45, 0-49)
    5.016068, 5.025445, 5.040023, 5.06117, 5.090047, 5.127151, 5.171838, 
    5.22204, 5.274341, 5.324514, 5.368355, 5.402508, 5.425014, 5.435463, 
    5.434813, 5.426049, 5.418765, 5.398278, 5.373139, 5.345995, 5.318683, 
    5.296079, 5.275944, 5.259601, 5.246169, 5.237257, 5.233617, 5.23592, 
    5.243749, 5.258614, 5.279437, 5.307597, 5.338169, 5.369109, 5.398049, 
    5.4224, 5.439507, 5.446893, 5.442554, 5.425341, 5.395344, 5.354149, 
    5.304817, 5.251482, 5.198609, 5.150136, 5.108815, 5.075948, 5.051572, 
    5.034879,
  // height(8,46, 0-49)
    5.010371, 5.016713, 5.026895, 5.042174, 5.063859, 5.092983, 5.129908, 
    5.173916, 5.222999, 5.273985, 5.323053, 5.366474, 5.401325, 5.425965, 
    5.440145, 5.44553, 5.448809, 5.439283, 5.423095, 5.402858, 5.380724, 
    5.361625, 5.344312, 5.33029, 5.318596, 5.310812, 5.307542, 5.309251, 
    5.315293, 5.327178, 5.343702, 5.365603, 5.388121, 5.409129, 5.4263, 
    5.437255, 5.439753, 5.431987, 5.41292, 5.382617, 5.342471, 5.295172, 
    5.244368, 5.194016, 5.147643, 5.107752, 5.075573, 5.051174, 5.03382, 
    5.022387,
  // height(8,47, 0-49)
    5.006379, 5.010458, 5.017199, 5.027631, 5.042955, 5.064367, 5.092776, 
    5.128459, 5.170724, 5.217763, 5.2668, 5.314528, 5.357748, 5.393965, 
    5.421778, 5.441412, 5.456867, 5.46001, 5.454927, 5.44398, 5.429455, 
    5.416289, 5.403948, 5.393989, 5.385193, 5.379011, 5.375869, 5.37608, 
    5.378881, 5.385936, 5.396016, 5.409431, 5.421616, 5.430514, 5.434071, 
    5.430398, 5.418005, 5.396079, 5.364757, 5.325294, 5.280035, 5.23211, 
    5.184909, 5.141459, 5.10393, 5.073397, 5.049934, 5.032877, 5.021182, 
    5.013739,
  // height(8,48, 0-49)
    5.003644, 5.006086, 5.010241, 5.016864, 5.02692, 5.041507, 5.061704, 
    5.088339, 5.121694, 5.161249, 5.20556, 5.252367, 5.298956, 5.342635, 
    5.381233, 5.413701, 5.441738, 5.458355, 5.465828, 5.466006, 5.46107, 
    5.455938, 5.450424, 5.446013, 5.441033, 5.436764, 5.433451, 5.431307, 
    5.42953, 5.430123, 5.431936, 5.435133, 5.435347, 5.430807, 5.42, 
    5.401847, 5.375895, 5.342507, 5.302944, 5.259302, 5.21424, 5.17055, 
    5.13068, 5.096348, 5.068379, 5.046762, 5.030877, 5.019772, 5.012416, 
    5.007883,
  // height(8,49, 0-49)
    5.001472, 5.002565, 5.00451, 5.007768, 5.012981, 5.020984, 5.032765, 
    5.049376, 5.071753, 5.100489, 5.135601, 5.176348, 5.22122, 5.268123, 
    5.314735, 5.359285, 5.403051, 5.435205, 5.457379, 5.470873, 5.477746, 
    5.48514, 5.4914, 5.497845, 5.49962, 5.498258, 5.49363, 5.486034, 
    5.474223, 5.463232, 5.452115, 5.442515, 5.428285, 5.40822, 5.38172, 
    5.348891, 5.31062, 5.268536, 5.22482, 5.181884, 5.141978, 5.106841, 
    5.077487, 5.054176, 5.036537, 5.023789, 5.01498, 5.009157, 5.005493, 
    5.003342,
  // height(9,0, 0-49)
    5.013042, 5.019694, 5.029954, 5.044734, 5.064919, 5.091146, 5.123545, 
    5.161498, 5.203522, 5.247341, 5.290179, 5.329203, 5.361989, 5.386886, 
    5.403194, 5.411325, 5.413615, 5.407965, 5.397056, 5.382667, 5.366389, 
    5.350346, 5.335258, 5.322433, 5.312547, 5.306667, 5.305348, 5.308775, 
    5.316498, 5.328191, 5.342663, 5.358954, 5.37482, 5.38847, 5.398046, 
    5.401766, 5.398109, 5.386037, 5.365193, 5.336077, 5.300086, 5.259408, 
    5.216734, 5.174833, 5.136135, 5.102393, 5.074556, 5.052821, 5.03683, 
    5.025922,
  // height(9,1, 0-49)
    5.018539, 5.027684, 5.041417, 5.060682, 5.086233, 5.118349, 5.15655, 
    5.19942, 5.244636, 5.289235, 5.330095, 5.364451, 5.390327, 5.406764, 
    5.413841, 5.412899, 5.408258, 5.395083, 5.37753, 5.357601, 5.33689, 
    5.31798, 5.300873, 5.28678, 5.275898, 5.269395, 5.267859, 5.271605, 
    5.28021, 5.293866, 5.31147, 5.332596, 5.354544, 5.375515, 5.393538, 
    5.406585, 5.412741, 5.410409, 5.398545, 5.376884, 5.346107, 5.307889, 
    5.264752, 5.219728, 5.175877, 5.135812, 5.10137, 5.073483, 5.052285, 
    5.037354,
  // height(9,2, 0-49)
    5.026684, 5.039216, 5.057403, 5.082047, 5.113499, 5.151348, 5.194202, 
    5.239692, 5.284729, 5.326012, 5.360569, 5.386237, 5.401902, 5.407519, 
    5.403984, 5.393466, 5.38223, 5.362339, 5.339471, 5.315671, 5.292365, 
    5.272373, 5.254879, 5.240854, 5.229998, 5.223449, 5.221773, 5.225418, 
    5.234077, 5.248452, 5.26766, 5.291913, 5.318253, 5.345037, 5.370354, 
    5.392126, 5.40825, 5.416761, 5.416035, 5.405025, 5.383495, 5.35221, 
    5.312987, 5.268557, 5.222194, 5.177207, 5.136419, 5.101797, 5.074339, 
    5.054193,
  // height(9,3, 0-49)
    5.037796, 5.054545, 5.077931, 5.108358, 5.145469, 5.18788, 5.233158, 
    5.278073, 5.319133, 5.353187, 5.377922, 5.392138, 5.395739, 5.389587, 
    5.375238, 5.355539, 5.338708, 5.313167, 5.286374, 5.260293, 5.236083, 
    5.216662, 5.200305, 5.187636, 5.177845, 5.171894, 5.170265, 5.173514, 
    5.181518, 5.195473, 5.21482, 5.240509, 5.269487, 5.300368, 5.331426, 
    5.360679, 5.385998, 5.405237, 5.416381, 5.417744, 5.408212, 5.3875, 
    5.356378, 5.316756, 5.271558, 5.224334, 5.17869, 5.137706, 5.103526, 
    5.07722,
  // height(9,4, 0-49)
    5.052035, 5.073641, 5.102532, 5.138441, 5.180034, 5.224841, 5.269492, 
    5.310276, 5.3438, 5.367561, 5.380238, 5.381697, 5.372798, 5.355103, 
    5.330607, 5.30267, 5.281563, 5.251438, 5.221951, 5.194925, 5.171211, 
    5.153751, 5.139843, 5.129701, 5.121983, 5.117336, 5.116074, 5.11881, 
    5.125641, 5.138234, 5.156425, 5.182015, 5.211965, 5.245227, 5.280334, 
    5.31548, 5.34862, 5.37757, 5.400111, 5.414134, 5.417838, 5.409997, 
    5.390258, 5.359409, 5.319504, 5.273733, 5.225988, 5.18022, 5.139762, 
    5.106874,
  // height(9,5, 0-49)
    5.06927, 5.096024, 5.130133, 5.170412, 5.21444, 5.258764, 5.299453, 
    5.332823, 5.356091, 5.367723, 5.367478, 5.356185, 5.335419, 5.307194, 
    5.273708, 5.238726, 5.214715, 5.180921, 5.149723, 5.122785, 5.100636, 
    5.086227, 5.075836, 5.069233, 5.064543, 5.061961, 5.061525, 5.063834, 
    5.069201, 5.079716, 5.095667, 5.119814, 5.149218, 5.18323, 5.220694, 
    5.260019, 5.299302, 5.336403, 5.369049, 5.394906, 5.411742, 5.417627, 
    5.411244, 5.392218, 5.361438, 5.321201, 5.275047, 5.227249, 5.182064, 
    5.142961,
  // height(9,6, 0-49)
    5.088974, 5.120697, 5.159075, 5.201886, 5.245714, 5.28647, 5.320168, 
    5.343662, 5.355105, 5.354039, 5.341181, 5.318075, 5.28674, 5.249392, 
    5.208251, 5.167442, 5.141766, 5.105011, 5.072841, 5.046739, 5.026933, 
    5.016384, 5.01034, 5.008129, 5.007359, 5.007643, 5.008629, 5.010802, 
    5.014644, 5.022597, 5.035425, 5.056958, 5.084433, 5.117664, 5.155847, 
    5.197634, 5.241279, 5.284737, 5.325753, 5.361929, 5.390816, 5.410064, 
    5.417652, 5.412226, 5.393486, 5.362525, 5.321963, 5.275724, 5.22841, 
    5.184418,
  // height(9,7, 0-49)
    5.110209, 5.146196, 5.187303, 5.230341, 5.2712, 5.305634, 5.330105, 
    5.342353, 5.341588, 5.328314, 5.30397, 5.270539, 5.230231, 5.185272, 
    5.137776, 5.092242, 5.065883, 5.026673, 4.994061, 4.969322, 4.952398, 
    4.94629, 4.94522, 4.948102, 4.952066, 4.956038, 4.959166, 4.961686, 
    4.96418, 4.969313, 4.978322, 4.996211, 5.020468, 5.051454, 5.088767, 
    5.131334, 5.177573, 5.225541, 5.273042, 5.317697, 5.356995, 5.388387, 
    5.409444, 5.418111, 5.413079, 5.394205, 5.362855, 5.321998, 5.275874, 
    5.22923,
  // height(9,8, 0-49)
    5.131696, 5.170769, 5.212703, 5.253581, 5.289032, 5.315145, 5.329186, 
    5.329929, 5.317555, 5.293313, 5.25909, 5.217057, 5.16942, 5.118283, 
    5.06558, 5.016235, 4.989789, 4.94848, 4.915803, 4.892795, 4.879127, 
    4.877858, 4.882214, 4.890742, 4.900167, 4.908644, 4.914731, 4.918277, 
    4.919837, 4.922133, 4.926813, 4.940151, 4.959956, 4.987245, 5.022112, 
    5.063804, 5.110915, 5.161597, 5.213713, 5.264927, 5.312754, 5.354599, 
    5.387856, 5.410053, 5.419156, 5.413955, 5.394502, 5.362439, 5.321009, 
    5.274606,
  // height(9,9, 0-49)
    5.152001, 5.192673, 5.233472, 5.270114, 5.29842, 5.315174, 5.318628, 
    5.308538, 5.285864, 5.252336, 5.21005, 5.161165, 5.107756, 5.051719, 
    4.994766, 4.942291, 4.915819, 4.872682, 4.84023, 4.81922, 4.809059, 
    4.812881, 4.822952, 4.837524, 4.85301, 4.866771, 4.876707, 4.882144, 
    4.883457, 4.883184, 4.883249, 4.891264, 4.905428, 4.927546, 4.95835, 
    4.997493, 5.043778, 5.095445, 5.150386, 5.2063, 5.260748, 5.311169, 
    5.354927, 5.389367, 5.412012, 5.420855, 5.414785, 5.39402, 5.360405, 
    5.317352,
  // height(9,10, 0-49)
    5.169785, 5.210491, 5.248452, 5.279398, 5.299693, 5.307023, 5.300615, 
    5.281043, 5.249805, 5.208882, 5.160379, 5.106323, 5.048559, 4.988734, 
    4.928304, 4.873112, 4.845929, 4.801261, 4.769295, 4.750492, 4.743991, 
    4.753007, 4.768904, 4.789725, 4.811697, 4.831421, 4.846126, 4.854508, 
    4.856575, 4.854371, 4.849869, 4.852006, 4.859412, 4.874855, 4.899894, 
    4.934735, 4.978467, 5.029416, 5.085478, 5.144336, 5.203576, 5.260691, 
    5.313084, 5.358071, 5.392953, 5.41521, 5.422825, 5.414724, 5.391241, 
    5.354405,
  // height(9,11, 0-49)
    5.184051, 5.223395, 5.257313, 5.281863, 5.294163, 5.292828, 5.27793, 
    5.25065, 5.212797, 5.166412, 5.113485, 5.055821, 4.994998, 4.932372, 
    4.869107, 4.811265, 4.781673, 4.735917, 4.704734, 4.688303, 4.685516, 
    4.699636, 4.72124, 4.748251, 4.776879, 4.803067, 4.823434, 4.835981, 
    4.840165, 4.837159, 4.828632, 4.824708, 4.824437, 4.831717, 4.849192, 
    4.877854, 4.917208, 4.965708, 5.021219, 5.081358, 5.143673, 5.205681, 
    5.264839, 5.318503, 5.363908, 5.398248, 5.41888, 5.423704, 5.411665, 
    5.383304,
  // height(9,12, 0-49)
    5.194335, 5.231282, 5.260574, 5.278791, 5.28386, 5.275225, 5.253618, 
    5.220604, 5.178126, 5.128154, 5.072487, 5.012671, 4.949991, 4.885493, 
    4.82, 4.759103, 4.724104, 4.677974, 4.647959, 4.634027, 4.634865, 
    4.653734, 4.680614, 4.713413, 4.74852, 4.781399, 4.808202, 4.826231, 
    4.834251, 4.832163, 4.82086, 4.811296, 4.802845, 4.800652, 4.808741, 
    4.829211, 4.862217, 4.906439, 4.959705, 5.019504, 5.083271, 5.148478, 
    5.212607, 5.273064, 5.327098, 5.371778, 5.404087, 5.421196, 5.420952, 
    5.402519,
  // height(9,13, 0-49)
    5.20077, 5.234771, 5.259482, 5.27208, 5.271227, 5.25703, 5.230669, 
    5.19392, 5.148717, 5.09689, 5.04002, 4.97939, 4.916002, 4.850582, 
    4.783556, 4.718486, 4.673654, 4.628222, 4.599886, 4.588519, 4.592689, 
    4.615596, 4.646937, 4.684716, 4.725712, 4.765153, 4.798926, 4.823727, 
    4.837541, 4.838665, 4.826695, 4.812769, 4.796377, 4.783873, 4.780921, 
    4.791139, 4.815689, 4.853671, 4.902922, 4.960753, 5.024401, 5.091208, 
    5.158616, 5.22405, 5.284799, 5.337901, 5.380161, 5.408309, 5.419418, 
    5.411558,
  // height(9,14, 0-49)
    5.204044, 5.235059, 5.255784, 5.26395, 5.258807, 5.240928, 5.211757, 
    5.173126, 5.126891, 5.074712, 5.01796, 4.9577, 4.894693, 4.829371, 
    4.761736, 4.690343, 4.630024, 4.586733, 4.560706, 4.551862, 4.558817, 
    4.584635, 4.619225, 4.660789, 4.706684, 4.75217, 4.793106, 4.82573, 
    4.84728, 4.85427, 4.84457, 4.828547, 4.805531, 4.782758, 4.767636, 
    4.765727, 4.779678, 4.809348, 4.852722, 4.90692, 4.968901, 5.035783, 
    5.104878, 5.173582, 5.2392, 5.2988, 5.349137, 5.386735, 5.408215, 5.410872,
  // height(9,15, 0-49)
    5.205245, 5.233704, 5.251448, 5.256646, 5.248955, 5.229216, 5.198977, 
    5.160035, 5.114126, 5.062756, 5.007135, 4.948183, 4.886503, 4.822322, 
    4.75529, 4.674098, 4.592133, 4.552732, 4.529696, 4.523179, 4.532108, 
    4.559325, 4.595654, 4.639558, 4.689092, 4.739789, 4.787691, 4.828758, 
    4.859601, 4.875039, 4.871017, 4.856003, 4.828897, 4.797172, 4.769747, 
    4.754407, 4.755836, 4.775146, 4.810735, 4.859603, 4.918382, 4.983872, 
    5.053164, 5.123552, 5.192328, 5.2566, 5.31316, 5.358506, 5.389058, 5.40165,
  // height(9,16, 0-49)
    5.205641, 5.232349, 5.248367, 5.25215, 5.243571, 5.223566, 5.193663, 
    5.155571, 5.1109, 5.061044, 5.007129, 4.950017, 4.890282, 4.828084, 
    4.762897, 4.667199, 4.558082, 4.524595, 4.505179, 4.500589, 4.510473, 
    4.537367, 4.573853, 4.618652, 4.670533, 4.725457, 4.779788, 4.82938, 
    4.870381, 4.896234, 4.90115, 4.890569, 4.862889, 4.82492, 4.786451, 
    4.75743, 4.745025, 4.7522, 4.7782, 4.820086, 4.874176, 4.936878, 
    5.004986, 5.075613, 5.145999, 5.21328, 5.274343, 5.325768, 5.363969, 
    5.385563,
  // height(9,17, 0-49)
    5.206429, 5.23244, 5.24809, 5.25195, 5.243927, 5.22491, 5.196322, 
    5.159752, 5.116711, 5.068528, 5.016322, 4.960996, 4.903182, 4.84309, 
    4.780164, 4.665139, 4.525096, 4.499957, 4.484663, 4.481379, 4.491128, 
    4.516054, 4.551351, 4.595904, 4.649085, 4.707342, 4.767391, 4.825082, 
    4.876275, 4.913509, 4.929801, 4.926649, 4.902213, 4.861757, 4.814963, 
    4.77341, 4.746902, 4.740796, 4.755741, 4.789182, 4.837222, 4.895868, 
    4.96155, 5.03114, 5.101774, 5.170614, 5.234653, 5.290627, 5.335063, 
    5.36453,
  // height(9,18, 0-49)
    5.208497, 5.234978, 5.251599, 5.256881, 5.250602, 5.233477, 5.206757, 
    5.171896, 5.13033, 5.083377, 5.032204, 4.977786, 4.920807, 4.861402, 
    4.798707, 4.662005, 4.489505, 4.475817, 4.465091, 4.462282, 4.47091, 
    4.492671, 4.525987, 4.569733, 4.623669, 4.684685, 4.74978, 4.814837, 
    4.875535, 4.924022, 4.952873, 4.959058, 4.941103, 4.902152, 4.850769, 
    4.799243, 4.759669, 4.740109, 4.743153, 4.767068, 4.80796, 4.861491, 
    4.9237, 4.991181, 5.060933, 5.130117, 5.195842, 5.255026, 5.304377, 
    5.340523,
  // height(9,19, 0-49)
    5.212205, 5.240322, 5.25919, 5.267125, 5.263608, 5.249043, 5.224416, 
    5.191014, 5.150217, 5.103388, 5.051769, 4.996344, 4.937584, 4.874966, 
    4.806328, 4.651233, 4.447761, 4.448816, 4.443101, 4.439723, 4.446472, 
    4.464695, 4.496089, 4.539269, 4.594101, 4.657805, 4.727543, 4.799196, 
    4.868299, 4.927033, 4.968306, 4.984324, 4.974784, 4.940611, 4.888542, 
    4.830527, 4.780185, 4.748146, 4.739299, 4.753189, 4.786242, 4.833904, 
    4.891861, 4.956418, 5.024415, 5.092998, 5.159379, 5.220663, 5.273758, 
    5.315415,
  // height(9,20, 0-49)
    5.212728, 5.239095, 5.257136, 5.265122, 5.262591, 5.250175, 5.229265, 
    5.201706, 5.169541, 5.134852, 5.099675, 5.065902, 5.035129, 5.008301, 
    4.984965, 0, 4.281867, 4.296238, 4.319592, 4.349007, 4.384036, 4.42006, 
    4.463272, 4.513869, 4.573604, 4.641306, 4.715052, 4.791258, 4.865699, 
    4.931174, 4.981727, 5.005177, 5.003088, 4.974547, 4.924257, 4.862964, 
    4.804741, 4.762134, 4.742292, 4.746347, 4.771365, 4.812787, 4.866036, 
    4.927151, 4.99281, 5.06013, 5.12641, 5.188928, 5.244792, 5.290888,
  // height(9,21, 0-49)
    5.21802, 5.246518, 5.267158, 5.277958, 5.278198, 5.26831, 5.249588, 
    5.223853, 5.193182, 5.159711, 5.125531, 5.092601, 5.062645, 5.036921, 
    5.015751, 0, 4.280171, 4.286097, 4.301404, 4.32449, 4.355588, 4.38597, 
    4.42638, 4.475754, 4.535542, 4.604822, 4.681754, 4.762756, 4.84341, 
    4.91684, 4.978211, 5.011083, 5.019394, 5.000573, 4.957034, 4.897546, 
    4.835649, 4.785192, 4.75563, 4.750137, 4.766894, 4.801638, 4.849658, 
    4.906757, 4.969437, 5.034751, 5.100053, 5.162745, 5.22009, 5.269087,
  // height(9,22, 0-49)
    5.22302, 5.253256, 5.275841, 5.288589, 5.290601, 5.282212, 5.264708, 
    5.239964, 5.210128, 5.177406, 5.143931, 5.111705, 5.082527, 5.057864, 
    5.038573, 0, 4.278119, 4.278525, 4.288034, 4.306596, 4.335303, 4.361061, 
    4.399333, 4.447818, 4.507654, 4.578084, 4.657235, 4.741405, 4.825919, 
    4.904216, 4.972783, 5.011243, 5.026633, 5.015471, 4.978484, 4.922526, 
    4.859972, 4.804983, 4.768548, 4.755605, 4.765541, 4.794574, 4.838022, 
    4.891535, 4.95148, 5.014856, 5.079045, 5.141546, 5.199745, 5.250741,
  // height(9,23, 0-49)
    5.226744, 5.258028, 5.281734, 5.295559, 5.298512, 5.290893, 5.27401, 
    5.249787, 5.220436, 5.188205, 5.155255, 5.1236, 5.095076, 5.07127, 
    5.053352, 0, 4.279414, 4.276551, 4.281965, 4.297147, 4.32407, 4.345681, 
    4.381749, 4.428933, 4.488155, 4.558842, 4.639098, 4.725091, 4.811872, 
    4.893102, 4.966422, 5.00808, 5.028121, 5.022609, 4.991148, 4.939076, 
    4.877542, 4.820482, 4.779746, 4.76159, 4.766459, 4.791107, 4.830965, 
    4.881619, 4.93934, 5.001071, 5.064211, 5.126318, 5.184858, 5.237008,
  // height(9,24, 0-49)
    5.228496, 5.259939, 5.283836, 5.297881, 5.301076, 5.293717, 5.277114, 
    5.253204, 5.224204, 5.192366, 5.159845, 5.128648, 5.100616, 5.077384, 
    5.060251, 0, 4.283651, 4.279233, 4.282315, 4.295458, 4.321284, 4.339952, 
    4.374256, 4.42016, 4.47849, 4.548845, 4.629343, 4.716074, 4.803885, 
    4.886553, 4.962506, 5.005624, 5.028133, 5.025902, 4.997901, 4.948527, 
    4.888073, 4.830173, 4.787071, 4.765799, 4.767502, 4.789327, 4.826833, 
    4.875592, 4.931826, 4.992456, 5.054884, 5.116711, 5.175456, 5.228333,
  // height(9,25, 0-49)
    5.22796, 5.258594, 5.281716, 5.295139, 5.297939, 5.290426, 5.27388, 
    5.250185, 5.221498, 5.190021, 5.157872, 5.127028, 5.099308, 5.07633, 
    5.059365, 0, 4.289196, 4.284725, 4.287505, 4.300285, 4.325872, 4.343461, 
    4.376945, 4.422066, 4.479642, 4.549365, 4.629392, 4.715792, 4.803343, 
    4.885863, 4.962089, 5.004999, 5.027723, 5.026116, 4.998996, 4.950472, 
    4.89053, 4.832613, 4.789001, 4.766916, 4.767715, 4.788686, 4.825451, 
    4.87359, 4.929327, 4.989579, 5.051758, 5.113479, 5.17228, 5.22539,
  // height(9,26, 0-49)
    5.225247, 5.254143, 5.275551, 5.287515, 5.289261, 5.281141, 5.26438, 
    5.240758, 5.21231, 5.18114, 5.149289, 5.11869, 5.091106, 5.068068, 
    5.050664, 0, 4.295433, 4.292458, 4.29705, 4.311205, 4.33739, 4.355901, 
    4.389616, 4.434559, 4.491645, 4.560555, 4.639478, 4.724538, 4.810594, 
    4.891437, 4.965577, 5.006762, 5.027511, 5.023829, 4.99484, 4.945057, 
    4.88476, 4.827417, 4.78503, 4.764428, 4.766649, 4.788824, 4.826549, 
    4.875436, 4.931742, 4.99241, 5.054859, 5.116698, 5.175449, 5.22833,
  // height(9,27, 0-49)
    5.220861, 5.247246, 5.266091, 5.275759, 5.275703, 5.266364, 5.248924, 
    5.225036, 5.196589, 5.16555, 5.133861, 5.103376, 5.075775, 5.052415, 
    5.034029, 0, 4.302463, 4.302832, 4.311277, 4.328385, 4.355904, 4.377017, 
    4.411754, 4.456905, 4.513578, 4.58136, 4.658477, 4.741166, 4.824496, 
    4.902151, 4.97192, 5.009845, 5.026492, 5.018219, 4.984942, 4.932204, 
    4.871093, 4.815196, 4.775881, 4.759018, 4.764867, 4.790172, 4.830435, 
    4.881328, 4.939181, 5.000987, 5.064165, 5.126294, 5.184847, 5.237001,
  // height(9,28, 0-49)
    5.215629, 5.238973, 5.254549, 5.261092, 5.258357, 5.246945, 5.228058, 
    5.203263, 5.174317, 5.143045, 5.111273, 5.080747, 5.053013, 5.029168, 
    5.009374, 0, 4.311146, 4.317119, 4.331298, 4.35264, 4.382026, 4.406691, 
    4.442622, 4.4878, 4.543655, 4.609676, 4.684156, 4.763472, 4.842965, 
    4.916097, 4.979532, 5.0127, 5.023324, 5.008373, 4.969041, 4.912435, 
    4.850762, 4.797608, 4.763256, 4.75213, 4.763408, 4.793327, 4.837316, 
    4.891145, 4.951268, 5.014741, 5.078983, 5.141513, 5.199726, 5.250731,
  // height(9,29, 0-49)
    5.210575, 5.230656, 5.242446, 5.245065, 5.238635, 5.224026, 5.202578, 
    5.175876, 5.145615, 5.11352, 5.081297, 5.050559, 5.022669, 4.99836, 
    4.977002, 0, 4.32097, 4.335202, 4.357126, 4.384002, 4.415863, 4.444396, 
    4.481161, 4.525657, 4.579839, 4.643129, 4.713893, 4.78861, 4.862862, 
    4.929764, 4.984661, 5.011045, 5.013606, 4.990396, 4.944409, 4.88464, 
    4.824273, 4.776336, 4.749413, 4.746114, 4.764445, 4.80021, 4.84885, 
    4.906308, 4.96919, 5.034617, 5.099981, 5.162707, 5.22007, 5.269075,
  // height(9,30, 0-49)
    5.211185, 5.232265, 5.243868, 5.245254, 5.236584, 5.218601, 5.192334, 
    5.158899, 5.119413, 5.074954, 5.0265, 4.974833, 4.92029, 4.862335, 
    4.799018, 4.650102, 4.46623, 4.474145, 4.474097, 4.474111, 4.482029, 
    4.496277, 4.523712, 4.562758, 4.613616, 4.67399, 4.741224, 4.811243, 
    4.879523, 4.938704, 4.982891, 5.000132, 4.992626, 4.960247, 4.908324, 
    4.847715, 4.791922, 4.752495, 4.735684, 4.742134, 4.768816, 4.811302, 
    4.865192, 4.926679, 4.992549, 5.059987, 5.126332, 5.188886, 5.244769, 
    5.290876,
  // height(9,31, 0-49)
    5.20908, 5.227884, 5.236427, 5.234247, 5.221874, 5.200438, 5.171289, 
    5.135762, 5.095062, 5.050255, 5.002267, 4.951888, 4.899677, 4.845722, 
    4.789222, 4.658228, 4.501397, 4.496706, 4.493328, 4.495354, 4.506206, 
    4.525119, 4.554814, 4.594297, 4.643971, 4.701432, 4.764091, 4.828028, 
    4.888942, 4.939219, 4.972041, 4.980291, 4.964257, 4.925714, 4.87197, 
    4.814879, 4.767239, 4.738547, 4.732779, 4.749048, 4.783735, 4.832435, 
    4.89102, 4.955945, 5.024151, 5.092851, 5.159298, 5.220619, 5.273735, 
    5.315403,
  // height(9,32, 0-49)
    5.209422, 5.227388, 5.234317, 5.229859, 5.214752, 5.190379, 5.15834, 
    5.120173, 5.077215, 5.030576, 4.981167, 4.929723, 4.876769, 4.822464, 
    4.766259, 4.657221, 4.530038, 4.515179, 4.508562, 4.511379, 4.524328, 
    4.547682, 4.579953, 4.620469, 4.669526, 4.724418, 4.782448, 4.839732, 
    4.892161, 4.932154, 4.95264, 4.951416, 4.927637, 4.885253, 4.833202, 
    4.783412, 4.747004, 4.730926, 4.736993, 4.76317, 4.805598, 4.860101, 
    4.922898, 4.990724, 5.060675, 5.129973, 5.195764, 5.254982, 5.304353, 
    5.340511,
  // height(9,33, 0-49)
    5.211784, 5.230331, 5.23714, 5.231805, 5.215128, 5.188638, 5.154125, 
    5.113319, 5.067709, 5.018507, 4.966658, 4.912882, 4.857656, 4.801088, 
    4.742635, 4.653386, 4.555256, 4.532505, 4.522496, 4.524918, 4.538918, 
    4.565711, 4.600144, 4.641606, 4.68998, 4.742125, 4.795075, 4.84495, 
    4.887879, 4.916761, 4.925084, 4.915268, 4.8861, 4.843475, 4.797151, 
    4.758084, 4.735029, 4.73236, 4.75014, 4.785647, 4.835072, 4.894595, 
    4.960809, 5.030715, 5.101532, 5.170478, 5.234578, 5.290584, 5.33504, 
    5.364517,
  // height(9,34, 0-49)
    5.215219, 5.235668, 5.243885, 5.23924, 5.222435, 5.195026, 5.158927, 
    5.11603, 5.067999, 5.016191, 4.961662, 4.905194, 4.847309, 4.788183, 
    4.727444, 4.6529, 4.580625, 4.55162, 4.538008, 4.538926, 4.552721, 
    4.581357, 4.616908, 4.658594, 4.70565, 4.754443, 4.80167, 4.843497, 
    4.87642, 4.894343, 4.89206, 4.875939, 4.844918, 4.806159, 4.769204, 
    4.743195, 4.734305, 4.744707, 4.773262, 4.816971, 4.872271, 4.935742, 
    5.004318, 5.075227, 5.145776, 5.213154, 5.274272, 5.325727, 5.363947, 
    5.38555,
  // height(9,35, 0-49)
    5.218414, 5.241881, 5.252987, 5.250708, 5.235466, 5.208694, 5.172336, 
    5.12841, 5.078754, 5.02491, 4.968103, 4.90927, 4.849085, 4.787934, 
    4.725807, 4.660797, 4.609091, 4.575197, 4.557967, 4.556472, 4.56875, 
    4.597325, 4.632507, 4.673204, 4.717884, 4.762468, 4.803359, 4.83689, 
    4.860095, 4.868361, 4.85827, 4.839107, 4.810142, 4.778883, 4.753745, 
    4.741656, 4.746446, 4.768659, 4.806472, 4.856906, 4.916722, 4.98287, 
    5.052571, 5.123204, 5.192127, 5.256485, 5.313095, 5.358469, 5.389037, 
    5.401639,
  // height(9,36, 0-49)
    5.219895, 5.247176, 5.262488, 5.264244, 5.252396, 5.228087, 5.193159, 
    5.149686, 5.099665, 5.044836, 4.98664, 4.926233, 4.864524, 4.80219, 
    4.739642, 4.680242, 4.642906, 4.605454, 4.584847, 4.580313, 4.589905, 
    4.616549, 4.649711, 4.687962, 4.729007, 4.768494, 4.802673, 4.828212, 
    4.842849, 4.843726, 4.829322, 4.810611, 4.787079, 4.765726, 4.753314, 
    4.754615, 4.771617, 4.803811, 4.849074, 4.904593, 4.967452, 5.034897, 
    5.104344, 5.173264, 5.239013, 5.29869, 5.349073, 5.3867, 5.408195, 
    5.410862,
  // height(9,37, 0-49)
    5.218255, 5.249717, 5.27024, 5.277552, 5.270936, 5.25105, 5.219474, 
    5.178236, 5.129437, 5.075015, 5.016646, 4.955743, 4.893483, 4.830852, 
    4.76865, 4.712382, 4.683611, 4.643882, 4.620321, 4.612436, 4.618487, 
    4.641649, 4.671282, 4.705679, 4.741915, 4.775605, 4.803057, 4.82145, 
    4.829312, 4.825551, 4.810279, 4.794975, 4.779095, 4.768571, 4.768416, 
    4.7816, 4.808813, 4.848932, 4.899767, 4.958707, 5.023099, 5.090394, 
    5.158112, 5.223743, 5.284613, 5.33779, 5.380095, 5.408271, 5.419396, 
    5.411546,
  // height(9,38, 0-49)
    5.212383, 5.247881, 5.274166, 5.288225, 5.288517, 5.274992, 5.248788, 
    5.21174, 5.165967, 5.113562, 5.056436, 4.996264, 4.934503, 4.87243, 
    4.811168, 4.756728, 4.73197, 4.691082, 4.665075, 4.653807, 4.65584, 
    4.674464, 4.699435, 4.72888, 4.759443, 4.786973, 4.808064, 4.820529, 
    4.823663, 4.81791, 4.804527, 4.794577, 4.787253, 4.787226, 4.797941, 
    4.821002, 4.856258, 4.902263, 4.956853, 5.017594, 5.082009, 5.147655, 
    5.212077, 5.272727, 5.326886, 5.371646, 5.404006, 5.421148, 5.420925, 
    5.402503,
  // height(9,39, 0-49)
    5.20167, 5.240501, 5.272511, 5.294001, 5.302503, 5.297089, 5.278226, 
    5.247378, 5.20655, 5.157911, 5.103568, 5.045445, 4.985273, 4.924599, 
    4.864816, 4.811718, 4.787943, 4.746778, 4.718848, 4.70439, 4.702281, 
    4.715828, 4.73548, 4.759322, 4.783782, 4.805178, 4.82057, 4.828451, 
    4.828772, 4.823126, 4.813404, 4.809672, 4.810735, 4.820044, 4.839785, 
    4.870599, 4.911798, 4.96177, 5.018401, 5.079369, 5.142285, 5.204723, 
    5.264188, 5.318067, 5.363621, 5.398062, 5.418763, 5.423631, 5.411623, 
    5.383276,
  // height(9,40, 0-49)
    5.186132, 5.22708, 5.264103, 5.293013, 5.310456, 5.314495, 5.304725, 
    5.282016, 5.248078, 5.205032, 5.155106, 5.100437, 5.043005, 4.984615, 
    4.926899, 4.87519, 4.850765, 4.809989, 4.780656, 4.763356, 4.757268, 
    4.765635, 4.779768, 4.797813, 4.816178, 4.8318, 4.84232, 4.846885, 
    4.845916, 4.841768, 4.836526, 4.838995, 4.847562, 4.864634, 4.891436, 
    4.927948, 4.973135, 5.025293, 5.082327, 5.141959, 5.201804, 5.259393, 
    5.312152, 5.357416, 5.392503, 5.414909, 5.422629, 5.414599, 5.391162, 
    5.354355,
  // height(9,41, 0-49)
    5.166451, 5.207902, 5.248558, 5.28407, 5.310394, 5.324593, 5.325236, 
    5.312375, 5.287194, 5.251593, 5.207793, 5.158082, 5.10465, 5.049539, 
    4.994611, 4.944724, 4.91911, 4.879265, 4.849064, 4.829385, 4.819679, 
    4.823095, 4.831874, 4.844314, 4.856938, 4.867391, 4.873917, 4.876226, 
    4.875024, 4.873092, 4.872416, 4.880478, 4.895287, 4.918398, 4.950332, 
    4.990605, 5.037953, 5.090587, 5.146398, 5.203084, 5.258206, 5.309211, 
    5.353455, 5.388292, 5.41125, 5.42033, 5.414435, 5.393792, 5.360259, 
    5.317256,
  // height(9,42, 0-49)
    5.143857, 5.184021, 5.226386, 5.266863, 5.301079, 5.325276, 5.336976, 
    5.335222, 5.320437, 5.294066, 5.258155, 5.215016, 5.166993, 5.116336, 
    5.06512, 5.017797, 4.99126, 4.952888, 4.922406, 4.90091, 4.888094, 
    4.887012, 4.890862, 4.898168, 4.905657, 4.911681, 4.915056, 4.915931, 
    4.915131, 4.915613, 4.919096, 4.931798, 4.951411, 4.978819, 5.014019, 
    5.056201, 5.103926, 5.155319, 5.208214, 5.260242, 5.308877, 5.35149, 
    5.38544, 5.408236, 5.417833, 5.413025, 5.393868, 5.362019, 5.320735, 
    5.274421,
  // height(9,43, 0-49)
    5.119925, 5.157089, 5.198948, 5.24208, 5.282256, 5.315266, 5.337736, 
    5.347641, 5.344442, 5.32887, 5.302574, 5.267717, 5.226689, 5.18188, 
    5.135561, 5.09184, 5.065246, 5.028996, 4.998917, 4.976262, 4.960958, 
    4.95599, 4.955519, 4.958347, 4.961455, 4.963848, 4.964833, 4.96487, 
    4.964771, 4.967505, 4.974444, 4.990649, 5.013561, 5.043531, 5.080167, 
    5.122412, 5.168684, 5.217022, 5.265179, 5.3107, 5.350989, 5.383418, 
    5.405475, 5.415052, 5.410805, 5.392574, 5.361722, 5.321233, 5.275365, 
    5.228883,
  // height(9,44, 0-49)
    5.096272, 5.129057, 5.168241, 5.211352, 5.254784, 5.29438, 5.326228, 
    5.34737, 5.35621, 5.352563, 5.337418, 5.312571, 5.280278, 5.24296, 
    5.203005, 5.164229, 5.138921, 5.105624, 5.076772, 5.053725, 5.036647, 
    5.028522, 5.024458, 5.023581, 5.023133, 5.022689, 5.021945, 5.021548, 
    5.022201, 5.026792, 5.036315, 5.054803, 5.079486, 5.110286, 5.146511, 
    5.186906, 5.22978, 5.273088, 5.314514, 5.351556, 5.381634, 5.402251, 
    5.411257, 5.407187, 5.389662, 5.359727, 5.319985, 5.274365, 5.22749, 
    5.183779,
  // height(9,45, 0-49)
    5.074281, 5.101814, 5.136524, 5.17699, 5.220571, 5.263685, 5.302406, 
    5.333194, 5.353523, 5.36219, 5.359307, 5.346044, 5.324288, 5.296298, 
    5.264447, 5.232249, 5.209951, 5.180675, 5.154027, 5.131465, 5.113417, 
    5.102954, 5.096113, 5.092372, 5.089212, 5.08668, 5.084756, 5.084169, 
    5.085434, 5.091334, 5.102482, 5.122004, 5.14693, 5.17682, 5.210737, 
    5.247275, 5.284656, 5.320791, 5.353364, 5.379928, 5.39808, 5.405691, 
    5.401236, 5.384155, 5.355194, 5.316544, 5.271692, 5.224903, 5.180446, 
    5.141823,
  // height(9,46, 0-49)
    5.0549, 5.07686, 5.105901, 5.141548, 5.18226, 5.22542, 5.26764, 5.305339, 
    5.335418, 5.355771, 5.36553, 5.365007, 5.355437, 5.338662, 5.316822, 
    5.293051, 5.275785, 5.251806, 5.228491, 5.207395, 5.189259, 5.177374, 
    5.168643, 5.162926, 5.157879, 5.153938, 5.151259, 5.150574, 5.152169, 
    5.158724, 5.17048, 5.189789, 5.213448, 5.240694, 5.270373, 5.30097, 
    5.330666, 5.357411, 5.379015, 5.393284, 5.398237, 5.392398, 5.375129, 
    5.346938, 5.309633, 5.26622, 5.22047, 5.176284, 5.136996, 5.104896,
  // height(9,47, 0-49)
    5.038558, 5.055104, 5.07795, 5.107332, 5.142719, 5.182619, 5.224613, 
    5.265657, 5.302625, 5.332863, 5.354623, 5.367231, 5.371015, 5.367095, 
    5.3571, 5.343633, 5.333583, 5.316318, 5.297566, 5.279008, 5.261748, 
    5.249465, 5.23981, 5.233042, 5.226902, 5.222136, 5.219, 5.218166, 
    5.219665, 5.226124, 5.237422, 5.255292, 5.276211, 5.299119, 5.322676, 
    5.345291, 5.365184, 5.380476, 5.389296, 5.389965, 5.381234, 5.362558, 
    5.334355, 5.298147, 5.256485, 5.212605, 5.169889, 5.131297, 5.098928, 
    5.073874,
  // height(9,48, 0-49)
    5.025191, 5.036808, 5.053524, 5.076003, 5.104483, 5.138533, 5.17689, 
    5.217495, 5.257764, 5.295023, 5.326963, 5.351994, 5.369394, 5.379289, 
    5.382505, 5.380936, 5.380241, 5.371087, 5.358146, 5.343263, 5.327931, 
    5.316406, 5.306894, 5.300048, 5.293569, 5.288468, 5.285032, 5.28385, 
    5.284679, 5.29018, 5.29989, 5.31511, 5.331882, 5.348882, 5.364614, 
    5.377472, 5.385822, 5.388123, 5.38307, 5.369785, 5.348024, 5.318344, 
    5.282197, 5.241826, 5.199984, 5.1595, 5.122818, 5.091662, 5.06691, 
    5.048687,
  // height(9,49, 0-49)
    5.012385, 5.018913, 5.028864, 5.043107, 5.062448, 5.087427, 5.118075, 
    5.153737, 5.193004, 5.233839, 5.273879, 5.31083, 5.342823, 5.368688, 
    5.388059, 5.402215, 5.418763, 5.421006, 5.415788, 5.405649, 5.392869, 
    5.385442, 5.379874, 5.377387, 5.372908, 5.368307, 5.363704, 5.359727, 
    5.355256, 5.355647, 5.359989, 5.371101, 5.38187, 5.390671, 5.395897, 
    5.396035, 5.389802, 5.3763, 5.355184, 5.326793, 5.292233, 5.253324, 
    5.212403, 5.171985, 5.134371, 5.101318, 5.073847, 5.052252, 5.036246, 
    5.025198,
  // height(10,0, 0-49)
    5.063582, 5.085031, 5.112928, 5.146696, 5.184947, 5.225497, 5.265574, 
    5.302221, 5.332746, 5.355133, 5.368267, 5.371976, 5.366912, 5.354355, 
    5.335983, 5.3139, 5.291661, 5.267425, 5.244224, 5.223267, 5.205225, 
    5.190944, 5.179907, 5.172104, 5.167113, 5.164995, 5.165788, 5.169702, 
    5.176876, 5.187829, 5.202584, 5.221438, 5.243492, 5.268015, 5.293913, 
    5.31977, 5.34392, 5.364543, 5.379786, 5.387915, 5.38752, 5.377726, 
    5.358419, 5.3304, 5.295416, 5.256012, 5.215207, 5.176044, 5.141145, 
    5.112394,
  // height(10,1, 0-49)
    5.079928, 5.105417, 5.137311, 5.174423, 5.214681, 5.255301, 5.293159, 
    5.325284, 5.349298, 5.363727, 5.368092, 5.362825, 5.349079, 5.32849, 
    5.302971, 5.274961, 5.249591, 5.22163, 5.19565, 5.1729, 5.153946, 
    5.139993, 5.129792, 5.123188, 5.119247, 5.117973, 5.119292, 5.123413, 
    5.130458, 5.141384, 5.156361, 5.176321, 5.200119, 5.227235, 5.256737, 
    5.287312, 5.31734, 5.344975, 5.368256, 5.385231, 5.394138, 5.393606, 
    5.382902, 5.362143, 5.332445, 5.295923, 5.255486, 5.214435, 5.175961, 
    5.142664,
  // height(10,2, 0-49)
    5.100276, 5.12977, 5.1649, 5.203756, 5.243615, 5.281312, 5.313743, 
    5.338332, 5.35337, 5.358143, 5.352868, 5.338513, 5.316582, 5.288897, 
    5.257421, 5.224789, 5.197577, 5.167107, 5.139554, 5.116156, 5.097363, 
    5.084681, 5.076171, 5.071518, 5.069331, 5.069472, 5.071693, 5.076145, 
    5.082903, 5.093283, 5.107612, 5.127469, 5.151559, 5.179631, 5.210985, 
    5.244498, 5.27869, 5.311812, 5.34193, 5.367047, 5.385226, 5.394764, 
    5.394402, 5.383549, 5.362504, 5.332596, 5.296147, 5.256245, 5.216292, 
    5.179459,
  // height(10,3, 0-49)
    5.123564, 5.156494, 5.193518, 5.232036, 5.268888, 5.30088, 5.325299, 
    5.340286, 5.344973, 5.33944, 5.324524, 5.3016, 5.27236, 5.238668, 
    5.202416, 5.166353, 5.138496, 5.1065, 5.078358, 5.055256, 5.03751, 
    5.026891, 5.020802, 5.018765, 5.018983, 5.021102, 5.024645, 5.029631, 
    5.036055, 5.045497, 5.058444, 5.077137, 5.100204, 5.127726, 5.159303, 
    5.194069, 5.230758, 5.267785, 5.303344, 5.335496, 5.362273, 5.381793, 
    5.39242, 5.392964, 5.382909, 5.362636, 5.33356, 5.298093, 5.259374, 
    5.220767,
  // height(10,4, 0-49)
    5.148277, 5.183551, 5.220681, 5.256588, 5.288019, 5.312116, 5.326862, 
    5.331258, 5.325281, 5.309696, 5.285806, 5.25523, 5.219736, 5.181118, 
    5.141133, 5.102629, 5.075132, 5.042326, 5.01433, 4.99224, 4.976225, 
    4.968293, 4.965206, 4.966337, 4.969534, 4.974173, 4.979482, 4.985287, 
    4.991461, 4.999736, 5.010735, 5.027388, 5.048301, 5.073945, 5.104287, 
    5.138782, 5.176426, 5.215847, 5.255407, 5.293285, 5.327562, 5.356293, 
    5.377622, 5.389924, 5.392003, 5.383332, 5.364291, 5.336296, 5.301751, 
    5.263733,
  // height(10,5, 0-49)
    5.17261, 5.208737, 5.244016, 5.275208, 5.299335, 5.314187, 5.318586, 
    5.31239, 5.29629, 5.271561, 5.239791, 5.202709, 5.162052, 5.119503, 
    5.076645, 5.036462, 5.010109, 4.97695, 4.949606, 4.929027, 4.91522, 
    4.910427, 4.91076, 4.915475, 4.92213, 4.929779, 4.937321, 4.944317, 
    4.950469, 4.957533, 4.96622, 4.980175, 4.998003, 5.020619, 5.048433, 
    5.081285, 5.118479, 5.158883, 5.201038, 5.243255, 5.283694, 5.320426, 
    5.351492, 5.375001, 5.389269, 5.393025, 5.385661, 5.367476, 5.339813, 
    5.305001,
  // height(10,6, 0-49)
    5.194726, 5.230039, 5.261647, 5.286497, 5.302191, 5.307335, 5.301603, 
    5.285583, 5.260492, 5.227921, 5.189589, 5.147222, 5.102467, 5.056863, 
    5.011828, 4.97053, 4.945855, 4.912601, 4.886216, 4.867458, 4.85615, 
    4.854763, 4.858765, 4.867326, 4.877797, 4.888885, 4.899129, 4.907778, 
    4.914294, 4.920318, 4.926564, 4.9374, 4.951415, 4.97002, 4.994144, 
    5.024087, 5.059518, 5.099563, 5.142944, 5.188095, 5.233257, 5.276544, 
    5.315973, 5.349518, 5.375189, 5.391176, 5.396054, 5.389062, 5.370367, 
    5.341236,
  // height(10,7, 0-49)
    5.213053, 5.245964, 5.27248, 5.290026, 5.296961, 5.292734, 5.27777, 
    5.253204, 5.220595, 5.181672, 5.138168, 5.091727, 5.04387, 4.995987, 
    4.949328, 4.907313, 4.88458, 4.851351, 4.826089, 4.809305, 4.800615, 
    4.802724, 4.810457, 4.822952, 4.837451, 4.852314, 4.865723, 4.876563, 
    4.88401, 4.889411, 4.893355, 4.900923, 4.910622, 4.924387, 4.94375, 
    4.969565, 5.001939, 5.040301, 5.083554, 5.130239, 5.178657, 5.226962, 
    5.27318, 5.315236, 5.350972, 5.378225, 5.394969, 5.399563, 5.391072, 
    5.369621,
  // height(10,8, 0-49)
    5.226548, 5.255755, 5.276319, 5.286304, 5.284873, 5.272231, 5.249386, 
    5.217844, 5.179329, 5.135591, 5.088283, 5.038926, 4.98889, 4.939411, 
    4.891582, 4.849094, 4.828224, 4.795094, 4.771032, 4.756248, 4.750131, 
    4.755633, 4.766952, 4.783258, 4.801815, 4.820665, 4.837659, 4.851306, 
    4.860435, 4.865911, 4.868018, 4.872491, 4.877636, 4.885912, 4.899523, 
    4.919997, 4.947987, 4.983297, 5.02504, 5.071846, 5.122056, 5.173835, 
    5.225216, 5.274106, 5.318265, 5.355324, 5.38286, 5.39859, 5.40069, 
    5.388237,
  // height(10,9, 0-49)
    5.234836, 5.259479, 5.273821, 5.276622, 5.26777, 5.248077, 5.218955, 
    5.182111, 5.139313, 5.09224, 5.042422, 4.991228, 4.93987, 4.889423, 
    4.840813, 4.797938, 4.778379, 4.745469, 4.722646, 4.709779, 4.706027, 
    4.714598, 4.729111, 4.748862, 4.77128, 4.794157, 4.815078, 4.832183, 
    4.843925, 4.850475, 4.851599, 4.853556, 4.854271, 4.856665, 4.863659, 
    4.877585, 4.899804, 4.930608, 4.969382, 5.014863, 5.0654, 5.119133, 
    5.17407, 5.228092, 5.27892, 5.324071, 5.360898, 5.386709, 5.399065, 
    5.396215,
  // height(10,10, 0-49)
    5.238247, 5.257951, 5.266341, 5.262815, 5.247848, 5.222678, 5.188955, 
    5.148462, 5.102916, 5.053882, 5.002743, 4.950707, 4.898828, 4.848012, 
    4.798991, 4.755602, 4.736162, 4.703743, 4.682203, 4.671069, 4.66929, 
    4.68035, 4.697388, 4.71993, 4.745744, 4.772466, 4.797513, 4.818703, 
    4.834116, 4.843032, 4.844454, 4.844961, 4.841871, 4.838394, 4.838163, 
    4.844429, 4.859446, 4.88419, 4.918439, 4.961081, 5.01046, 5.064648, 
    5.121579, 5.17908, 5.234825, 5.286284, 5.330706, 5.365195, 5.38696, 
    5.393692,
  // height(10,11, 0-49)
    5.237722, 5.252574, 5.255694, 5.247005, 5.227397, 5.198365, 5.161659, 
    5.119038, 5.072123, 5.022343, 4.970935, 4.918961, 4.86732, 4.81674, 
    4.767717, 4.723385, 4.702055, 4.670654, 4.650481, 4.64079, 4.640394, 
    4.653071, 4.671667, 4.696053, 4.724506, 4.754633, 4.783804, 4.809594, 
    4.829752, 4.842523, 4.845928, 4.846569, 4.840914, 4.832191, 4.824595, 
    4.822354, 4.828823, 4.845907, 4.873978, 4.912177, 4.958867, 5.012014, 
    5.069425, 5.128822, 5.187816, 5.243847, 5.294146, 5.335773, 5.365799, 
    5.381611,
  // height(10,12, 0-49)
    5.234626, 5.245103, 5.243909, 5.231354, 5.20858, 5.177192, 5.138937, 
    5.095491, 5.048359, 4.998839, 4.948044, 4.896914, 4.84622, 4.796515, 
    4.748018, 4.701878, 4.675796, 4.646248, 4.627597, 4.618956, 4.619151, 
    4.632289, 4.651206, 4.676237, 4.706321, 4.739155, 4.772195, 4.802876, 
    4.828703, 4.846828, 4.854155, 4.856939, 4.85062, 4.838054, 4.82369, 
    4.812641, 4.809513, 4.817426, 4.837632, 4.869717, 4.912129, 4.962729, 
    5.019142, 5.078934, 5.139617, 5.198605, 5.253157, 5.300396, 5.33741, 
    5.361478,
  // height(10,13, 0-49)
    5.230535, 5.237388, 5.232965, 5.21782, 5.193212, 5.160748, 5.122097, 
    5.078829, 5.032333, 4.983805, 4.934273, 4.884608, 4.835494, 4.787343, 
    4.740097, 4.690714, 4.656355, 4.629813, 4.612917, 4.604844, 4.60468, 
    4.616896, 4.634736, 4.65907, 4.689609, 4.724247, 4.760649, 4.796208, 
    4.828288, 4.853024, 4.866192, 4.873289, 4.868722, 4.854521, 4.834921, 
    4.81561, 4.802438, 4.8, 4.810771, 4.835072, 4.871596, 4.918133, 4.972108, 
    5.030878, 5.091822, 5.152305, 5.209641, 5.261067, 5.303789, 5.335109,
  // height(10,14, 0-49)
    5.22699, 5.231134, 5.224566, 5.207964, 5.182598, 5.150006, 5.111754, 
    5.069297, 5.023933, 4.976803, 4.928903, 4.881094, 4.834053, 4.788131, 
    4.743088, 4.688396, 4.642111, 4.619964, 4.605116, 4.597078, 4.595531, 
    4.605345, 4.620689, 4.643006, 4.672795, 4.708239, 4.747289, 4.787376, 
    4.82584, 4.857959, 4.878545, 4.891905, 4.89165, 4.878604, 4.856218, 
    4.830238, 4.807499, 4.794166, 4.79429, 4.80929, 4.838372, 4.879369, 
    4.929523, 4.985952, 5.04586, 5.106551, 5.16538, 5.219721, 5.266939, 
    5.304432,
  // height(10,15, 0-49)
    5.225293, 5.227697, 5.219958, 5.202792, 5.177416, 5.145269, 5.107808, 
    5.066401, 5.02229, 4.976607, 4.930377, 4.88452, 4.839792, 4.79663, 
    4.75483, 4.69235, 4.631154, 4.614925, 4.602443, 4.593904, 4.58998, 
    4.595966, 4.607544, 4.62669, 4.65465, 4.689934, 4.730808, 4.7748, 
    4.819294, 4.85896, 4.887938, 4.908922, 4.915213, 4.906217, 4.884106, 
    4.854033, 4.823288, 4.799448, 4.788349, 4.792909, 4.813193, 4.847295, 
    4.892347, 4.94524, 5.002972, 5.062758, 5.12198, 5.17813, 5.228736, 
    5.271329,
  // height(10,16, 0-49)
    5.226336, 5.227925, 5.219817, 5.202703, 5.177724, 5.146221, 5.109568, 
    5.06908, 5.025991, 4.981462, 4.936589, 4.892404, 4.84983, 4.809532, 
    4.771629, 4.699264, 4.621652, 4.61295, 4.603134, 4.593575, 4.586397, 
    4.587306, 4.594104, 4.609207, 4.634496, 4.668808, 4.710706, 4.757823, 
    4.807619, 4.854417, 4.892068, 4.921228, 4.935552, 4.933044, 4.914313, 
    4.883314, 4.847099, 4.81419, 4.792173, 4.785765, 4.796284, 4.822381, 
    4.861237, 4.909564, 4.964163, 5.022121, 5.08082, 5.137845, 5.190862, 
    5.237532,
  // height(10,17, 0-49)
    5.230514, 5.23212, 5.224253, 5.207549, 5.183083, 5.152126, 5.116007, 
    5.076031, 5.033445, 4.989463, 4.945265, 4.902009, 4.860803, 4.822589, 
    4.787977, 4.705591, 4.612271, 4.612747, 4.605839, 4.594719, 4.583512, 
    4.578328, 4.579618, 4.590136, 4.612224, 4.645008, 4.687278, 4.736743, 
    4.790919, 4.844021, 4.890014, 4.927098, 4.949994, 4.955523, 4.94271, 
    4.913936, 4.875333, 4.835699, 4.804019, 4.7869, 4.787251, 4.804621, 
    4.836472, 4.879438, 4.930146, 4.985555, 5.04301, 5.100143, 5.154733, 
    5.204546,
  // height(10,18, 0-49)
    5.237718, 5.240082, 5.232924, 5.216834, 5.19283, 5.162156, 5.126127, 
    5.086053, 5.043212, 4.998859, 4.954231, 4.910549, 4.86899, 4.830619, 
    4.796376, 4.707914, 4.602833, 4.613844, 4.60993, 4.59652, 4.580455, 
    4.568354, 4.563672, 4.569397, 4.588124, 4.619167, 4.66143, 4.712628, 
    4.770273, 4.82866, 4.882247, 4.92637, 4.957467, 4.971514, 4.966166, 
    4.942143, 4.904187, 4.860658, 4.821369, 4.794617, 4.785073, 4.793501, 
    4.817908, 4.85501, 4.901318, 4.953671, 5.009349, 5.066003, 5.121474, 
    5.173612,
  // height(10,19, 0-49)
    5.247415, 5.251267, 5.245289, 5.230013, 5.20642, 5.175728, 5.139245, 
    5.098292, 5.054173, 5.008155, 4.961453, 4.915181, 4.870294, 4.827582, 
    4.788054, 4.702839, 4.595904, 4.617163, 4.615731, 4.598713, 4.576507, 
    4.556717, 4.545831, 4.546948, 4.562612, 4.592149, 4.634409, 4.687026, 
    4.747424, 4.810097, 4.870316, 4.920206, 4.958426, 4.980475, 4.982996, 
    4.965231, 4.930353, 4.885727, 4.841322, 4.806689, 4.788195, 4.788025, 
    4.80498, 4.836047, 4.87772, 4.926739, 4.980312, 5.036072, 5.091892, 
    5.14567,
  // height(10,20, 0-49)
    5.253863, 5.255918, 5.248505, 5.232355, 5.208736, 5.179231, 5.145556, 
    5.109469, 5.072702, 5.036943, 5.003791, 4.974656, 4.950539, 4.931577, 
    4.916345, 0, 4.529047, 4.533604, 4.533447, 4.529254, 4.524078, 4.517531, 
    4.516744, 4.524277, 4.543463, 4.574782, 4.617994, 4.671397, 4.732827, 
    4.797443, 4.86176, 4.91475, 4.957507, 4.985386, 4.994432, 4.982762, 
    4.952068, 4.908407, 4.861261, 4.820816, 4.794822, 4.786893, 4.796811, 
    4.82201, 4.859082, 4.904712, 4.956047, 5.010677, 5.066474, 5.121367,
  // height(10,21, 0-49)
    5.263675, 5.267076, 5.260616, 5.245088, 5.221847, 5.192562, 5.159019, 
    5.122997, 5.086214, 5.050299, 5.016766, 4.986938, 4.961788, 4.941614, 
    4.925509, 0, 4.57267, 4.567389, 4.555607, 4.539651, 4.524162, 4.505689, 
    4.496675, 4.498558, 4.514233, 4.543977, 4.587254, 4.642064, 4.705884, 
    4.773979, 4.843802, 4.901035, 4.949372, 4.984136, 5.000959, 4.997036, 
    4.972662, 4.932421, 4.884916, 4.840544, 4.808241, 4.793121, 4.796153, 
    4.815408, 4.847692, 4.889668, 4.938398, 4.991401, 5.046501, 5.101614,
  // height(10,22, 0-49)
    5.271476, 5.27575, 5.269802, 5.254496, 5.231293, 5.201962, 5.168361, 
    5.132299, 5.095483, 5.059496, 5.025783, 4.995612, 4.969961, 4.949296, 
    4.933185, 0, 4.606127, 4.593786, 4.574115, 4.550414, 4.528358, 4.500781, 
    4.48548, 4.482813, 4.495416, 4.523509, 4.566337, 4.621633, 4.686522, 
    4.756358, 4.829571, 4.888551, 4.939791, 4.978797, 5.001094, 5.003343, 
    4.984809, 4.94875, 4.902673, 4.85667, 4.820312, 4.799883, 4.797452, 
    4.8118, 4.840026, 4.878856, 4.925291, 4.976785, 5.031116, 5.086174,
  // height(10,23, 0-49)
    5.276399, 5.281113, 5.275375, 5.260115, 5.236866, 5.207469, 5.173829, 
    5.13778, 5.101011, 5.065071, 5.031356, 5.001098, 4.975291, 4.954518, 
    4.93868, 0, 4.630615, 4.613832, 4.58922, 4.560673, 4.534565, 4.500163, 
    4.480029, 4.473634, 4.483511, 4.509951, 4.552076, 4.607405, 4.672744, 
    4.743471, 4.818842, 4.878325, 4.930957, 4.972464, 4.998406, 5.005173, 
    4.991349, 4.959182, 4.915194, 4.868976, 4.830346, 4.80637, 4.800004, 
    4.810667, 4.83577, 4.87212, 4.916699, 4.966904, 5.020463, 5.075243,
  // height(10,24, 0-49)
    5.277895, 5.282643, 5.276915, 5.261662, 5.238444, 5.20912, 5.175599, 
    5.139707, 5.103124, 5.067368, 5.033813, 5.003671, 4.977938, 4.957258, 
    4.941692, 0, 4.644578, 4.625749, 4.598795, 4.567974, 4.540061, 4.501756, 
    4.478832, 4.470163, 4.478271, 4.503554, 4.545105, 4.600323, 4.665806, 
    4.736924, 4.813501, 4.87292, 4.926011, 4.96866, 4.996484, 5.005741, 
    4.994654, 4.964887, 4.922336, 4.876217, 4.836404, 4.810391, 4.801668, 
    4.810068, 4.83323, 4.868037, 4.911464, 4.96088, 5.013984, 5.068623,
  // height(10,25, 0-49)
    5.275751, 5.280137, 5.274252, 5.259029, 5.235986, 5.20693, 5.173734, 
    5.138188, 5.10195, 5.066529, 5.033287, 5.003433, 4.977952, 4.957484, 
    4.942075, 0, 4.646362, 4.627713, 4.600918, 4.57033, 4.542782, 4.504051, 
    4.480865, 4.47187, 4.479598, 4.504527, 4.545787, 4.600784, 4.666057, 
    4.736995, 4.813643, 4.872583, 4.925354, 4.967914, 4.995914, 5.005612, 
    4.995152, 4.966033, 4.923948, 4.877962, 4.837917, 4.81139, 4.802017, 
    4.809758, 4.832334, 4.866657, 4.909718, 4.958877, 5.011829, 5.066416,
  // height(10,26, 0-49)
    5.270087, 5.273705, 5.267471, 5.252261, 5.229498, 5.200881, 5.168194, 
    5.133167, 5.097431, 5.062489, 5.029718, 5.00033, 4.975293, 4.955161, 
    4.939804, 0, 4.636261, 4.619933, 4.595723, 4.567776, 4.542617, 4.506954, 
    4.486037, 4.478699, 4.487489, 4.512912, 4.554196, 4.60886, 4.67358, 
    4.743774, 4.819333, 4.877504, 4.92928, 4.970582, 4.997083, 5.005145, 
    4.993102, 4.962729, 4.919972, 4.874004, 4.834575, 4.809024, 4.800726, 
    4.809459, 4.832855, 4.867812, 4.911335, 4.960805, 5.013942, 5.0686,
  // height(10,27, 0-49)
    5.261351, 5.26376, 5.256897, 5.241565, 5.219057, 5.190928, 5.158837, 
    5.124437, 5.089321, 5.054998, 5.022872, 4.994169, 4.969829, 4.950259, 
    4.934984, 0, 4.616155, 4.604306, 4.585077, 4.56209, 4.541208, 4.511642, 
    4.495096, 4.490992, 4.501941, 4.528447, 4.569895, 4.624023, 4.687788, 
    4.756649, 4.829976, 4.887001, 4.937045, 4.975907, 4.999275, 5.003732, 
    4.988097, 4.954829, 4.910524, 4.864675, 4.826832, 4.803771, 4.798227, 
    4.809523, 4.835066, 4.871701, 4.916456, 4.966763, 5.020384, 5.0752,
  // height(10,28, 0-49)
    5.250287, 5.251001, 5.243098, 5.227319, 5.204828, 5.177031, 5.145455, 
    5.111665, 5.077218, 5.043633, 5.012346, 4.984618, 4.961354, 4.942771, 
    4.927911, 0, 4.589266, 4.58401, 4.572131, 4.556344, 4.541521, 4.520256, 
    4.509414, 4.509357, 4.5229, 4.55061, 4.592104, 4.645408, 4.707838, 
    4.774844, 4.844988, 4.900376, 4.947849, 4.983022, 5.001625, 5.000618, 
    4.979618, 4.942165, 4.895842, 4.850533, 4.815399, 4.796301, 4.795027, 
    4.81025, 4.839077, 4.87829, 4.924963, 4.976596, 5.031007, 5.086114,
  // height(10,29, 0-49)
    5.237892, 5.236384, 5.226872, 5.210082, 5.187092, 5.159198, 5.127821, 
    5.094449, 5.060609, 5.027836, 4.997607, 4.971239, 4.949625, 4.9328, 
    4.919292, 0, 4.557674, 4.560971, 4.558987, 4.552932, 4.546215, 4.534846, 
    4.530406, 4.534475, 4.550333, 4.578779, 4.61976, 4.671615, 4.73202, 
    4.796323, 4.862085, 4.914719, 4.958258, 4.988181, 5.000409, 4.992544, 
    4.965331, 4.923674, 4.876193, 4.832937, 4.80229, 4.788859, 4.793301, 
    4.813599, 4.846585, 4.889009, 4.938014, 4.991178, 5.046374, 5.101542,
  // height(10,30, 0-49)
    5.229731, 5.229138, 5.220243, 5.203627, 5.180113, 5.150661, 5.116294, 
    5.078084, 5.037141, 4.994608, 4.951617, 4.909244, 4.868432, 4.829989, 
    4.794954, 4.714292, 4.616234, 4.637926, 4.637839, 4.622587, 4.602194, 
    4.580849, 4.568728, 4.568097, 4.581463, 4.608438, 4.648096, 4.698241, 
    4.756376, 4.817419, 4.877771, 4.926244, 4.964109, 4.986963, 4.99125, 
    4.975613, 4.942276, 4.897612, 4.851018, 4.812195, 4.788252, 4.782269, 
    4.793753, 4.820078, 4.857902, 4.904008, 4.955632, 5.010437, 5.066337, 
    5.121289,
  // height(10,31, 0-49)
    5.219232, 5.216277, 5.205369, 5.187213, 5.162733, 5.132943, 5.098883, 
    5.061612, 5.022202, 4.98176, 4.94143, 4.902367, 4.865702, 4.832438, 
    4.803414, 4.719196, 4.623185, 4.63613, 4.634095, 4.622359, 4.607735, 
    4.594142, 4.588014, 4.591664, 4.607731, 4.635858, 4.675278, 4.723969, 
    4.779628, 4.836938, 4.891286, 4.934981, 4.966794, 4.982536, 4.979336, 
    4.957036, 4.91935, 4.873874, 4.830328, 4.797622, 4.781393, 4.783288, 
    4.801867, 4.834084, 4.87652, 4.926019, 4.979887, 5.035825, 5.091748, 
    5.145588,
  // height(10,32, 0-49)
    5.212204, 5.207666, 5.195166, 5.175536, 5.149817, 5.119109, 5.084501, 
    5.047058, 5.007833, 4.967883, 4.928288, 4.890134, 4.854459, 4.822115, 
    4.793561, 4.715725, 4.631017, 4.635134, 4.631091, 4.622012, 4.61214, 
    4.605616, 4.605232, 4.613331, 4.632458, 4.662114, 4.70151, 4.748676, 
    4.801376, 4.854101, 4.901446, 4.939006, 4.963384, 4.970959, 4.959958, 
    4.931739, 4.891537, 4.847791, 4.809901, 4.785426, 4.77831, 4.788849, 
    4.814866, 4.853093, 4.900144, 4.952962, 5.008929, 5.065755, 5.121329, 
    5.173527,
  // height(10,33, 0-49)
    5.20914, 5.203825, 5.190194, 5.169207, 5.142048, 5.109946, 5.074082, 
    5.035568, 4.995455, 4.954757, 4.914469, 4.875549, 4.838848, 4.804925, 
    4.77372, 4.706617, 4.637273, 4.633828, 4.628059, 4.621222, 4.615577, 
    4.615524, 4.620589, 4.633079, 4.655277, 4.686444, 4.725629, 4.770813, 
    4.819751, 4.866857, 4.906264, 4.936515, 4.952563, 4.951732, 4.933675, 
    4.901386, 4.861358, 4.822259, 4.792506, 4.777924, 4.780762, 4.800201, 
    4.83359, 4.877619, 4.929025, 4.984875, 5.042601, 5.0999, 5.154591, 
    5.204463,
  // height(10,34, 0-49)
    5.210141, 5.204962, 5.190825, 5.168797, 5.140215, 5.106468, 5.068875, 
    5.028635, 4.986836, 4.944474, 4.902484, 4.861712, 4.82285, 4.786231, 
    4.751455, 4.695054, 4.642087, 4.632432, 4.625143, 4.620174, 4.618269, 
    4.623944, 4.634017, 4.650625, 4.67562, 4.707963, 4.746448, 4.788954, 
    4.833173, 4.873645, 4.904438, 4.926645, 4.934232, 4.925783, 4.902545, 
    4.868981, 4.83229, 4.800661, 4.780991, 4.77725, 4.790213, 4.818267, 
    4.858552, 4.907861, 4.963102, 5.021472, 5.080428, 5.137609, 5.190722, 
    5.237449,
  // height(10,35, 0-49)
    5.214813, 5.2108, 5.196992, 5.174516, 5.144845, 5.109542, 5.070085, 
    5.0278, 4.983854, 4.939272, 4.894969, 4.851746, 4.810218, 4.770653, 
    4.732632, 4.684653, 4.646751, 4.632051, 4.62333, 4.619743, 4.620919, 
    4.631336, 4.64574, 4.665937, 4.693183, 4.726111, 4.763205, 4.802227, 
    4.84081, 4.873873, 4.895854, 4.909962, 4.909899, 4.895682, 4.870054, 
    4.838493, 4.808202, 4.78625, 4.777755, 4.784982, 4.807583, 4.843489, 
    4.889846, 4.943633, 5.00196, 5.062129, 5.121593, 5.177893, 5.228593, 
    5.271242,
  // height(10,36, 0-49)
    5.222264, 5.220515, 5.208066, 5.186024, 5.155957, 5.119577, 5.078528, 
    5.03429, 4.988141, 4.941181, 4.894366, 4.848512, 4.804265, 4.76197, 
    4.721433, 4.679046, 4.653185, 4.63448, 4.62433, 4.621491, 4.624862, 
    4.638769, 4.656545, 4.67952, 4.708213, 4.740936, 4.775853, 4.810642, 
    4.842913, 4.868268, 4.881892, 4.888682, 4.882713, 4.865387, 4.840581, 
    4.814148, 4.792623, 4.781571, 4.784374, 4.801928, 4.833148, 4.875787, 
    4.927128, 4.984381, 5.044846, 5.105902, 5.164972, 5.219464, 5.266778, 
    5.30433,
  // height(10,37, 0-49)
    5.231169, 5.232775, 5.222847, 5.202373, 5.172933, 5.13634, 5.094387, 
    5.048704, 5.000711, 4.951622, 4.902481, 4.854186, 4.807487, 4.762895, 
    4.720541, 4.681284, 4.663596, 4.641848, 4.63024, 4.627433, 4.631958, 
    4.647927, 4.667863, 4.692542, 4.721674, 4.753293, 4.785275, 4.815282, 
    4.840997, 4.858955, 4.865395, 4.866431, 4.85696, 4.839487, 4.818485, 
    4.799541, 4.78807, 4.788061, 4.801427, 4.82809, 4.86656, 4.914594, 
    4.969669, 5.029223, 5.090712, 5.15157, 5.209159, 5.260755, 5.303586, 
    5.334973,
  // height(10,38, 0-49)
    5.239892, 5.24584, 5.239644, 5.222045, 5.194521, 5.158906, 5.117092, 
    5.070849, 5.021742, 4.971128, 4.920183, 4.869933, 4.821266, 4.774899, 
    4.73128, 4.693408, 4.680095, 4.656179, 4.643091, 4.639637, 4.644267, 
    4.660845, 4.6816, 4.706756, 4.735232, 4.764845, 4.793278, 4.818267, 
    4.837685, 4.849177, 4.850168, 4.847516, 4.837119, 4.822165, 4.80716, 
    4.796963, 4.795705, 4.805967, 4.828554, 4.862772, 4.906951, 4.958941, 
    5.016412, 5.076992, 5.138256, 5.197663, 5.252513, 5.29996, 5.337116, 
    5.361272,
  // height(10,39, 0-49)
    5.246655, 5.257724, 5.256416, 5.243073, 5.218928, 5.18572, 5.145367, 
    5.099737, 5.050538, 4.999286, 4.947315, 4.895807, 4.845814, 4.798248, 
    4.753822, 4.71631, 4.704317, 4.678978, 4.664438, 4.659803, 4.663629, 
    4.679513, 4.699796, 4.724214, 4.750978, 4.777809, 4.802306, 4.822383, 
    4.83622, 4.842612, 4.840141, 4.835948, 4.826879, 4.816355, 4.808491, 
    4.8072, 4.815392, 4.83454, 4.864683, 4.904767, 4.953069, 5.007549, 
    5.066037, 5.126289, 5.185953, 5.242501, 5.293189, 5.335102, 5.365329, 
    5.381271,
  // height(10,40, 0-49)
    5.249744, 5.266394, 5.270947, 5.263197, 5.243958, 5.214726, 5.177338, 
    5.133704, 5.085651, 5.034855, 4.982824, 4.930913, 4.880349, 4.832219, 
    4.787439, 4.749863, 4.737173, 4.711016, 4.69513, 4.68898, 4.691325, 
    4.705497, 4.724216, 4.746839, 4.771021, 4.794501, 4.81493, 4.830498, 
    4.839759, 4.842586, 4.838536, 4.834641, 4.828501, 4.823401, 4.822832, 
    4.829747, 4.846045, 4.872379, 4.908298, 4.952549, 5.003408, 5.058919, 
    5.117007, 5.175501, 5.232083, 5.284229, 5.329195, 5.364105, 5.386174, 
    5.393111,
  // height(10,41, 0-49)
    5.247719, 5.269979, 5.281053, 5.280043, 5.267168, 5.243511, 5.210688, 
    5.170568, 5.125053, 5.075967, 5.024994, 4.973671, 4.923398, 4.875422, 
    4.830817, 4.79321, 4.778804, 4.752316, 4.735268, 4.727466, 4.727908, 
    4.739669, 4.756018, 4.776052, 4.797035, 4.816849, 4.833313, 4.844961, 
    4.85074, 4.851439, 4.847338, 4.845059, 4.842711, 4.843216, 4.849365, 
    4.863264, 4.886032, 4.917758, 4.95768, 5.004436, 5.056305, 5.111372, 
    5.167601, 5.222831, 5.274746, 5.320846, 5.358463, 5.384906, 5.397736, 
    5.395216,
  // height(10,42, 0-49)
    5.239619, 5.267014, 5.284798, 5.291317, 5.286037, 5.269451, 5.242799, 
    5.207787, 5.166325, 5.120343, 5.071693, 5.02209, 4.973096, 4.926105, 
    4.88232, 4.845045, 4.828703, 4.802299, 4.784326, 4.774885, 4.773208, 
    4.78215, 4.795608, 4.812541, 4.829976, 4.846041, 4.858818, 4.867209, 
    4.870528, 4.870278, 4.867199, 4.867313, 4.869003, 4.87472, 4.886584, 
    4.906005, 4.933528, 4.968866, 5.01106, 5.058681, 5.109999, 5.1631, 
    5.215928, 5.266298, 5.311891, 5.350265, 5.378949, 5.395628, 5.398466, 
    5.386536,
  // height(10,43, 0-49)
    5.225125, 5.256631, 5.280723, 5.295022, 5.298166, 5.289894, 5.270908, 
    5.242608, 5.206801, 5.165462, 5.120562, 5.073971, 5.027399, 4.982369, 
    4.940185, 4.903838, 4.885886, 4.85994, 4.841307, 4.830328, 4.826455, 
    4.832383, 4.842665, 4.856229, 4.869998, 4.882415, 4.891881, 4.897665, 
    4.899386, 4.899063, 4.897659, 4.900507, 4.90607, 4.916288, 4.932685, 
    4.956121, 4.986723, 5.023946, 5.066707, 5.113532, 5.16267, 5.212178, 
    5.259955, 5.303786, 5.34137, 5.370416, 5.388793, 5.394788, 5.38742, 
    5.366787,
  // height(10,44, 0-49)
    5.204635, 5.238729, 5.268057, 5.289697, 5.30149, 5.302343, 5.292276, 
    5.272214, 5.243718, 5.20869, 5.169145, 5.127045, 5.08421, 5.042264, 
    5.0026, 4.967926, 4.949046, 4.92391, 4.904885, 4.892501, 4.88643, 
    4.88929, 4.896282, 4.906398, 4.916552, 4.925547, 4.932125, 4.93589, 
    4.936687, 4.936886, 4.937493, 4.94312, 4.952159, 4.966044, 4.985777, 
    5.011779, 5.043863, 5.081303, 5.122929, 5.167236, 5.212452, 5.256604, 
    5.297564, 5.333117, 5.361072, 5.379413, 5.386541, 5.381553, 5.364513, 
    5.336632,
  // height(10,45, 0-49)
    5.179212, 5.214012, 5.246877, 5.274645, 5.294554, 5.304733, 5.304421, 
    5.293918, 5.274354, 5.247395, 5.214958, 5.179004, 5.14139, 5.103791, 
    5.067675, 5.035524, 5.016601, 4.992625, 4.973468, 4.959824, 4.951601, 
    4.951439, 4.955157, 4.961893, 4.9686, 4.974474, 4.978585, 4.980832, 
    4.981196, 4.982283, 4.985005, 4.993274, 5.005284, 5.021986, 5.043922, 
    5.071142, 5.103206, 5.139245, 5.178025, 5.218019, 5.257449, 5.294353, 
    5.326642, 5.352213, 5.369123, 5.375821, 5.371424, 5.355994, 5.330694, 
    5.29772,
  // height(10,46, 0-49)
    5.15041, 5.183906, 5.218145, 5.250115, 5.276795, 5.295731, 5.305416, 
    5.305406, 5.296213, 5.27905, 5.255547, 5.227502, 5.196701, 5.164815, 
    5.133346, 5.104626, 5.08668, 5.064239, 5.04522, 5.03049, 5.020214, 
    5.017181, 5.017759, 5.021304, 5.024827, 5.027922, 5.029962, 5.031085, 
    5.031336, 5.033477, 5.038228, 5.048871, 5.063292, 5.081979, 5.10506, 
    5.132253, 5.162891, 5.19597, 5.230196, 5.264036, 5.295753, 5.323472, 
    5.345274, 5.359347, 5.364205, 5.358969, 5.343636, 5.319263, 5.287948, 
    5.25254,
  // height(10,47, 0-49)
    5.119985, 5.150326, 5.183611, 5.217366, 5.248749, 5.275069, 5.294239, 
    5.305062, 5.307268, 5.30139, 5.288529, 5.270121, 5.247734, 5.222944, 
    5.197252, 5.1729, 5.157071, 5.136595, 5.11804, 5.102479, 5.090351, 
    5.084734, 5.082446, 5.08311, 5.083791, 5.084471, 5.08479, 5.085076, 
    5.085362, 5.088531, 5.095047, 5.107666, 5.123862, 5.143695, 5.166904, 
    5.192897, 5.220782, 5.249414, 5.27744, 5.303342, 5.32549, 5.342224, 
    5.351979, 5.353467, 5.345912, 5.329299, 5.304561, 5.273603, 5.239101, 
    5.204047,
  // height(10,48, 0-49)
    5.089595, 5.115337, 5.145545, 5.178566, 5.212147, 5.243782, 5.271115, 
    5.29231, 5.306252, 5.312603, 5.311698, 5.304386, 5.291848, 5.275453, 
    5.25664, 5.23762, 5.225192, 5.207209, 5.189566, 5.173572, 5.159956, 
    5.152224, 5.147508, 5.145734, 5.143994, 5.142636, 5.141529, 5.141139, 
    5.141435, 5.145405, 5.153227, 5.167259, 5.184483, 5.204558, 5.226863, 
    5.250508, 5.274375, 5.297177, 5.317502, 5.333895, 5.344922, 5.349295, 
    5.346019, 5.33458, 5.315123, 5.288604, 5.256801, 5.222151, 5.187412, 
    5.155191,
  // height(10,49, 0-49)
    5.053679, 5.072524, 5.096591, 5.125384, 5.157755, 5.191944, 5.225796, 
    5.257071, 5.283777, 5.304451, 5.318295, 5.325191, 5.325613, 5.320494, 
    5.311103, 5.300251, 5.299141, 5.285053, 5.268355, 5.251288, 5.235315, 
    5.227765, 5.223431, 5.222784, 5.22031, 5.217353, 5.213843, 5.210539, 
    5.206765, 5.208167, 5.214479, 5.229855, 5.247833, 5.267559, 5.287977, 
    5.307836, 5.32576, 5.340317, 5.350102, 5.353841, 5.350516, 5.339516, 
    5.320797, 5.295008, 5.263525, 5.228363, 5.191968, 5.156848, 5.125219, 
    5.098701,
  // height(11,0, 0-49)
    5.173462, 5.206308, 5.240257, 5.272574, 5.300474, 5.321579, 5.334246, 
    5.337715, 5.33208, 5.318138, 5.297173, 5.270765, 5.240604, 5.208375, 
    5.175654, 5.144077, 5.116427, 5.090436, 5.068562, 5.051296, 5.038685, 
    5.030923, 5.027062, 5.026567, 5.028524, 5.032345, 5.037494, 5.043713, 
    5.050945, 5.059712, 5.070448, 5.084126, 5.100892, 5.121141, 5.144976, 
    5.172139, 5.202004, 5.233603, 5.265666, 5.296687, 5.325003, 5.348888, 
    5.366683, 5.376942, 5.378628, 5.371307, 5.355311, 5.331816, 5.302765, 
    5.270608,
  // height(11,1, 0-49)
    5.194742, 5.228152, 5.26071, 5.289646, 5.312393, 5.32699, 5.332311, 
    5.328114, 5.314935, 5.29389, 5.266475, 5.234376, 5.199319, 5.162972, 
    5.126867, 5.092795, 5.064954, 5.037652, 5.015035, 4.997619, 4.985379, 
    4.97889, 4.976613, 4.977965, 4.981647, 4.987005, 4.993341, 5.000309, 
    5.007703, 5.0163, 5.026547, 5.039942, 5.056371, 5.076459, 5.100532, 
    5.128533, 5.160006, 5.194112, 5.229676, 5.265248, 5.299183, 5.329723, 
    5.355093, 5.373639, 5.383974, 5.385177, 5.376961, 5.359829, 5.335091, 
    5.304753,
  // height(11,2, 0-49)
    5.215133, 5.247335, 5.276393, 5.299809, 5.315543, 5.322279, 5.319528, 
    5.307566, 5.287278, 5.259983, 5.227242, 5.190721, 5.152076, 5.112883, 
    5.074576, 5.039062, 5.011899, 4.983998, 4.961249, 4.944171, 4.93268, 
    4.927715, 4.927212, 4.93057, 4.936181, 4.943317, 4.951117, 4.959096, 
    4.966879, 4.975387, 4.985026, 4.997762, 5.013227, 5.032263, 5.055445, 
    5.082962, 5.114574, 5.149624, 5.187086, 5.225627, 5.263697, 5.299596, 
    5.33156, 5.357855, 5.376884, 5.387331, 5.388323, 5.37959, 5.3616, 5.335593,
  // height(11,3, 0-49)
    5.23278, 5.262092, 5.285949, 5.302372, 5.310034, 5.308362, 5.297498, 
    5.278173, 5.251532, 5.218977, 5.182038, 5.142278, 5.101216, 5.060287, 
    5.020789, 4.984736, 4.959036, 4.931108, 4.908727, 4.892389, 4.881948, 
    4.878703, 4.880101, 4.885571, 4.893275, 4.902404, 4.911927, 4.921201, 
    4.929637, 4.9382, 4.947193, 4.959, 4.972971, 4.990158, 5.011407, 
    5.037199, 5.067567, 5.102092, 5.139944, 5.17996, 5.220726, 5.260663, 
    5.298082, 5.331253, 5.358465, 5.378115, 5.388823, 5.389595, 5.380008, 
    5.360395,
  // height(11,4, 0-49)
    5.246124, 5.271151, 5.28868, 5.297393, 5.296728, 5.286824, 5.26838, 
    5.242476, 5.21042, 5.173625, 5.133534, 5.091561, 5.049062, 5.007304, 
    4.967432, 4.931567, 4.908005, 4.880484, 4.858866, 4.843581, 4.83441, 
    4.833011, 4.836378, 4.843999, 4.853899, 4.86519, 4.876671, 4.887522, 
    4.896918, 4.905757, 4.914163, 4.924904, 4.936983, 4.951648, 4.970031, 
    4.992957, 5.020799, 5.053441, 5.090303, 5.130426, 5.172563, 5.215267, 
    5.256948, 5.295912, 5.330392, 5.358579, 5.378705, 5.389174, 5.388783, 
    5.376987,
  // height(11,5, 0-49)
    5.254175, 5.273928, 5.284616, 5.285609, 5.277045, 5.259663, 5.234583, 
    5.203132, 5.1667, 5.126667, 5.08436, 5.041042, 4.997897, 4.956021, 
    4.916396, 4.881262, 4.860361, 4.83355, 4.812981, 4.798963, 4.791189, 
    4.79168, 4.796989, 4.80671, 4.818825, 4.832373, 4.846004, 4.858711, 
    4.86942, 4.878846, 4.88686, 4.896566, 4.906542, 4.918179, 4.932914, 
    4.951959, 4.976102, 5.005606, 5.040208, 5.079185, 5.121468, 5.165733, 
    5.210474, 5.254028, 5.294588, 5.330204, 5.358836, 5.378459, 5.387281, 
    5.384035,
  // height(11,6, 0-49)
    5.256631, 5.270588, 5.274484, 5.268309, 5.25277, 5.229043, 5.198534, 
    5.162709, 5.122982, 5.080671, 5.036992, 4.993062, 4.949906, 4.90846, 
    4.869534, 4.835497, 4.817565, 4.791654, 4.772311, 4.759662, 4.753291, 
    4.755591, 4.762683, 4.77432, 4.788547, 4.804348, 4.820257, 4.835084, 
    4.847507, 4.857955, 4.865939, 4.874877, 4.882786, 4.891138, 4.901649, 
    4.915957, 4.935346, 4.960551, 4.991693, 5.028335, 5.069591, 5.114242, 
    5.160832, 5.2077, 5.252995, 5.294673, 5.33052, 5.358258, 5.375719, 
    5.381134,
  // height(11,7, 0-49)
    5.253899, 5.261981, 5.259573, 5.247164, 5.225865, 5.197128, 5.162515, 
    5.123538, 5.081592, 5.037923, 4.993641, 4.949739, 4.907105, 4.866518, 
    4.828615, 4.795863, 4.780922, 4.756021, 4.737971, 4.726662, 4.721548, 
    4.72541, 4.733949, 4.747142, 4.763211, 4.781125, 4.799346, 4.816528, 
    4.831117, 4.843144, 4.851673, 4.860385, 4.866592, 4.871735, 4.877743, 
    4.88669, 4.900416, 4.920234, 4.94675, 4.979874, 5.018923, 5.062773, 
    5.109976, 5.158839, 5.207454, 5.253706, 5.295303, 5.329849, 5.355006, 
    5.36871,
  // height(11,8, 0-49)
    5.246972, 5.249469, 5.241543, 5.224041, 5.198316, 5.165953, 5.128552, 
    5.087615, 5.044479, 5.000314, 4.956141, 4.912849, 4.871207, 4.831842, 
    4.795206, 4.763745, 4.751428, 4.727627, 4.710842, 4.700696, 4.696517, 
    4.701485, 4.710924, 4.725105, 4.742551, 4.762268, 4.782706, 4.802408, 
    4.81963, 4.83391, 4.843769, 4.853097, 4.858361, 4.860801, 4.86244, 
    4.865728, 4.873104, 4.886553, 4.907292, 4.935679, 4.971288, 5.01309, 
    5.059626, 5.109141, 5.159651, 5.208991, 5.254846, 5.29482, 5.326542, 
    5.347835,
  // height(11,9, 0-49)
    5.237248, 5.234728, 5.222235, 5.200835, 5.17199, 5.1373, 5.09833, 
    5.056515, 5.013119, 4.96924, 4.925823, 4.883679, 4.843467, 4.805668, 
    4.770514, 4.740153, 4.729591, 4.707032, 4.691422, 4.682123, 4.678374, 
    4.683771, 4.693341, 4.707723, 4.725875, 4.746894, 4.769297, 4.791569, 
    4.811847, 4.829095, 4.841227, 4.852277, 4.857747, 4.858494, 4.856425, 
    4.854231, 4.854913, 4.861206, 4.875076, 4.897473, 4.92833, 4.966763, 
    5.011302, 5.060114, 5.111127, 5.162135, 5.210836, 5.254894, 5.292007, 
    5.319999,
  // height(11,10, 0-49)
    5.226325, 5.219534, 5.203464, 5.179299, 5.148501, 5.112608, 5.073096, 
    5.031306, 4.988426, 4.94549, 4.903389, 4.862872, 4.824508, 4.788627, 
    4.755206, 4.725522, 4.715262, 4.694233, 4.679683, 4.670805, 4.666822, 
    4.671776, 4.680524, 4.694141, 4.712152, 4.733792, 4.757727, 4.782455, 
    4.806074, 4.826941, 4.84233, 4.856339, 4.863483, 4.86403, 4.859515, 
    4.852623, 4.846785, 4.845483, 4.851567, 4.866756, 4.891508, 4.925184, 
    4.966353, 5.013109, 5.063296, 5.114656, 5.164914, 5.211822, 5.253187, 
    5.286903,
  // height(11,11, 0-49)
    5.215777, 5.205538, 5.186835, 5.160881, 5.129076, 5.092853, 5.05357, 
    5.01247, 4.970669, 4.929159, 4.888799, 4.850304, 4.814176, 4.780593, 
    4.749253, 4.719546, 4.70758, 4.688578, 4.67502, 4.666077, 4.661113, 
    4.664628, 4.671499, 4.683293, 4.700191, 4.72163, 4.746493, 4.773363, 
    4.800385, 4.825321, 4.844834, 4.86298, 4.873383, 4.875564, 4.870417, 
    4.860304, 4.848796, 4.840018, 4.837758, 4.844696, 4.862033, 4.889554, 
    4.925972, 4.969349, 5.01745, 5.067966, 5.118637, 5.167293, 5.211854, 
    5.250307,
  // height(11,12, 0-49)
    5.206971, 5.194101, 5.173579, 5.146593, 5.114454, 5.078471, 5.039887, 
    4.99986, 4.959449, 4.919629, 4.88126, 4.845059, 4.811492, 4.78062, 
    4.751868, 4.72114, 4.705098, 4.688858, 4.676319, 4.666856, 4.660173, 
    4.661228, 4.665177, 4.674097, 4.688881, 4.709216, 4.734272, 4.762765, 
    4.792983, 4.822137, 4.846368, 4.869545, 4.884646, 4.890373, 4.886761, 
    4.875495, 4.859918, 4.844513, 4.833935, 4.83196, 4.84078, 4.860842, 
    4.891177, 4.929914, 4.974764, 5.023362, 5.073436, 5.12287, 5.169671, 
    5.211904,
  // height(11,13, 0-49)
    5.200899, 5.186135, 5.164429, 5.136922, 5.104827, 5.069341, 5.031617, 
    4.992749, 4.953773, 4.915673, 4.879345, 4.845548, 4.814764, 4.787011, 
    4.761545, 4.728561, 4.7061, 4.693552, 4.682205, 4.671872, 4.662838, 
    4.660499, 4.66059, 4.665687, 4.677411, 4.695735, 4.72017, 4.749611, 
    4.782543, 4.815727, 4.844905, 4.873561, 4.8944, 4.905334, 4.90543, 
    4.895422, 4.878002, 4.857599, 4.839486, 4.828537, 4.828136, 4.839681, 
    4.862757, 4.895705, 4.936254, 4.981984, 5.030586, 5.079952, 5.128131, 
    5.173246,
  // height(11,14, 0-49)
    5.198095, 5.182048, 5.159592, 5.13182, 5.099866, 5.064854, 5.027873, 
    4.989992, 4.952253, 4.915678, 4.881233, 4.849756, 4.82182, 4.797526, 
    4.776157, 4.739671, 4.70902, 4.701211, 4.69137, 4.679989, 4.668147, 
    4.661624, 4.657088, 4.65757, 4.665394, 4.680862, 4.703853, 4.733477, 
    4.768441, 4.805169, 4.839162, 4.873245, 4.9003, 4.917571, 4.923186, 
    4.916782, 4.900061, 4.876922, 4.852844, 4.83361, 4.823883, 4.826264, 
    4.841175, 4.867381, 4.902731, 4.944778, 4.991159, 5.039723, 5.088521, 
    5.135692,
  // height(11,15, 0-49)
    5.198611, 5.181742, 5.158781, 5.130789, 5.098861, 5.064082, 5.027527, 
    4.990268, 4.953382, 4.917949, 4.885024, 4.855564, 4.83031, 4.809587, 
    4.793001, 4.752295, 4.712822, 4.710817, 4.702914, 4.690477, 4.67556, 
    4.664219, 4.654443, 4.649671, 4.652883, 4.664748, 4.685534, 4.714571, 
    4.750784, 4.790377, 4.82878, 4.867803, 4.900972, 4.92504, 4.93734, 
    4.936428, 4.922827, 4.899501, 4.871641, 4.845568, 4.827119, 4.820251, 
    4.826494, 4.845283, 4.874737, 4.912448, 4.955987, 5.003134, 5.051886, 
    5.100367,
  // height(11,16, 0-49)
    5.202085, 5.184723, 5.161361, 5.133057, 5.10091, 5.066013, 5.029459, 
    4.99235, 4.955808, 4.920977, 4.889006, 4.860992, 4.837896, 4.820388, 
    4.808672, 4.76449, 4.717262, 4.722044, 4.716553, 4.703173, 4.685042, 
    4.668344, 4.652804, 4.642239, 4.640246, 4.647893, 4.665833, 4.693597, 
    4.730288, 4.771996, 4.814262, 4.857442, 4.896148, 4.926826, 4.946223, 
    4.951967, 4.943392, 4.922285, 4.893093, 4.862197, 4.836313, 4.820743, 
    4.818316, 4.829373, 4.852494, 4.885402, 4.925627, 4.970856, 5.019004, 
    5.068143,
  // height(11,17, 0-49)
    5.207882, 5.190274, 5.166554, 5.137811, 5.105181, 5.069798, 5.032796, 
    4.995312, 4.95851, 4.923584, 4.891758, 4.864257, 4.842258, 4.826826, 
    4.818871, 4.77463, 4.723094, 4.735348, 4.732672, 4.718445, 4.696949, 
    4.674356, 4.652512, 4.635655, 4.627968, 4.630945, 4.645575, 4.671546, 
    4.708066, 4.751193, 4.796754, 4.843171, 4.886521, 4.923114, 4.949328, 
    4.962093, 4.959697, 4.942693, 4.914481, 4.881027, 4.849508, 4.826371, 
    4.815795, 4.819218, 4.835872, 4.863728, 4.900331, 4.943276, 4.990375, 
    5.039623,
  // height(11,18, 0-49)
    5.215275, 5.197681, 5.173691, 5.144443, 5.111129, 5.074939, 5.037043, 
    4.998607, 4.960812, 4.924872, 4.892043, 4.863613, 4.840909, 4.825321, 
    4.818491, 4.781203, 4.73237, 4.751977, 4.752251, 4.737044, 4.711777, 
    4.682581, 4.653769, 4.630121, 4.616386, 4.614459, 4.625572, 4.649482, 
    4.685395, 4.729392, 4.777759, 4.826488, 4.873441, 4.914927, 4.947153, 
    4.966595, 4.970727, 4.958978, 4.933579, 4.899727, 4.8646, 4.835458, 
    4.817726, 4.814026, 4.824396, 4.847192, 4.880045, 4.920485, 4.966215, 
    5.015142,
  // height(11,19, 0-49)
    5.223647, 5.206471, 5.182448, 5.152765, 5.118663, 5.081373, 5.042089, 
    5.001988, 4.962242, 4.924037, 4.888577, 4.857102, 4.830956, 4.811839, 
    4.802468, 4.782428, 4.748799, 4.774101, 4.776849, 4.759989, 4.72988, 
    4.692934, 4.656215, 4.62528, 4.605374, 4.598666, 4.606437, 4.628368, 
    4.663541, 4.708077, 4.758886, 4.809097, 4.858589, 4.903782, 4.940869, 
    4.966106, 4.976411, 4.9703, 4.948884, 4.916395, 4.87963, 4.846251, 
    4.822695, 4.812732, 4.817303, 4.835267, 4.864427, 4.902291, 4.94647, 
    4.994776,
  // height(11,20, 0-49)
    5.228605, 5.209377, 5.183713, 5.153066, 5.118945, 5.08285, 5.046243, 
    5.010551, 4.977164, 4.947405, 4.922451, 4.903156, 4.889757, 4.881487, 
    4.876232, 0, 4.74619, 4.746288, 4.737542, 4.720608, 4.697607, 4.668127, 
    4.638677, 4.612827, 4.595506, 4.58938, 4.596458, 4.617135, 4.651025, 
    4.694868, 4.746641, 4.79661, 4.846766, 4.893705, 4.933717, 4.963015, 
    4.978206, 4.977147, 4.959987, 4.929938, 4.893122, 4.857208, 4.829299, 
    4.814166, 4.813659, 4.827224, 4.852918, 4.888282, 4.930861, 4.978384,
  // height(11,21, 0-49)
    5.2353, 5.216488, 5.190962, 5.160259, 5.125952, 5.089577, 5.052596, 
    5.016393, 4.982272, 4.951435, 4.92492, 4.903454, 4.887238, 4.875626, 
    4.866798, 0, 4.797721, 4.792305, 4.77688, 4.75208, 4.720561, 4.678942, 
    4.639472, 4.605354, 4.581752, 4.571404, 4.576097, 4.595869, 4.629888, 
    4.674782, 4.72919, 4.780305, 4.832267, 4.881819, 4.925358, 4.959108, 
    4.979494, 4.983882, 4.97161, 4.944922, 4.909168, 4.871809, 4.840419, 
    4.820678, 4.815356, 4.824558, 4.846657, 4.879263, 4.919861, 4.966089,
  // height(11,22, 0-49)
    5.239971, 5.221348, 5.19583, 5.165015, 5.130526, 5.093925, 5.056665, 
    5.020096, 4.985459, 4.95387, 4.926275, 4.903344, 4.885296, 4.871654, 
    4.860947, 0, 4.835303, 4.825794, 4.806291, 4.777096, 4.740961, 4.690882, 
    4.644479, 4.604306, 4.575753, 4.561767, 4.564087, 4.582548, 4.615982, 
    4.660958, 4.716836, 4.767711, 4.819979, 4.870557, 4.915993, 4.952604, 
    4.976768, 4.985557, 4.977713, 4.954643, 4.920895, 4.883494, 4.850173, 
    4.82724, 4.818252, 4.823944, 4.84304, 4.873272, 4.912107, 4.957114,
  // height(11,23, 0-49)
    5.242476, 5.223934, 5.198411, 5.167542, 5.132972, 5.096276, 5.058898, 
    5.022161, 4.987256, 4.95525, 4.927035, 4.903254, 4.884159, 4.869406, 
    4.857812, 0, 4.860757, 4.848539, 4.826694, 4.795172, 4.756673, 4.700799, 
    4.649669, 4.605175, 4.572934, 4.556139, 4.556563, 4.573909, 4.606749, 
    4.651597, 4.708432, 4.75862, 4.810601, 4.861441, 4.90783, 4.9462, 
    4.97295, 4.984998, 4.980686, 4.960799, 4.929197, 4.892447, 4.858245, 
    4.833289, 4.82172, 4.824795, 4.841565, 4.869889, 4.907241, 4.951149,
  // height(11,24, 0-49)
    5.242755, 5.224256, 5.198783, 5.167976, 5.133484, 5.096869, 5.059566, 
    5.022881, 4.987978, 4.955898, 4.927505, 4.903431, 4.883943, 4.868771, 
    4.856884, 0, 4.873823, 4.860311, 4.837456, 4.80504, 4.765738, 4.706779, 
    4.653216, 4.606438, 4.572193, 4.55386, 4.553253, 4.570012, 4.602548, 
    4.647337, 4.704798, 4.75439, 4.805976, 4.856723, 4.903411, 4.942552, 
    4.970578, 4.984347, 4.981996, 4.963964, 4.933707, 4.897477, 4.862895, 
    4.836847, 4.823806, 4.825346, 4.840734, 4.867923, 4.904401, 4.947665,
  // height(11,25, 0-49)
    5.240794, 5.22232, 5.196975, 5.166369, 5.132127, 5.095788, 5.058773, 
    5.022375, 4.987755, 4.955944, 4.927806, 4.903964, 4.884675, 4.869664, 
    4.8579, 0, 4.873703, 4.860322, 4.837665, 4.805562, 4.766716, 4.707583, 
    4.654046, 4.607269, 4.572984, 4.554605, 4.553962, 4.570693, 4.603181, 
    4.647916, 4.705504, 4.754699, 4.80592, 4.856369, 4.902862, 4.941946, 
    4.970081, 4.984127, 4.982181, 4.964595, 4.934705, 4.898656, 4.864019, 
    4.837709, 4.824278, 4.825392, 4.84038, 4.86723, 4.903439, 4.946502,
  // height(11,26, 0-49)
    5.236609, 5.218122, 5.192966, 5.162689, 5.128861, 5.092988, 5.056469, 
    5.020595, 4.98654, 4.955349, 4.927902, 4.904818, 4.886321, 4.872047, 
    4.860817, 0, 4.860604, 4.848742, 4.827468, 4.796851, 4.759639, 4.703284, 
    4.652233, 4.607754, 4.575406, 4.558476, 4.558778, 4.576014, 4.608685, 
    4.653347, 4.710508, 4.75958, 4.810529, 4.860532, 4.90638, 4.944607, 
    4.971689, 4.984544, 4.981393, 4.962756, 4.932151, 4.895843, 4.8614, 
    4.835618, 4.82288, 4.824695, 4.8403, 4.867644, 4.904226, 4.947563,
  // height(11,27, 0-49)
    5.230247, 5.211652, 5.186687, 5.156816, 5.12353, 5.088286, 5.052456, 
    5.017334, 4.984122, 4.953905, 4.927598, 4.90583, 4.888774, 4.875917, 
    4.8658, 0, 4.835612, 4.826562, 4.807929, 4.780112, 4.745865, 4.695104, 
    4.648843, 4.608716, 4.580005, 4.565769, 4.567803, 4.585944, 4.618935, 
    4.663445, 4.719617, 4.768734, 4.819421, 4.868762, 4.913473, 4.950031, 
    4.97492, 4.985185, 4.979329, 4.958301, 4.926076, 4.889226, 4.855335, 
    4.83092, 4.819949, 4.823555, 4.84074, 4.869361, 4.906916, 4.950954,
  // height(11,28, 0-49)
    5.221816, 5.202913, 5.178044, 5.148566, 5.115879, 5.081367, 5.046379, 
    5.012208, 4.980105, 4.951216, 4.926524, 4.906692, 4.891847, 4.881296, 
    4.873246, 0, 4.800921, 4.795757, 4.781104, 4.757642, 4.728002, 4.685359, 
    4.64586, 4.611671, 4.58779, 4.577054, 4.5813, 4.600579, 4.633968, 
    4.678254, 4.733004, 4.782204, 4.832494, 4.880813, 4.923745, 4.957682, 
    4.979128, 4.985353, 4.975339, 4.950729, 4.91621, 4.878789, 4.846007, 
    4.823902, 4.815784, 4.822229, 4.841906, 4.872549, 4.91166, 4.956846,
  // height(11,29, 0-49)
    5.211528, 5.191969, 5.166947, 5.13771, 5.105555, 5.071788, 5.037718, 
    5.004653, 4.97389, 4.946674, 4.924098, 4.906909, 4.895241, 4.888247, 
    4.883862, 0, 4.758096, 4.757624, 4.74851, 4.73148, 4.7087, 4.676564, 
    4.645609, 4.618504, 4.600053, 4.593021, 4.59944, 4.61967, 4.653188, 
    4.696864, 4.749561, 4.798358, 4.847646, 4.894192, 4.934445, 4.964732, 
    4.981649, 4.982831, 4.967932, 4.939481, 4.902971, 4.865784, 4.835213, 
    4.816581, 4.812366, 4.8225, 4.845302, 4.8784, 4.919327, 4.965767,
  // height(11,30, 0-49)
    5.203184, 5.185256, 5.161644, 5.13331, 5.101258, 5.066503, 5.030076, 
    4.993026, 4.956442, 4.921446, 4.889181, 4.860801, 4.837526, 4.82086, 
    4.81322, 4.793564, 4.759291, 4.783369, 4.786592, 4.771524, 4.744068, 
    4.707412, 4.671654, 4.641252, 4.621176, 4.613644, 4.620066, 4.640306, 
    4.673593, 4.716428, 4.766704, 4.814546, 4.862028, 4.905797, 4.942236, 
    4.967708, 4.97907, 4.974526, 4.954614, 4.922864, 4.885518, 4.850087, 
    4.823308, 4.809544, 4.810329, 4.82495, 4.851427, 4.887334, 4.930273, 
    4.978027,
  // height(11,31, 0-49)
    5.191897, 5.173043, 5.149139, 5.121112, 5.08991, 5.056485, 5.021814, 
    4.986914, 4.952852, 4.920757, 4.891789, 4.867128, 4.847923, 4.835331, 
    4.830701, 4.793941, 4.74672, 4.765321, 4.765812, 4.751783, 4.728415, 
    4.699248, 4.671027, 4.647578, 4.633379, 4.630328, 4.639804, 4.661777, 
    4.695667, 4.737928, 4.785717, 4.832349, 4.877781, 4.918511, 4.950845, 
    4.971227, 4.976875, 4.966708, 4.942261, 4.908067, 4.87096, 4.838338, 
    4.81617, 4.807773, 4.813767, 4.832868, 4.862859, 4.901292, 4.945847, 
    4.994394,
  // height(11,32, 0-49)
    5.182117, 5.162619, 5.138494, 5.110645, 5.079966, 5.047355, 5.013735, 
    4.980078, 4.947419, 4.916849, 4.889486, 4.866421, 4.848642, 4.836962, 
    4.832007, 4.788759, 4.739945, 4.751895, 4.749567, 4.736239, 4.716129, 
    4.69341, 4.671788, 4.654728, 4.646223, 4.647764, 4.660519, 4.684406, 
    4.718903, 4.760376, 4.805366, 4.850052, 4.892422, 4.928905, 4.955868, 
    4.970041, 4.969263, 4.95342, 4.925176, 4.889977, 4.854934, 4.826926, 
    4.810857, 4.808888, 4.820767, 4.844739, 4.87844, 4.919459, 4.965571, 
    5.014742,
  // height(11,33, 0-49)
    5.174572, 5.154589, 5.13018, 5.102248, 5.071674, 5.039321, 5.00607, 
    4.972849, 4.940649, 4.910503, 4.883449, 4.860447, 4.842265, 4.829318, 
    4.82152, 4.779136, 4.735283, 4.740807, 4.736142, 4.723701, 4.706699, 
    4.689884, 4.674292, 4.663169, 4.660039, 4.665985, 4.681876, 4.707491, 
    4.742249, 4.782453, 4.824167, 4.866026, 4.904251, 4.935326, 4.955851, 
    4.96308, 4.955732, 4.934846, 4.90422, 4.869962, 4.83904, 4.817427, 
    4.808751, 4.814018, 4.832221, 4.861261, 4.898711, 4.942233, 4.989711, 
    5.039204,
  // height(11,34, 0-49)
    5.170084, 5.149796, 5.125022, 5.096713, 5.065773, 5.033074, 4.999493, 
    4.965929, 4.933328, 4.902668, 4.874899, 4.850855, 4.831088, 4.815667, 
    4.803902, 4.766072, 4.730641, 4.730635, 4.724333, 4.713195, 4.699438, 
    4.68818, 4.678235, 4.672667, 4.674529, 4.684519, 4.703167, 4.730061, 
    4.764484, 4.802741, 4.840598, 4.878656, 4.91169, 4.936383, 4.949773, 
    4.949892, 4.936552, 4.912015, 4.881037, 4.849986, 4.825233, 4.811538, 
    4.81119, 4.824152, 4.848831, 4.882911, 4.923972, 4.969772, 5.0183, 
    5.067683,
  // height(11,35, 0-49)
    5.16936, 5.149054, 5.123928, 5.095007, 5.063273, 5.029659, 4.99507, 
    4.960418, 4.926631, 4.894642, 4.865333, 4.839435, 4.817364, 4.798974, 
    4.783234, 4.750862, 4.725138, 4.7207, 4.713482, 4.704073, 4.693744, 
    4.687737, 4.683125, 4.682759, 4.689171, 4.702719, 4.723572, 4.751113, 
    4.784435, 4.819942, 4.853301, 4.886603, 4.913572, 4.931258, 4.937376, 
    4.930943, 4.912982, 4.886868, 4.857957, 4.832395, 4.815557, 4.810833, 
    4.819266, 4.839981, 4.870982, 4.909855, 4.954227, 5.001952, 5.051094, 
    5.099827,
  // height(11,36, 0-49)
    5.172808, 5.152929, 5.127627, 5.098027, 5.065219, 5.030244, 4.994094, 
    4.95773, 4.922098, 4.888113, 4.856624, 4.828312, 4.803537, 4.782102, 
    4.762949, 4.735329, 4.718907, 4.711125, 4.703607, 4.696209, 4.689353, 
    4.688214, 4.688584, 4.693012, 4.703455, 4.719961, 4.742342, 4.769779, 
    4.801148, 4.833087, 4.861357, 4.889116, 4.909484, 4.920085, 4.919499, 
    4.907862, 4.887349, 4.862151, 4.837749, 4.819602, 4.811847, 4.816537, 
    4.833683, 4.861814, 4.898704, 4.941922, 4.989157, 5.038332, 5.08755, 
    5.134997,
  // height(11,37, 0-49)
    5.180398, 5.161556, 5.136457, 5.106329, 5.072402, 5.035862, 4.997823, 
    4.959341, 4.921418, 4.884993, 4.850913, 4.819863, 4.792229, 4.767898, 
    4.746009, 4.72179, 4.713002, 4.702868, 4.695462, 4.6901, 4.686528, 
    4.689706, 4.694558, 4.703251, 4.717091, 4.735848, 4.758998, 4.785535, 
    4.814129, 4.841794, 4.864573, 4.886342, 4.900098, 4.904203, 4.898227, 
    4.883398, 4.862806, 4.841026, 4.823173, 4.813704, 4.815465, 4.829372, 
    4.854675, 4.889541, 4.931647, 4.978592, 5.028115, 5.07816, 5.126826, 
    5.172269,
  // height(11,38, 0-49)
    5.191592, 5.174534, 5.150224, 5.119972, 5.085162, 5.047144, 5.007191, 
    4.966487, 4.926123, 4.887098, 4.850299, 4.816452, 4.786022, 4.759057, 
    4.735008, 4.712789, 4.70924, 4.697576, 4.690451, 4.686867, 4.686113, 
    4.692836, 4.701461, 4.713706, 4.730173, 4.750387, 4.773516, 4.798402, 
    4.82355, 4.846487, 4.86371, 4.879532, 4.88728, 4.886151, 4.876693, 
    4.861042, 4.842818, 4.826513, 4.816519, 4.816159, 4.827136, 4.849496, 
    4.882006, 4.922656, 4.969118, 5.019029, 5.070147, 5.120387, 5.167787, 
    5.210437,
  // height(11,39, 0-49)
    5.205347, 5.190912, 5.168145, 5.138416, 5.103247, 5.064161, 5.022605, 
    4.979915, 4.937297, 4.895839, 4.856494, 4.820059, 4.787104, 4.757856, 
    4.732081, 4.710703, 4.709868, 4.697269, 4.690359, 4.688056, 4.689408, 
    4.698699, 4.710176, 4.72507, 4.743271, 4.764093, 4.786444, 4.809061, 
    4.830353, 4.848471, 4.860497, 4.870972, 4.873897, 4.869296, 4.858545, 
    4.844366, 4.830497, 4.82097, 4.819266, 4.827655, 4.846931, 4.876558, 
    4.915043, 4.960332, 5.010135, 5.06212, 5.114024, 5.163682, 5.209023, 
    5.248034,
  // height(11,40, 0-49)
    5.220186, 5.209238, 5.188896, 5.160541, 5.125803, 5.086365, 5.043848, 
    4.999744, 4.955394, 4.911988, 4.870568, 4.832009, 4.796983, 4.765884, 
    4.73874, 4.717393, 4.717087, 4.703911, 4.69698, 4.695314, 4.697904, 
    4.708665, 4.721914, 4.738419, 4.75739, 4.777978, 4.798889, 4.81882, 
    4.836173, 4.849782, 4.857394, 4.863602, 4.863284, 4.857172, 4.847208, 
    4.836345, 4.828079, 4.825771, 4.831997, 4.848148, 4.874382, 4.90982, 
    4.95287, 5.001508, 5.053501, 5.106535, 5.158285, 5.206468, 5.248866, 
    5.283354,
  // height(11,41, 0-49)
    5.23431, 5.227661, 5.210699, 5.184736, 5.151451, 5.112651, 5.070111, 
    5.025473, 4.980214, 4.935633, 4.892861, 4.852852, 4.816367, 4.783926, 
    4.755749, 4.733974, 4.732622, 4.719017, 4.711739, 4.710033, 4.712957, 
    4.724083, 4.737983, 4.755019, 4.773808, 4.793388, 4.812348, 4.829412, 
    4.84305, 4.852812, 4.85709, 4.860407, 4.858553, 4.852761, 4.845245, 
    4.838876, 4.836684, 4.841298, 4.854504, 4.87704, 4.908657, 4.948308, 
    4.994401, 5.044983, 5.097881, 5.150779, 5.201279, 5.246957, 5.285442, 
    5.314502,
  // height(11,42, 0-49)
    5.245757, 5.244094, 5.231469, 5.209024, 5.178406, 5.141475, 5.100114, 
    5.056091, 5.011003, 4.966255, 4.923054, 4.882427, 4.845201, 4.811985, 
    4.783129, 4.76075, 4.75743, 4.7434, 4.735441, 4.733069, 4.735492, 
    4.745985, 4.759491, 4.776057, 4.793811, 4.811748, 4.828418, 4.84264, 
    4.853035, 4.859815, 4.861965, 4.863824, 4.861996, 4.857988, 4.854019, 
    4.852657, 4.856369, 4.867102, 4.886012, 4.913383, 4.948726, 4.99094, 
    5.038484, 5.089493, 5.141856, 5.193256, 5.241224, 5.283213, 5.316723, 
    5.33947,
  // height(11,43, 0-49)
    5.252583, 5.256382, 5.248981, 5.231237, 5.20464, 5.171007, 5.132254, 
    5.090226, 5.046606, 5.002879, 4.96032, 4.92001, 4.882821, 4.849424, 
    4.820261, 4.797302, 4.791629, 4.777101, 4.768164, 4.764614, 4.765842, 
    4.774894, 4.787142, 4.802403, 4.818435, 4.834261, 4.848473, 4.860041, 
    4.867776, 4.872492, 4.873652, 4.875337, 4.87478, 4.873552, 4.873688, 
    4.877326, 4.886364, 4.902164, 4.925396, 4.95604, 4.993475, 5.036603, 
    5.083958, 5.133768, 5.18399, 5.232327, 5.276277, 5.313229, 5.340635, 
    5.356261,
  // height(11,44, 0-49)
    5.253074, 5.262515, 5.261069, 5.249179, 5.228035, 5.199276, 5.164745, 
    5.12628, 5.085594, 5.044218, 5.003467, 4.964456, 4.928098, 4.895112, 
    4.866016, 4.842618, 4.834599, 4.819472, 4.809327, 4.804217, 4.803734, 
    4.810767, 4.821117, 4.834463, 4.848287, 4.861711, 4.873432, 4.882618, 
    4.888287, 4.891765, 4.892875, 4.89539, 4.896967, 4.89908, 4.90345, 
    4.911751, 4.925344, 4.945101, 4.971322, 5.003768, 5.041742, 5.084168, 
    5.129661, 5.176544, 5.222858, 5.266371, 5.304625, 5.335056, 5.355216, 
    5.363077,
  // height(11,45, 0-49)
    5.245976, 5.260865, 5.26584, 5.260825, 5.246549, 5.224311, 5.19573, 
    5.162527, 5.126361, 5.08875, 5.05102, 5.014307, 4.97956, 4.947553, 
    4.918889, 4.895254, 4.885153, 4.869344, 4.85784, 4.850928, 4.848397, 
    4.853063, 4.861111, 4.872155, 4.883486, 4.894375, 4.903677, 4.910774, 
    4.914892, 4.917789, 4.919525, 4.923557, 4.927764, 4.933413, 4.941857, 
    4.954303, 4.971632, 4.994293, 5.02229, 5.055206, 5.092278, 5.13245, 
    5.174401, 5.216556, 5.257073, 5.293852, 5.324604, 5.34698, 5.358833, 
    5.358551,
  // height(11,46, 0-49)
    5.230698, 5.250425, 5.261923, 5.264531, 5.258378, 5.244246, 5.223355, 
    5.197155, 5.167138, 5.134735, 5.101245, 5.067813, 5.035434, 5.004955, 
    4.977088, 4.953472, 4.941727, 4.925207, 4.912287, 4.903466, 4.898721, 
    4.900876, 4.90643, 4.914997, 4.923724, 4.932077, 4.939089, 4.944373, 
    4.94734, 4.950113, 4.952881, 4.958815, 4.965834, 4.974938, 4.987098, 
    5.003079, 5.023328, 5.047932, 5.076622, 5.108816, 5.143669, 5.180115, 
    5.216885, 5.252507, 5.285301, 5.313405, 5.334856, 5.347742, 5.35046, 
    5.342037,
  // height(11,47, 0-49)
    5.207477, 5.23103, 5.248695, 5.259253, 5.262141, 5.257459, 5.24584, 
    5.228285, 5.205985, 5.18019, 5.152124, 5.122934, 5.093671, 5.065282, 
    5.03861, 5.015327, 5.00253, 4.985361, 4.971079, 4.96038, 4.953408, 
    4.953086, 4.956131, 4.962209, 4.968366, 4.974279, 4.979176, 4.982888, 
    4.984988, 4.987902, 4.991867, 4.999817, 5.009564, 5.021826, 5.037194, 
    5.056029, 5.07839, 5.104032, 5.132427, 5.162814, 5.194239, 5.225595, 
    5.255641, 5.283024, 5.306286, 5.323929, 5.334507, 5.336784, 5.329955, 
    5.313877,
  // height(11,48, 0-49)
    5.177426, 5.203481, 5.226476, 5.244749, 5.257052, 5.262691, 5.261548, 
    5.253999, 5.240782, 5.222868, 5.201346, 5.177341, 5.151967, 5.126286, 
    5.101289, 5.078762, 5.06565, 5.04801, 5.03255, 5.020142, 5.011084, 
    5.008462, 5.009127, 5.012832, 5.016562, 5.020209, 5.023188, 5.025537, 
    5.026949, 5.030105, 5.035226, 5.045074, 5.057245, 5.072175, 5.090107, 
    5.111032, 5.134658, 5.16043, 5.187572, 5.215123, 5.242, 5.267024, 
    5.288981, 5.30666, 5.318905, 5.324718, 5.323361, 5.314494, 5.298303, 
    5.275572,
  // height(11,49, 0-49)
    5.130487, 5.157133, 5.184359, 5.21029, 5.233043, 5.250996, 5.26301, 
    5.268517, 5.267499, 5.260395, 5.247995, 5.231311, 5.211483, 5.189702, 
    5.167173, 5.146682, 5.140685, 5.122538, 5.104847, 5.089356, 5.0769, 
    5.074059, 5.074942, 5.079597, 5.082418, 5.084044, 5.083921, 5.082497, 
    5.079126, 5.079224, 5.082874, 5.095003, 5.110043, 5.128022, 5.148745, 
    5.171737, 5.196276, 5.221437, 5.24613, 5.269165, 5.289305, 5.305318, 
    5.316079, 5.32065, 5.318389, 5.309089, 5.293078, 5.271255, 5.245065, 
    5.216325,
  // height(12,0, 0-49)
    5.283156, 5.303393, 5.315825, 5.319623, 5.31465, 5.301387, 5.280786, 
    5.254111, 5.222781, 5.188264, 5.151982, 5.115261, 5.079288, 5.045088, 
    5.013504, 4.985375, 4.962522, 4.942296, 4.926528, 4.915215, 4.908121, 
    4.905272, 4.90585, 4.909438, 4.915286, 4.922814, 4.93137, 4.940413, 
    4.949502, 4.958674, 4.967987, 4.978175, 4.989471, 5.002637, 5.018452, 
    5.037585, 5.060488, 5.087313, 5.117883, 5.15169, 5.18792, 5.225489, 
    5.263074, 5.299156, 5.332043, 5.359944, 5.381062, 5.393738, 5.396669, 
    5.389134,
  // height(12,1, 0-49)
    5.289672, 5.306209, 5.313846, 5.31217, 5.301459, 5.28255, 5.256652, 
    5.225194, 5.189679, 5.15159, 5.112332, 5.073187, 5.035285, 4.999592, 
    4.966884, 4.938138, 4.916506, 4.896032, 4.880301, 4.86932, 4.862805, 
    4.861174, 4.863127, 4.868292, 4.875661, 4.884639, 4.894459, 4.904496, 
    4.91414, 4.923573, 4.932739, 4.942745, 4.953437, 4.965678, 4.980408, 
    4.998491, 5.020582, 5.047031, 5.077825, 5.112586, 5.150586, 5.19079, 
    5.231888, 5.272332, 5.310356, 5.344034, 5.371366, 5.390417, 5.399523, 
    5.397548,
  // height(12,2, 0-49)
    5.289351, 5.301156, 5.303457, 5.296273, 5.280246, 5.256473, 5.226311, 
    5.191248, 5.152781, 5.112347, 5.071281, 5.030792, 4.991937, 4.955608, 
    4.922512, 4.893762, 4.873818, 4.853418, 4.837952, 4.827422, 4.821506, 
    4.821013, 4.824201, 4.830774, 4.839534, 4.849892, 4.860994, 4.872135, 
    4.882534, 4.892459, 4.901697, 4.911676, 4.921791, 4.932947, 4.946202, 
    4.962606, 4.983036, 5.008065, 5.037891, 5.072294, 5.110664, 5.152039, 
    5.195147, 5.238437, 5.280128, 5.318251, 5.350725, 5.375486, 5.390674, 
    5.394858,
  // height(12,3, 0-49)
    5.282612, 5.289087, 5.285932, 5.273549, 5.252862, 5.225129, 5.191766, 
    5.154241, 5.113979, 5.072326, 5.030522, 4.989674, 4.950751, 4.914566, 
    4.881744, 4.85353, 4.835714, 4.815639, 4.800602, 4.790585, 4.785224, 
    4.785729, 4.789946, 4.797691, 4.807655, 4.819279, 4.831649, 4.843991, 
    4.855368, 4.866057, 4.875648, 4.885847, 4.895519, 4.905539, 4.917031, 
    4.931207, 4.949178, 4.971781, 4.999463, 5.032219, 5.069589, 5.110712, 
    5.154368, 5.199042, 5.24297, 5.2842, 5.320669, 5.350304, 5.37118, 5.381702,
  // height(12,4, 0-49)
    5.270433, 5.271401, 5.263016, 5.245987, 5.221428, 5.190666, 5.15511, 
    5.116154, 5.07512, 5.033241, 4.991632, 4.951296, 4.9131, 4.877757, 
    4.845793, 4.818586, 4.803279, 4.783717, 4.769216, 4.759707, 4.754789, 
    4.756079, 4.761035, 4.769634, 4.780541, 4.793252, 4.806829, 4.820447, 
    4.833023, 4.844786, 4.855074, 4.865842, 4.87534, 4.884321, 4.893908, 
    4.905432, 4.92024, 4.93947, 4.963875, 4.993721, 5.02876, 5.068261, 
    5.111091, 5.155785, 5.200624, 5.243716, 5.283067, 5.316677, 5.342657, 
    5.359342,
  // height(12,5, 0-49)
    5.254186, 5.249829, 5.236703, 5.215734, 5.188132, 5.155237, 5.118395, 
    5.078903, 5.037965, 4.996687, 4.956069, 4.916993, 4.880211, 4.84632, 
    4.815726, 4.789899, 4.777379, 4.758461, 4.744543, 4.735467, 4.730793, 
    4.732566, 4.737878, 4.74691, 4.758401, 4.771935, 4.786589, 4.801508, 
    4.815494, 4.828657, 4.840042, 4.851838, 4.861586, 4.869823, 4.877574, 
    4.886226, 4.897335, 4.912361, 4.932431, 4.958163, 4.989584, 5.026161, 
    5.066878, 5.110339, 5.154894, 5.19872, 5.239929, 5.276628, 5.30701, 
    5.329417,
  // height(12,6, 0-49)
    5.235466, 5.226234, 5.209022, 5.184886, 5.155065, 5.120851, 5.083508, 
    5.044224, 5.004089, 4.964089, 4.925107, 4.88791, 4.853123, 4.821205, 
    4.792401, 4.768209, 4.758565, 4.740386, 4.727033, 4.718237, 4.713521, 
    4.715374, 4.720548, 4.729478, 4.741088, 4.755076, 4.770578, 4.786751, 
    4.802309, 4.817187, 4.830103, 4.84348, 4.854072, 4.862099, 4.868368, 
    4.874223, 4.881364, 4.891574, 4.906406, 4.926915, 4.953505, 4.985915, 
    5.023302, 5.064378, 5.107562, 5.151116, 5.193247, 5.232182, 5.266211, 
    5.293715,
  // height(12,7, 0-49)
    5.215919, 5.202434, 5.181869, 5.155337, 5.124051, 5.089231, 5.052039, 
    5.013558, 4.974773, 4.936571, 4.899731, 4.864904, 4.832586, 4.803066, 
    4.776391, 4.753929, 4.746964, 4.729606, 4.716753, 4.708011, 4.702882, 
    4.704314, 4.708754, 4.716944, 4.728096, 4.742053, 4.758061, 4.775326, 
    4.792534, 4.809388, 4.824256, 4.839813, 4.851985, 4.860579, 4.86606, 
    4.869582, 4.872879, 4.878002, 4.88695, 4.901301, 4.921952, 4.949025, 
    4.981931, 5.019534, 5.060344, 5.102702, 5.144898, 5.185256, 5.222154, 
    5.254018,
  // height(12,8, 0-49)
    5.197084, 5.180053, 5.15687, 5.128651, 5.096552, 5.0617, 5.02516, 
    4.987918, 4.950877, 4.914841, 4.880503, 4.848413, 4.818925, 4.792144, 
    4.76786, 4.747036, 4.742175, 4.725766, 4.713326, 4.70436, 4.698389, 
    4.698829, 4.701871, 4.708604, 4.71863, 4.731961, 4.748012, 4.766073, 
    4.784878, 4.803852, 4.82102, 4.839316, 4.853869, 4.863999, 4.869711, 
    4.871802, 4.871869, 4.872107, 4.874922, 4.882471, 4.896258, 4.916928, 
    4.944264, 4.977354, 5.014838, 5.055129, 5.096582, 5.137584, 5.17657, 
    5.212003,
  // height(12,9, 0-49)
    5.180264, 5.160401, 5.13527, 5.105958, 5.07355, 5.03908, 5.003524, 
    4.967793, 4.932725, 4.899067, 4.86745, 4.838332, 4.811933, 4.788154, 
    4.766489, 4.747004, 4.743248, 4.728023, 4.715933, 4.706465, 4.699218, 
    4.698076, 4.699035, 4.70357, 4.711748, 4.723778, 4.739289, 4.757714, 
    4.777895, 4.798965, 4.818629, 4.840088, 4.857762, 4.870472, 4.877666, 
    4.879622, 4.877593, 4.873718, 4.870685, 4.871213, 4.877508, 4.890886, 
    4.911653, 4.939244, 4.972483, 5.00987, 5.049802, 5.090693, 5.131, 5.169196,
  // height(12,10, 0-49)
    5.166411, 5.144372, 5.117849, 5.087887, 5.0555, 5.021643, 4.987225, 
    4.9531, 4.920068, 4.888845, 4.86002, 4.833982, 4.810833, 4.790262, 
    4.771456, 4.752806, 4.748785, 4.735146, 4.723433, 4.713244, 4.704352, 
    4.701074, 4.699321, 4.700947, 4.706553, 4.716559, 4.730864, 4.749084, 
    4.770245, 4.79319, 4.815342, 4.840149, 4.861498, 4.877731, 4.887707, 
    4.891069, 4.888515, 4.881875, 4.873897, 4.867746, 4.866354, 4.871841, 
    4.885215, 4.906405, 4.934523, 4.968196, 5.005853, 5.045899, 5.086775, 
    5.126939,
  // height(12,11, 0-49)
    5.156057, 5.132392, 5.104886, 5.074547, 5.042329, 5.009131, 4.975822, 
    4.943227, 4.912133, 4.883249, 4.85715, 4.83418, 4.814344, 4.797164, 
    4.781535, 4.763055, 4.757185, 4.745727, 4.734569, 4.723561, 4.712773, 
    4.706907, 4.701915, 4.700012, 4.70236, 4.709619, 4.721997, 4.739341, 
    4.760933, 4.785336, 4.809756, 4.837816, 4.863089, 4.883525, 4.89742, 
    4.90373, 4.902445, 4.894832, 4.883407, 4.871558, 4.862848, 4.860272, 
    4.865705, 4.879758, 4.901966, 4.931159, 4.965813, 5.004309, 5.045033, 
    5.086396,
  // height(12,12, 0-49)
    5.149285, 5.12441, 5.096178, 5.065566, 5.033495, 5.000843, 4.968459, 
    4.937173, 4.907782, 4.881011, 4.857444, 4.837414, 4.820879, 4.807252, 
    4.795251, 4.776213, 4.766981, 4.758471, 4.748212, 4.73646, 4.723689, 
    4.714914, 4.706287, 4.700346, 4.698822, 4.702633, 4.712355, 4.728104, 
    4.74946, 4.774756, 4.801041, 4.831972, 4.861088, 4.886032, 4.904624, 
    4.915174, 4.916892, 4.910286, 4.897347, 4.881368, 4.866335, 4.856068, 
    4.853416, 4.859857, 4.875521, 4.899554, 4.930533, 4.966812, 5.006703, 
    5.048541,
  // height(12,13, 0-49)
    5.145769, 5.119963, 5.09112, 5.060205, 5.028135, 4.995795, 4.964047, 
    4.933748, 4.905724, 4.880737, 4.859405, 4.842088, 4.828754, 4.818828, 
    4.811018, 4.790828, 4.777141, 4.772433, 4.763588, 4.751352, 4.736684, 
    4.724803, 4.712266, 4.701881, 4.695943, 4.695662, 4.70202, 4.715442, 
    4.735847, 4.761384, 4.789021, 4.822229, 4.854795, 4.884152, 4.90777, 
    4.923401, 4.929517, 4.925776, 4.913407, 4.895278, 4.875484, 4.858485, 
    4.848105, 4.846823, 4.855548, 4.87389, 4.900612, 4.934071, 4.9725, 5.01414,
  // height(12,14, 0-49)
    5.144871, 5.118295, 5.088853, 5.057521, 5.02524, 4.992924, 4.961475, 
    4.931789, 4.904742, 4.881144, 4.861664, 4.846729, 4.836396, 4.830227, 
    4.827164, 4.805708, 4.787249, 4.787188, 4.780379, 4.768078, 4.751752, 
    4.736667, 4.720029, 4.704872, 4.694035, 4.689069, 4.691406, 4.701812, 
    4.720558, 4.745669, 4.774117, 4.808887, 4.844282, 4.877623, 4.906136, 
    4.927167, 4.938556, 4.939137, 4.929252, 4.911079, 4.888462, 4.866208, 
    4.848984, 4.840306, 4.842016, 4.854346, 4.876366, 4.906497, 4.942909, 
    4.983748,
  // height(12,15, 0-49)
    5.145796, 5.118527, 5.088447, 5.056561, 5.023852, 4.991281, 4.959796, 
    4.930346, 4.903856, 4.881192, 4.863095, 4.850088, 4.842387, 4.839818, 
    4.841783, 4.819959, 4.797536, 4.802824, 4.798692, 4.786848, 4.769209, 
    4.750873, 4.72998, 4.709755, 4.693579, 4.683396, 4.681126, 4.687901, 
    4.70434, 4.728413, 4.75718, 4.792764, 4.83025, 4.866904, 4.899821, 
    4.926082, 4.943048, 4.948842, 4.942933, 4.92663, 4.903234, 4.877543, 
    4.854808, 4.839509, 4.834488, 4.840753, 4.857808, 4.884229, 4.918171, 
    4.957691,
  // height(12,16, 0-49)
    5.14775, 5.119838, 5.089086, 5.056542, 5.023234, 4.99017, 4.958349, 
    4.928762, 4.902383, 4.88013, 4.862822, 4.851107, 4.845402, 4.84588, 
    4.852536, 4.832886, 4.808788, 4.819836, 4.818934, 4.808081, 4.789505, 
    4.767872, 4.742556, 4.716972, 4.695046, 4.67918, 4.671813, 4.674458, 
    4.688052, 4.710579, 4.739286, 4.774993, 4.813807, 4.852983, 4.889573, 
    4.920512, 4.942851, 4.954165, 4.953143, 4.940207, 4.917892, 4.890668, 
    4.864047, 4.843275, 4.83217, 4.832603, 4.844646, 4.867138, 4.898277, 
    4.936063,
  // height(12,17, 0-49)
    5.150093, 5.121617, 5.090219, 5.056981, 5.022968, 4.989228, 4.956792, 
    4.926682, 4.899899, 4.877413, 4.860113, 4.84878, 4.844049, 4.846456, 
    4.856596, 4.843801, 4.822259, 4.838977, 4.841652, 4.832212, 4.813004, 
    4.787975, 4.758004, 4.726743, 4.698685, 4.676764, 4.663949, 4.662121, 
    4.672501, 4.693131, 4.72155, 4.756793, 4.796225, 4.837117, 4.876529, 
    4.911358, 4.938486, 4.955118, 4.959318, 4.950685, 4.930918, 4.903908, 
    4.875101, 4.850234, 4.833983, 4.829096, 4.836311, 4.854834, 4.882985, 
    4.918743,
  // height(12,18, 0-49)
    5.152446, 5.123583, 5.091654, 5.057766, 5.023003, 4.988423, 4.955067, 
    4.923962, 4.896122, 4.872548, 4.854192, 4.841951, 4.836679, 4.839291, 
    4.851016, 4.851833, 4.839601, 4.861182, 4.867465, 4.859635, 4.839867, 
    4.81117, 4.776155, 4.738822, 4.704293, 4.676091, 4.657684, 4.651282, 
    4.65831, 4.676892, 4.704975, 4.739322, 4.778765, 4.820615, 4.861983, 
    4.8998, 4.930897, 4.952261, 4.961515, 4.957573, 4.941316, 4.915917, 
    4.886491, 4.85898, 4.838706, 4.829237, 4.832021, 4.846715, 4.871841, 
    4.905409,
  // height(12,19, 0-49)
    5.154763, 5.125841, 5.093623, 5.059199, 5.023643, 4.987998, 4.95329, 
    4.920535, 4.890742, 4.864912, 4.844035, 4.829114, 4.82127, 4.821993, 
    4.833523, 4.855882, 4.862566, 4.887558, 4.897141, 4.890828, 4.870145, 
    4.837114, 4.796288, 4.752288, 4.710979, 4.67649, 4.652683, 4.64197, 
    4.645842, 4.66249, 4.690382, 4.723572, 4.762553, 4.804698, 4.847201, 
    4.887078, 4.921197, 4.946469, 4.960234, 4.960886, 4.948586, 4.925761, 
    4.897009, 4.868209, 4.845094, 4.831927, 4.83085, 4.842024, 4.864239, 
    4.895589,
  // height(12,20, 0-49)
    5.154693, 5.1242, 5.09093, 5.056166, 5.021146, 4.987069, 4.955105, 
    4.926386, 4.901967, 4.88274, 4.869288, 4.861674, 4.859224, 4.860402, 
    4.862944, 0, 4.887241, 4.889175, 4.884861, 4.87331, 4.854144, 4.824542, 
    4.78899, 4.749675, 4.711314, 4.677715, 4.653001, 4.640221, 4.641569, 
    4.655976, 4.682993, 4.71405, 4.751464, 4.792706, 4.835068, 4.875674, 
    4.911485, 4.939419, 4.956679, 4.961297, 4.952844, 4.933036, 4.905849, 
    4.876883, 4.852042, 4.836103, 4.831837, 4.839926, 4.859478, 4.888717,
  // height(12,21, 0-49)
    5.155864, 5.125593, 5.092457, 5.057732, 5.02263, 4.988307, 4.955864, 
    4.926349, 4.90071, 4.879722, 4.863865, 4.853156, 4.846985, 4.843976, 
    4.841977, 0, 4.928431, 4.928067, 4.921334, 4.906662, 4.883474, 4.84574, 
    4.802858, 4.756638, 4.712227, 4.67375, 4.64543, 4.630235, 4.630127, 
    4.64397, 4.671875, 4.702372, 4.7396, 4.78107, 4.82414, 4.866025, 
    4.903787, 4.934397, 4.954999, 4.963388, 4.958678, 4.941965, 4.916625, 
    4.887901, 4.861739, 4.843331, 4.83602, 4.841007, 4.857741, 4.884601,
  // height(12,22, 0-49)
    5.156168, 5.126009, 5.092949, 5.05825, 5.023098, 4.988604, 4.955816, 
    4.925714, 4.899168, 4.876884, 4.859283, 4.846379, 4.837635, 4.831826, 
    4.826962, 0, 4.95737, 4.955109, 4.947015, 4.931, 4.906226, 4.863213, 
    4.81588, 4.765259, 4.716686, 4.674536, 4.643195, 4.62569, 4.623909, 
    4.63674, 4.664946, 4.694184, 4.7305, 4.771442, 4.814431, 4.856776, 
    4.895633, 4.928053, 4.951179, 4.962662, 4.96128, 4.947614, 4.924472, 
    4.896675, 4.870069, 4.850082, 4.840516, 4.843034, 4.857418, 4.882221,
  // height(12,23, 0-49)
    5.155862, 5.125789, 5.092804, 5.058161, 5.023019, 4.988459, 4.955489, 
    4.925042, 4.897942, 4.874845, 4.856148, 4.84187, 4.831531, 4.824033, 
    4.817537, 0, 4.976377, 4.972693, 4.963794, 4.947212, 4.921901, 4.875348, 
    4.825215, 4.771749, 4.720391, 4.675718, 4.642266, 4.623123, 4.620123, 
    4.632184, 4.660638, 4.688662, 4.724012, 4.764284, 4.806946, 4.849384, 
    4.888843, 4.92245, 4.947373, 4.961187, 4.962439, 4.951327, 4.930201, 
    4.903494, 4.876895, 4.855958, 4.8448, 4.845447, 4.857971, 4.881085,
  // height(12,24, 0-49)
    5.155117, 5.125144, 5.092268, 5.057733, 5.022682, 4.988179, 4.955212, 
    4.924688, 4.897405, 4.873996, 4.85484, 4.839958, 4.828905, 4.820646, 
    4.81344, 0, 4.985891, 4.981441, 4.972165, 4.95543, 4.930089, 4.881607, 
    4.830071, 4.775189, 4.722447, 4.676545, 4.642097, 4.622215, 4.618693, 
    4.630451, 4.65923, 4.686486, 4.721179, 4.760937, 4.803261, 4.84558, 
    4.885197, 4.919293, 4.945075, 4.960088, 4.962771, 4.953119, 4.93321, 
    4.907235, 4.880754, 4.85936, 4.84734, 4.846935, 4.858387, 4.880515,
  // height(12,25, 0-49)
    5.154003, 5.124162, 5.091442, 5.057076, 5.022206, 4.987893, 4.955125, 
    4.924804, 4.897723, 4.874507, 4.855525, 4.840787, 4.829843, 4.821658, 
    4.814504, 0, 4.985445, 4.981015, 4.971813, 4.955236, 4.930161, 4.881445, 
    4.829905, 4.775073, 4.722418, 4.676649, 4.642362, 4.622644, 4.61925, 
    4.63111, 4.66012, 4.687131, 4.721565, 4.761066, 4.803155, 4.84528, 
    4.884767, 4.918823, 4.94467, 4.959867, 4.962834, 4.953512, 4.933909, 
    4.908139, 4.88171, 4.860214, 4.847972, 4.847279, 4.858426, 4.880264,
  // height(12,26, 0-49)
    5.152479, 5.122794, 5.090271, 5.056139, 5.021544, 4.98756, 4.955191, 
    4.925356, 4.898864, 4.876347, 4.858164, 4.84431, 4.834285, 4.826993, 
    4.820641, 0, 4.975043, 4.971416, 4.962752, 4.946657, 4.92212, 4.874942, 
    4.824836, 4.771557, 4.72049, 4.676219, 4.64323, 4.624537, 4.621883, 
    4.634203, 4.663285, 4.690606, 4.725205, 4.764738, 4.80672, 4.848597, 
    4.887678, 4.921165, 4.946287, 4.960632, 4.962692, 4.952519, 4.932245, 
    4.906088, 4.879598, 4.858325, 4.846496, 4.846295, 4.857932, 4.880213,
  // height(12,27, 0-49)
    5.150397, 5.120863, 5.088561, 5.054716, 5.020484, 4.986965, 4.955193, 
    4.926123, 4.900596, 4.879271, 4.862515, 4.85029, 4.842027, 4.836516, 
    4.831839, 0, 4.955084, 4.952917, 4.945256, 4.930057, 4.906505, 4.862667, 
    4.815493, 4.76527, 4.717227, 4.67572, 4.645051, 4.628139, 4.626747, 
    4.639816, 4.668792, 4.696878, 4.731983, 4.77176, 4.813708, 4.855239, 
    4.893616, 4.925999, 4.949613, 4.96211, 4.962144, 4.950032, 4.928223, 
    4.901196, 4.874612, 4.853933, 4.843158, 4.844211, 4.857095, 4.880501,
  // height(12,28, 0-49)
    5.147523, 5.118073, 5.085974, 5.052443, 5.018648, 4.985715, 4.954721, 
    4.926675, 4.902474, 4.882824, 4.868122, 4.858309, 4.85273, 4.850033, 
    4.848179, 0, 4.926608, 4.926298, 4.920071, 4.906347, 4.884541, 4.845834, 
    4.803155, 4.757463, 4.713751, 4.676086, 4.648576, 4.634062, 4.63437, 
    4.648452, 4.677229, 4.706404, 4.742229, 4.782332, 4.82418, 4.865112, 
    4.902321, 4.932904, 4.95409, 4.963649, 4.960521, 4.945456, 4.921401, 
    4.893226, 4.866715, 4.847156, 4.838172, 4.84128, 4.85618, 4.881395,
  // height(12,29, 0-49)
    5.143562, 5.11403, 5.082041, 5.048799, 5.015478, 4.983227, 4.953168, 
    4.926374, 4.903827, 4.886317, 4.874309, 4.867758, 4.86593, 4.867328, 
    4.869853, 0, 4.889934, 4.891613, 4.88732, 4.875996, 4.857266, 4.825638, 
    4.789297, 4.749714, 4.711526, 4.678509, 4.654641, 4.642774, 4.644877, 
    4.659924, 4.688231, 4.718379, 4.754757, 4.794957, 4.836395, 4.876332, 
    4.911868, 4.940042, 4.958111, 4.964036, 4.957141, 4.938742, 4.912372, 
    4.883308, 4.857393, 4.839608, 4.833077, 4.838827, 4.856208, 4.883573,
  // height(12,30, 0-49)
    5.140514, 5.112536, 5.081708, 5.049011, 5.015432, 4.981946, 4.949521, 
    4.919111, 4.891653, 4.868042, 4.849143, 4.835805, 4.82899, 4.830027, 
    4.841019, 4.861464, 4.864655, 4.888956, 4.899061, 4.894265, 4.875897, 
    4.843383, 4.804152, 4.761779, 4.721758, 4.68805, 4.664435, 4.653369, 
    4.656442, 4.672151, 4.699848, 4.730855, 4.767568, 4.807538, 4.848127, 
    4.886528, 4.91977, 4.944874, 4.959198, 4.960996, 4.950107, 4.928501, 
    4.900321, 4.871173, 4.846792, 4.831698, 4.828403, 4.837403, 4.857709, 
    4.887527,
  // height(12,31, 0-49)
    5.134956, 5.106979, 5.076535, 5.044599, 5.012144, 4.980138, 4.949538, 
    4.921287, 4.896299, 4.875444, 4.859525, 4.84926, 4.845331, 4.848502, 
    4.859925, 4.859009, 4.845135, 4.865917, 4.872577, 4.866015, 4.848228, 
    4.820029, 4.786397, 4.750472, 4.717049, 4.68944, 4.671017, 4.664021, 
    4.67, 4.687367, 4.714871, 4.746837, 4.783939, 4.823677, 4.863338, 
    4.900009, 4.93064, 4.952261, 4.962398, 4.959703, 4.944641, 4.919906, 
    4.890231, 4.861438, 4.83902, 4.826921, 4.826994, 4.839206, 4.862264, 
    4.894248,
  // height(12,32, 0-49)
    5.129212, 5.101433, 5.071481, 5.040294, 5.008811, 4.97796, 4.948673, 
    4.921868, 4.898431, 4.87919, 4.864866, 4.856045, 4.853179, 4.856658, 
    4.867016, 4.852871, 4.831022, 4.847097, 4.850173, 4.841893, 4.824452, 
    4.79999, 4.771226, 4.741108, 4.713883, 4.692271, 4.679163, 4.676469, 
    4.685562, 4.704714, 4.732142, 4.764843, 4.801892, 4.840762, 4.878683, 
    4.912685, 4.939712, 4.956912, 4.96214, 4.954616, 4.93555, 4.908378, 
    4.878297, 4.851113, 4.831837, 4.823677, 4.827783, 4.84363, 4.869668, 
    4.90391,
  // height(12,33, 0-49)
    5.12343, 5.095872, 5.066374, 5.035829, 5.005118, 4.975122, 4.946723, 
    4.920801, 4.898202, 4.879708, 4.865957, 4.8574, 4.854257, 4.856545, 
    4.864198, 4.843874, 4.820434, 4.831309, 4.831038, 4.821383, 4.804472, 
    4.783561, 4.75934, 4.73466, 4.713286, 4.697415, 4.689446, 4.690929, 
    4.70299, 4.723768, 4.751048, 4.784074, 4.82048, 4.857722, 4.89301, 
    4.92337, 4.945841, 4.957834, 4.957703, 4.945395, 4.922944, 4.894461, 
    4.865391, 4.841245, 4.82632, 4.822978, 4.831672, 4.851446, 4.880571, 
    4.91704,
  // height(12,34, 0-49)
    5.118104, 5.090694, 5.0615, 5.031375, 5.001149, 4.971647, 4.943697, 
    4.918133, 4.895763, 4.877318, 4.863366, 4.854235, 4.849931, 4.850104, 
    4.854072, 4.83257, 4.811661, 4.817543, 4.81448, 4.804032, 4.788081, 
    4.770701, 4.75087, 4.731368, 4.715502, 4.705021, 4.701844, 4.707161, 
    4.721816, 4.74386, 4.770767, 4.803555, 4.838606, 4.873378, 4.905098, 
    4.930877, 4.947974, 4.954234, 4.948682, 4.932118, 4.907397, 4.87913, 
    4.852721, 4.83309, 4.823634, 4.825835, 4.8395, 4.863335, 4.895511, 
    4.934046,
  // height(12,35, 0-49)
    5.113986, 5.086621, 5.057515, 5.027502, 4.997377, 4.967923, 4.939924, 
    4.914174, 4.891447, 4.872436, 4.85766, 4.847354, 4.841359, 4.839027, 
    4.839162, 4.81933, 4.803371, 4.80494, 4.799863, 4.789345, 4.774886, 
    4.761084, 4.745565, 4.731028, 4.720322, 4.714813, 4.715966, 4.724633, 
    4.74135, 4.764152, 4.790324, 4.822191, 4.855091, 4.886513, 4.913769, 
    4.934159, 4.945316, 4.945704, 4.935174, 4.915422, 4.890007, 4.863766, 
    4.841733, 4.827977, 4.824899, 4.833127, 4.851935, 4.879796, 4.914845, 
    4.955168,
  // height(12,36, 0-49)
    5.111942, 5.084561, 5.055326, 5.025081, 4.994619, 4.964703, 4.936105, 
    4.909595, 4.885931, 4.865786, 4.849653, 4.83772, 4.829732, 4.824864, 
    4.821609, 4.804615, 4.794687, 4.792881, 4.786672, 4.776821, 4.764374, 
    4.754197, 4.742932, 4.733154, 4.727239, 4.726232, 4.731174, 4.742603, 
    4.760743, 4.7837, 4.808667, 4.838854, 4.868789, 4.896034, 4.918074, 
    4.932533, 4.937595, 4.932491, 4.91799, 4.896621, 4.872406, 4.850078, 
    4.833977, 4.827167, 4.831044, 4.845499, 4.8694, 4.901079, 4.938695, 
    4.980416,
  // height(12,37, 0-49)
    5.112801, 5.08544, 5.055923, 5.025138, 4.993912, 4.963036, 4.933292, 
    4.905466, 4.880316, 4.858521, 4.840577, 4.826664, 4.81651, 4.809246, 
    4.803285, 4.789212, 4.785302, 4.781154, 4.774646, 4.766088, 4.756061, 
    4.7495, 4.742392, 4.737138, 4.735608, 4.738574, 4.746701, 4.76024, 
    4.779102, 4.801551, 4.82479, 4.852537, 4.878767, 4.901183, 4.917546, 
    4.92596, 4.9253, 4.915676, 4.898742, 4.877671, 4.856634, 4.839904, 
    4.830922, 4.831695, 4.84272, 4.863298, 4.892019, 4.927155, 4.966915, 
    5.009552,
  // height(12,38, 0-49)
    5.117163, 5.089993, 5.060169, 5.028653, 4.996345, 4.964101, 4.932761, 
    4.903154, 4.876072, 4.852218, 4.83211, 4.815961, 4.803544, 4.794055, 
    4.786015, 4.774364, 4.77559, 4.770068, 4.763923, 4.757067, 4.749672, 
    4.746599, 4.743455, 4.742412, 4.744793, 4.75115, 4.761802, 4.776754, 
    4.795622, 4.81691, 4.837911, 4.862556, 4.884535, 4.90178, 4.912446, 
    4.915242, 4.909836, 4.897208, 4.879747, 4.860974, 4.844863, 4.834976, 
    4.833762, 4.842255, 4.86022, 4.886531, 4.919603, 4.957696, 4.999078, 
    5.042069,
  // height(12,39, 0-49)
    5.125264, 5.098615, 5.068628, 5.036368, 5.002841, 4.969013, 4.935816, 
    4.904154, 4.874874, 4.84872, 4.826249, 4.807725, 4.793006, 4.781432, 
    4.771742, 4.761746, 4.766644, 4.760505, 4.755105, 4.750071, 4.74527, 
    4.745384, 4.745862, 4.74859, 4.754327, 4.763429, 4.775914, 4.791576, 
    4.809772, 4.829317, 4.847673, 4.868758, 4.88626, 4.898421, 4.903902, 
    4.902092, 4.893451, 4.879701, 4.863706, 4.849003, 4.839085, 4.836678, 
    4.843287, 4.859147, 4.883482, 4.914883, 4.951668, 4.992102, 5.034494, 
    5.077206,
  // height(12,40, 0-49)
    5.136877, 5.111238, 5.081432, 5.048639, 5.014005, 4.978633, 4.943581, 
    4.909848, 4.878351, 4.849883, 4.825041, 4.804149, 4.787166, 4.773599, 
    4.76246, 4.753274, 4.760116, 4.753808, 4.749212, 4.745819, 4.743309, 
    4.746111, 4.749687, 4.755607, 4.764044, 4.775191, 4.788807, 4.804513, 
    4.821455, 4.83882, 4.854307, 4.871682, 4.884876, 4.892533, 4.893868, 
    4.888951, 4.878927, 4.866021, 4.853262, 4.843918, 4.840827, 4.845891, 
    4.859829, 4.882285, 4.912125, 4.94777, 4.987484, 5.029533, 5.072239, 
    5.113965,
  // height(12,41, 0-49)
    5.151308, 5.127309, 5.098226, 5.065358, 5.030005, 4.993429, 4.956825, 
    4.921301, 4.887843, 4.857288, 4.830274, 4.807172, 4.78804, 4.772555, 
    4.759991, 4.750806, 4.757907, 4.751545, 4.747518, 4.745323, 4.744565, 
    4.749381, 4.755365, 4.763759, 4.774164, 4.786629, 4.800695, 4.81586, 
    4.83112, 4.846073, 4.858711, 4.872571, 4.882043, 4.886209, 4.884839, 
    4.878588, 4.869079, 4.858769, 4.850559, 4.847245, 4.850982, 4.862956, 
    4.883301, 4.911276, 4.945533, 4.98441, 5.026139, 5.068966, 5.111191, 
    5.151146,
  // height(12,42, 0-49)
    5.167433, 5.145825, 5.118198, 5.085958, 5.05056, 5.013422, 4.975871, 
    4.939118, 4.904213, 4.872023, 4.84321, 4.818187, 4.797098, 4.779766, 
    4.765706, 4.755823, 4.761775, 4.755195, 4.751298, 4.749695, 4.749995, 
    4.756035, 4.763631, 4.773695, 4.7853, 4.798368, 4.81227, 4.826428, 
    4.839757, 4.852291, 4.862344, 4.873213, 4.879873, 4.881848, 4.879389, 
    4.873567, 4.866244, 4.859843, 4.856923, 4.859726, 4.86978, 4.887712, 
    4.91327, 4.945491, 4.982934, 5.023899, 5.066599, 5.109246, 5.150087, 
    5.187401,
  // height(12,43, 0-49)
    5.183809, 5.165433, 5.140165, 5.109489, 5.074985, 5.038198, 5.000572, 
    4.963393, 4.927755, 4.894545, 4.864434, 4.837869, 4.815063, 4.795979, 
    4.780333, 4.769211, 4.773004, 4.765872, 4.76158, 4.759906, 4.760523, 
    4.766987, 4.77537, 4.786294, 4.798351, 4.811367, 4.824594, 4.837421, 
    4.848752, 4.859057, 4.866989, 4.875616, 4.880549, 4.881706, 4.879692, 
    4.875801, 4.871909, 4.870196, 4.872773, 4.881325, 4.896852, 4.919589, 
    4.94904, 4.984147, 5.023449, 5.065253, 5.107759, 5.149135, 5.187568, 
    5.22127,
  // height(12,44, 0-49)
    5.198803, 5.184547, 5.162685, 5.134711, 5.102264, 5.066974, 5.03035, 
    4.993721, 4.9582, 4.924677, 4.893834, 4.866149, 4.841905, 4.821187, 
    4.803893, 4.791168, 4.792223, 4.784158, 4.778965, 4.776611, 4.77686, 
    4.783025, 4.79144, 4.802482, 4.814332, 4.826746, 4.838907, 4.85022, 
    4.859634, 4.868042, 4.874416, 4.881635, 4.88592, 4.887495, 4.887174, 
    4.886299, 4.886583, 4.889843, 4.897708, 4.911355, 4.931366, 4.957692, 
    4.989709, 5.026331, 5.066129, 5.10744, 5.148468, 5.187353, 5.222224, 
    5.251262,
  // height(12,45, 0-49)
    5.210752, 5.201502, 5.184183, 5.160196, 5.131147, 5.098663, 5.064255, 
    5.029252, 4.994759, 4.961669, 4.930681, 4.902313, 4.876929, 4.854733, 
    4.835791, 4.821271, 4.819385, 4.810057, 4.803559, 4.800041, 4.799366, 
    4.804659, 4.81249, 4.82304, 4.834153, 4.845552, 4.856387, 4.866125, 
    4.873801, 4.880695, 4.886077, 4.892675, 4.897229, 4.900172, 4.9024, 
    4.905163, 4.909904, 4.918032, 4.9307, 4.948648, 4.972125, 5.000875, 
    5.034193, 5.071006, 5.109934, 5.149368, 5.187541, 5.222595, 5.252655, 
    5.275915,
  // height(12,46, 0-49)
    5.218122, 5.214686, 5.20306, 5.184418, 5.160201, 5.131918, 5.101005, 
    5.068739, 5.036206, 5.004301, 4.973755, 4.945153, 4.91895, 4.895483, 
    4.874975, 4.858628, 4.853901, 4.843082, 4.835012, 4.830008, 4.828019, 
    4.832044, 4.838839, 4.848449, 4.858446, 4.868553, 4.87793, 4.886125, 
    4.892288, 4.898044, 4.902914, 4.909524, 4.915015, 4.919935, 4.925162, 
    4.93177, 4.940877, 4.953484, 4.970314, 4.991725, 5.017685, 5.047775, 
    5.081226, 5.116975, 5.153697, 5.189855, 5.223742, 5.253561, 5.277506, 
    5.293887,
  // height(12,47, 0-49)
    5.21968, 5.222688, 5.21781, 5.205827, 5.18786, 5.16517, 5.139026, 
    5.110605, 5.080956, 5.050987, 5.021486, 4.993125, 4.966475, 4.942011, 
    4.920112, 4.902047, 4.89479, 4.88238, 4.87262, 4.865965, 4.86244, 
    4.86497, 4.870446, 4.87882, 4.88747, 4.896142, 4.904027, 4.910778, 
    4.91566, 4.9206, 4.925312, 4.932374, 4.939193, 4.946368, 4.954691, 
    4.965012, 4.978126, 4.994638, 5.014892, 5.038917, 5.066428, 5.09685, 
    5.129348, 5.162853, 5.19609, 5.227598, 5.255783, 5.278975, 5.295548, 
    5.304067,
  // height(12,48, 0-49)
    5.214645, 5.224436, 5.227116, 5.222918, 5.212476, 5.196669, 5.176497, 
    5.152991, 5.127141, 5.099882, 5.07207, 5.044486, 5.017835, 4.992734, 
    4.969724, 4.950169, 4.940837, 4.926858, 4.91543, 4.907111, 4.90198, 
    4.902931, 4.906935, 4.913908, 4.921101, 4.9283, 4.934745, 4.940191, 
    4.944019, 4.94839, 4.953168, 4.960919, 4.969209, 4.978634, 4.989865, 
    5.003521, 5.020082, 5.039804, 5.062685, 5.088459, 5.11661, 5.146403, 
    5.176918, 5.207063, 5.235599, 5.261165, 5.28232, 5.297623, 5.305756, 
    5.305692,
  // height(12,49, 0-49)
    5.192284, 5.210041, 5.222421, 5.228807, 5.229014, 5.22324, 5.211989, 
    5.195982, 5.176065, 5.153151, 5.128168, 5.102034, 5.075628, 5.049784, 
    5.025281, 5.004552, 5.000236, 4.983833, 4.969202, 4.957649, 4.949624, 
    4.951151, 4.956371, 4.96534, 4.972784, 4.978915, 4.982822, 4.984548, 
    4.983208, 4.98358, 4.985592, 4.994268, 5.004465, 5.016714, 5.031483, 
    5.049073, 5.069549, 5.092734, 5.118204, 5.145324, 5.173291, 5.201159, 
    5.227886, 5.252362, 5.273417, 5.289875, 5.300619, 5.304664, 5.301308, 
    5.290269,
  // height(13,0, 0-49)
    5.302906, 5.297866, 5.283644, 5.261401, 5.232627, 5.198957, 5.162014, 
    5.123312, 5.084203, 5.045848, 5.009209, 4.975058, 4.943973, 4.916348, 
    4.892391, 4.872317, 4.857236, 4.844203, 4.834624, 4.828238, 4.824745, 
    4.82422, 4.826094, 4.830255, 4.836333, 4.844073, 4.853085, 4.862946, 
    4.873157, 4.88348, 4.893552, 4.903595, 4.913329, 4.923114, 4.933573, 
    4.945522, 4.959881, 4.977537, 4.999209, 5.025342, 5.056015, 5.090916, 
    5.129323, 5.170135, 5.211916, 5.252959, 5.291361, 5.325141, 5.352355, 
    5.371239,
  // height(13,1, 0-49)
    5.28951, 5.280722, 5.263025, 5.237669, 5.206186, 5.170209, 5.131349, 
    5.091095, 5.05077, 5.011506, 4.974237, 4.939699, 4.908432, 4.880779, 
    4.856899, 4.837128, 4.823848, 4.810921, 4.801519, 4.795393, 4.792206, 
    4.792432, 4.795098, 4.800194, 4.807179, 4.81584, 4.825731, 4.836394, 
    4.847203, 4.858047, 4.868423, 4.878859, 4.888578, 4.897897, 4.907441, 
    4.918092, 4.930884, 4.946864, 4.966928, 4.991677, 5.021327, 5.055649, 
    5.093979, 5.135242, 5.178015, 5.220617, 5.26118, 5.297764, 5.328457, 
    5.351484,
  // height(13,2, 0-49)
    5.270072, 5.257787, 5.237234, 5.209664, 5.176543, 5.139416, 5.099804, 
    5.059119, 5.018622, 4.979402, 4.942351, 4.90817, 4.877359, 4.850216, 
    4.826835, 4.807679, 4.796417, 4.78367, 4.774438, 4.768469, 4.765407, 
    4.766132, 4.769279, 4.774964, 4.782534, 4.791835, 4.802403, 4.813765, 
    4.825194, 4.836684, 4.847581, 4.858711, 4.868759, 4.877928, 4.886779, 
    4.896184, 4.907245, 4.921134, 4.938916, 4.961381, 4.988906, 5.021394, 
    5.058273, 5.098534, 5.14082, 5.18352, 5.224868, 5.263035, 5.29622, 
    5.322726,
  // height(13,3, 0-49)
    5.246368, 5.230927, 5.208125, 5.179145, 5.145323, 5.108055, 5.068716, 
    5.028602, 4.988883, 4.950584, 4.914549, 4.881436, 4.851695, 4.825564, 
    4.803069, 4.78479, 4.775711, 4.763161, 4.754032, 4.748058, 4.744871, 
    4.745768, 4.749006, 4.754856, 4.762612, 4.77221, 4.783199, 4.795122, 
    4.807179, 4.819442, 4.831099, 4.843277, 4.85408, 4.863536, 4.872057, 
    4.880424, 4.889727, 4.901223, 4.916138, 4.935462, 4.959786, 4.989203, 
    5.023292, 5.061168, 5.10159, 5.143067, 5.183972, 5.222636, 5.257412, 
    5.286727,
  // height(13,4, 0-49)
    5.220337, 5.202127, 5.177616, 5.147886, 5.114111, 5.077507, 5.039276, 
    5.000571, 4.962453, 4.925858, 4.89157, 4.860184, 4.83209, 4.80745, 
    4.786195, 4.768989, 4.762178, 4.749801, 4.740659, 4.734465, 4.730842, 
    4.731516, 4.734381, 4.73989, 4.747362, 4.756843, 4.767935, 4.780223, 
    4.792881, 4.806018, 4.818665, 4.832267, 4.844315, 4.854602, 4.863307, 
    4.871026, 4.878742, 4.887725, 4.899331, 4.91477, 4.934896, 4.960064, 
    4.990092, 5.024294, 5.061602, 5.100693, 5.140108, 5.178351, 5.21394, 
    5.245433,
  // height(13,5, 0-49)
    5.193888, 5.173308, 5.147536, 5.117548, 5.084359, 5.048999, 5.012493, 
    4.975842, 4.939978, 4.905743, 4.873834, 4.84477, 4.818851, 4.796136, 
    4.776439, 4.760425, 4.755842, 4.743599, 4.734304, 4.72764, 4.723233, 
    4.723243, 4.725216, 4.729818, 4.736472, 4.745353, 4.756155, 4.768545, 
    4.781706, 4.795761, 4.809578, 4.824949, 4.838744, 4.850475, 4.860016, 
    4.867673, 4.874217, 4.880829, 4.88893, 4.899941, 4.915029, 4.9349, 
    4.959711, 4.989072, 5.022166, 5.057874, 5.094924, 5.131988, 5.167728, 
    5.200819,
  // height(13,6, 0-49)
    5.168723, 5.146162, 5.119484, 5.089571, 5.057295, 5.023526, 4.989129, 
    4.954954, 4.92181, 4.890425, 4.861399, 4.835148, 4.811861, 4.791458, 
    4.773588, 4.758794, 4.756223, 4.744107, 4.734529, 4.727149, 4.721606, 
    4.720503, 4.721052, 4.724154, 4.729415, 4.737158, 4.74721, 4.759347, 
    4.772826, 4.78774, 4.802809, 4.820201, 4.836185, 4.849976, 4.861088, 
    4.869447, 4.875493, 4.880192, 4.884932, 4.891296, 4.900784, 4.914537, 
    4.933163, 4.956684, 4.984612, 5.016095, 5.050054, 5.085308, 5.12063, 
    5.154777,
  // height(13,7, 0-49)
    5.146191, 5.122014, 5.094694, 5.065038, 5.033816, 5.001769, 4.969636, 
    4.938137, 4.907962, 4.879731, 4.853929, 4.830854, 4.810551, 4.792776, 
    4.776973, 4.763321, 4.762328, 4.750426, 4.740496, 4.732202, 4.72523, 
    4.722604, 4.721231, 4.72226, 4.725554, 4.73159, 4.740366, 4.751813, 
    4.765307, 4.780891, 4.797148, 4.816651, 4.835127, 4.851506, 4.864916, 
    4.874842, 4.881288, 4.884869, 4.886801, 4.888733, 4.892467, 4.899627, 
    4.911375, 4.928267, 4.950256, 4.976807, 5.007057, 5.039953, 5.074344, 
    5.109021,
  // height(13,8, 0-49)
    5.12719, 5.101721, 5.073936, 5.044599, 5.01441, 4.984032, 4.95411, 
    4.92527, 4.898105, 4.873127, 4.850711, 4.831019, 4.81394, 4.799034, 
    4.785518, 4.77283, 4.772757, 4.761313, 4.751078, 4.74178, 4.733187, 
    4.728723, 4.725017, 4.723469, 4.724253, 4.728013, 4.734952, 4.745189, 
    4.758284, 4.7742, 4.791411, 4.812908, 4.833974, 4.853284, 4.869596, 
    4.881938, 4.889804, 4.893339, 4.893427, 4.891637, 4.889973, 4.890526, 
    4.895082, 4.90484, 4.920309, 4.941354, 4.96736, 4.997399, 5.030363, 
    5.06504,
  // height(13,9, 0-49)
    5.112118, 5.085622, 5.057474, 5.028415, 4.999117, 4.970207, 4.94228, 
    4.915903, 4.891597, 4.869787, 4.850737, 4.834479, 4.820738, 4.808884, 
    4.7979, 4.785911, 4.785915, 4.775369, 4.765037, 4.754792, 4.744537, 
    4.73805, 4.731728, 4.727205, 4.725008, 4.725948, 4.730473, 4.738923, 
    4.7511, 4.766879, 4.784646, 4.8078, 4.831308, 4.853636, 4.873232, 
    4.888683, 4.898961, 4.903659, 4.903191, 4.898856, 4.892699, 4.88718, 
    4.884699, 4.887177, 4.895783, 4.910887, 4.932183, 4.958889, 4.989927, 
    5.024058,
  // height(13,10, 0-49)
    5.100892, 5.073568, 5.045088, 5.016195, 4.987566, 4.959826, 4.933566, 
    4.909325, 4.887583, 4.868696, 4.852839, 4.839923, 4.829534, 4.820874, 
    4.812728, 4.801129, 4.800285, 4.791276, 4.781237, 4.770275, 4.758482, 
    4.749933, 4.740851, 4.733079, 4.727515, 4.725141, 4.726683, 4.732738, 
    4.743409, 4.758473, 4.776271, 4.800553, 4.826117, 4.851284, 4.874251, 
    4.893243, 4.906741, 4.913769, 4.914171, 4.908805, 4.899549, 4.88904, 
    4.880201, 4.875673, 4.877369, 4.886271, 4.902476, 4.925397, 4.954008, 
    4.987036,
  // height(13,11, 0-49)
    5.093023, 5.064999, 5.036164, 5.007285, 4.979065, 4.952162, 4.927186, 
    4.904684, 4.885119, 4.868808, 4.855855, 4.846086, 4.838981, 4.833637, 
    4.828726, 4.817231, 4.814683, 4.807994, 4.798809, 4.787527, 4.774482, 
    4.76396, 4.75211, 4.74093, 4.731703, 4.725581, 4.723604, 4.726661, 
    4.7352, 4.748919, 4.766147, 4.790886, 4.817931, 4.845511, 4.87165, 
    4.894293, 4.911518, 4.921821, 4.924446, 4.919686, 4.909037, 4.895079, 
    4.881061, 4.870255, 4.86534, 4.868004, 4.878853, 4.897589, 4.923282, 
    4.954648,
  // height(13,12, 0-49)
    5.087749, 5.05909, 5.029847, 5.00082, 4.972756, 4.946362, 4.92229, 
    4.901118, 4.883312, 4.869174, 4.858771, 4.851879, 4.847934, 4.846014, 
    4.844818, 4.833281, 4.828422, 4.824882, 4.817225, 4.80616, 4.792282, 
    4.779981, 4.765455, 4.75081, 4.737704, 4.727466, 4.721484, 4.720968, 
    4.72675, 4.738482, 4.754528, 4.778989, 4.806825, 4.836215, 4.865081, 
    4.891179, 4.912287, 4.926467, 4.932404, 4.92977, 4.919513, 4.903913, 
    4.886283, 4.870348, 4.859491, 4.856153, 4.861555, 4.875796, 4.898129, 
    4.927302,
  // height(13,13, 0-49)
    5.084192, 5.054919, 5.025204, 4.995886, 4.967764, 4.941601, 4.918097, 
    4.897873, 4.881418, 4.86904, 4.860798, 4.856464, 4.8555, 4.857069, 
    4.860056, 4.848661, 4.84133, 4.84169, 4.836272, 4.826051, 4.811856, 
    4.798031, 4.780994, 4.762904, 4.745772, 4.731121, 4.720706, 4.716094, 
    4.718533, 4.727675, 4.741975, 4.765423, 4.793318, 4.823824, 4.854806, 
    4.883918, 4.908742, 4.927023, 4.936974, 4.937667, 4.929421, 4.914011, 
    4.894545, 4.874947, 4.859157, 4.850342, 4.850424, 4.860008, 4.878631, 
    4.905142,
  // height(13,14, 0-49)
    5.081517, 5.05163, 5.021392, 4.991681, 4.963344, 4.937195, 4.913986, 
    4.89438, 4.878895, 4.867865, 4.861372, 4.85923, 4.860987, 4.865987, 
    4.87346, 4.863003, 4.853669, 4.858477, 4.855946, 4.847213, 4.833271, 
    4.818205, 4.798866, 4.777408, 4.756172, 4.736881, 4.721683, 4.712525, 
    4.7111, 4.717124, 4.729209, 4.750969, 4.778223, 4.809133, 4.841548, 
    4.873077, 4.901201, 4.923458, 4.937708, 4.942506, 4.937534, 4.923936, 
    4.904391, 4.882751, 4.863289, 4.849806, 4.844934, 4.849881, 4.864576, 
    4.888054,
  // height(13,15, 0-49)
    5.079049, 5.048556, 5.017774, 4.987615, 4.958967, 4.932677, 4.909543, 
    4.890262, 4.875388, 4.865291, 4.8601, 4.859703, 4.863788, 4.871943, 
    4.883821, 4.876032, 4.865983, 4.875477, 4.876322, 4.869667, 4.856545, 
    4.840522, 4.819111, 4.794412, 4.769051, 4.744977, 4.724737, 4.710681, 
    4.704965, 4.707441, 4.716984, 4.73648, 4.762472, 4.793127, 4.826293, 
    4.859575, 4.890423, 4.916268, 4.934734, 4.94397, 4.943079, 4.932546, 
    4.914461, 4.892363, 4.870615, 4.853478, 4.844249, 4.844784, 4.855497, 
    4.875701,
  // height(13,16, 0-49)
    5.076357, 5.04529, 5.013985, 4.983371, 4.954356, 4.927814, 4.90456, 
    4.885322, 4.870687, 4.861065, 4.85665, 4.857431, 4.863256, 4.873969, 
    4.889624, 4.887436, 4.878976, 4.892997, 4.897475, 4.893355, 4.881554, 
    4.864819, 4.841561, 4.813771, 4.784333, 4.755423, 4.729992, 4.710805, 
    4.700493, 4.699131, 4.705956, 4.722753, 4.746984, 4.776818, 4.810111, 
    4.844488, 4.877415, 4.906292, 4.928608, 4.942223, 4.945766, 4.939097, 
    4.923651, 4.902481, 4.879802, 4.860133, 4.84732, 4.843862, 4.850718, 
    4.867552,
  // height(13,17, 0-49)
    5.073276, 5.041718, 5.00995, 4.978906, 4.949494, 4.922585, 4.899002, 
    4.879483, 4.864644, 4.854941, 4.850645, 4.851858, 4.858593, 4.870928, 
    4.889231, 4.896774, 4.893412, 4.911368, 4.919476, 4.918165, 4.908042, 
    4.890761, 4.865815, 4.835064, 4.801618, 4.767901, 4.737255, 4.712861, 
    4.697815, 4.692492, 4.696613, 4.710435, 4.732548, 4.761121, 4.794013, 
    4.828882, 4.86324, 4.894509, 4.920127, 4.937771, 4.94571, 4.943258, 
    4.931211, 4.912036, 4.889621, 4.86853, 4.853006, 4.846128, 4.849413, 
    4.862942,
  // height(13,18, 0-49)
    5.069894, 5.037993, 5.005871, 4.974439, 4.94458, 4.917144, 4.89294, 
    4.872707, 4.857082, 4.846572, 4.841537, 4.842215, 4.848804, 4.861626, 
    4.881323, 4.903514, 4.910012, 4.930978, 4.94249, 4.944072, 4.935783, 
    4.917948, 4.891298, 4.857579, 4.820136, 4.781682, 4.745924, 4.716439, 
    4.696753, 4.687572, 4.689219, 4.699979, 4.719781, 4.746784, 4.778859, 
    4.813701, 4.848888, 4.881894, 4.910168, 4.931293, 4.943286, 4.945026, 
    4.936729, 4.920257, 4.899048, 4.877536, 4.860189, 4.850558, 4.850698, 
    4.861127,
  // height(13,19, 0-49)
    5.066533, 5.034526, 5.002198, 4.970406, 4.939985, 4.911748, 4.886477, 
    4.864903, 4.847689, 4.835394, 4.828495, 4.827422, 4.832679, 4.845, 
    4.865422, 4.907155, 4.92915, 4.952248, 4.966908, 4.971374, 4.964861, 
    4.946195, 4.917465, 4.88041, 4.838736, 4.795547, 4.754904, 4.720706, 
    4.696789, 4.684154, 4.683802, 4.691631, 4.709097, 4.734366, 4.765323, 
    4.799715, 4.83519, 4.869302, 4.899551, 4.923498, 4.939002, 4.944619, 
    4.940077, 4.926665, 4.907319, 4.886206, 4.86786, 4.856178, 4.853689, 
    4.861349,
  // height(13,20, 0-49)
    5.062326, 5.029428, 4.996673, 4.965066, 4.935573, 4.909109, 4.88653, 
    4.868585, 4.85582, 4.848474, 4.846332, 4.848631, 4.854045, 4.860835, 
    4.867209, 0, 4.960554, 4.96489, 4.966611, 4.9642, 4.956264, 4.938369, 
    4.913416, 4.881072, 4.843659, 4.803276, 4.763498, 4.72832, 4.70213, 
    4.68676, 4.684481, 4.689006, 4.70359, 4.72649, 4.755638, 4.788839, 
    4.823808, 4.858182, 4.88953, 4.915427, 4.93366, 4.942553, 4.941444, 
    4.931111, 4.913975, 4.893856, 4.875212, 4.86215, 4.857589, 4.862891,
  // height(13,21, 0-49)
    5.05939, 5.026729, 4.99416, 4.962648, 4.9331, 4.906367, 4.883225, 
    4.864333, 4.850152, 4.840854, 4.836205, 4.83551, 4.837572, 4.840788, 
    4.843318, 0, 4.988412, 4.991874, 4.992982, 4.989769, 4.980573, 4.958037, 
    4.92908, 4.892868, 4.851937, 4.808477, 4.766072, 4.728681, 4.700647, 
    4.683903, 4.681386, 4.684261, 4.697501, 4.719358, 4.747776, 4.780595, 
    4.815596, 4.850495, 4.882943, 4.910565, 4.93112, 4.942796, 4.944633, 
    4.936992, 4.921839, 4.902638, 4.883723, 4.869337, 4.862715, 4.865593,
  // height(13,22, 0-49)
    5.056715, 5.024198, 4.991746, 4.960288, 4.930684, 4.903732, 4.880151, 
    4.860536, 4.845291, 4.834549, 4.828082, 4.825235, 4.824912, 4.825584, 
    4.825378, 0, 5.007531, 5.01016, 5.010991, 5.007695, 4.998391, 4.972798, 
    4.941637, 4.903322, 4.860387, 4.814988, 4.770687, 4.731456, 4.701693, 
    4.683507, 4.680566, 4.681566, 4.693231, 4.713815, 4.741263, 4.773442, 
    4.808179, 4.843255, 4.876388, 4.905256, 4.92762, 4.941576, 4.94595, 
    4.940767, 4.927596, 4.90955, 4.890788, 4.875599, 4.867455, 4.868394,
  // height(13,23, 0-49)
    5.054629, 5.022224, 4.989868, 4.958463, 4.928839, 4.901758, 4.877898, 
    4.857814, 4.841877, 4.830197, 4.822548, 4.818313, 4.816451, 4.815497, 
    4.813565, 0, 5.020011, 5.021922, 5.022535, 5.019291, 5.010156, 4.982364, 
    4.949795, 4.910171, 4.86599, 4.819386, 4.773896, 4.733502, 4.702621, 
    4.683495, 4.680393, 4.679896, 4.690282, 4.709814, 4.73644, 4.768047, 
    4.802501, 4.837631, 4.871211, 4.900962, 4.924655, 4.940331, 4.946666, 
    4.94344, 4.931912, 4.914906, 4.89641, 4.880715, 4.871446, 4.870869,
  // height(13,24, 0-49)
    5.053342, 5.021052, 4.988799, 4.957475, 4.927895, 4.900801, 4.876853, 
    4.856582, 4.840339, 4.828224, 4.820012, 4.8151, 4.812484, 4.810732, 
    4.807968, 0, 5.026357, 5.027834, 5.028316, 5.025136, 5.016194, 4.987086, 
    4.953739, 4.913423, 4.868618, 4.821458, 4.775474, 4.734633, 4.703346, 
    4.683897, 4.680958, 4.67964, 4.689296, 4.708194, 4.734291, 4.765488, 
    4.799673, 4.834713, 4.868412, 4.898533, 4.92286, 4.939422, 4.946823, 
    4.944707, 4.934157, 4.91782, 4.899562, 4.883654, 4.873792, 4.872372,
  // height(13,25, 0-49)
    5.052937, 5.020776, 4.988652, 4.957452, 4.927993, 4.901019, 4.877185, 
    4.857019, 4.840869, 4.828824, 4.820656, 4.815761, 4.813137, 4.811367, 
    4.80859, 0, 5.026131, 5.027595, 5.028104, 5.025001, 5.016189, 4.986772, 
    4.953303, 4.912925, 4.868127, 4.821061, 4.775249, 4.73463, 4.703572, 
    4.684343, 4.681725, 4.680303, 4.68982, 4.708557, 4.734481, 4.76551, 
    4.799545, 4.834464, 4.868091, 4.898201, 4.922594, 4.939297, 4.946908, 
    4.945036, 4.934718, 4.918549, 4.900354, 4.884392, 4.874371, 4.872713,
  // height(13,26, 0-49)
    5.053365, 5.021352, 4.989378, 4.958348, 4.92909, 4.902367, 4.878851, 
    4.859085, 4.843421, 4.831948, 4.824425, 4.82023, 4.81834, 4.817324, 
    4.815344, 0, 5.019228, 5.021117, 5.02184, 5.018843, 5.010098, 4.981457, 
    4.948575, 4.908823, 4.864714, 4.818419, 4.773448, 4.7337, 4.703471, 
    4.684952, 4.682744, 4.681938, 4.691911, 4.710961, 4.737072, 4.768174, 
    4.802174, 4.836944, 4.870301, 4.900016, 4.923895, 4.939982, 4.946925, 
    4.944401, 4.933534, 4.917, 4.89867, 4.8828, 4.873055, 4.871789,
  // height(13,27, 0-49)
    5.054453, 5.022583, 4.990769, 4.959939, 4.930949, 4.904599, 4.881593, 
    4.862506, 4.847711, 4.837303, 4.831028, 4.82823, 4.827834, 4.828379, 
    4.828067, 0, 5.005809, 5.008458, 5.00954, 5.006703, 4.998044, 4.971261, 
    4.939735, 4.901355, 4.858659, 4.813832, 4.770372, 4.732119, 4.703287, 
    4.685929, 4.684206, 4.684655, 4.695604, 4.715379, 4.741986, 4.773363, 
    4.807406, 4.841971, 4.874848, 4.903781, 4.926571, 4.941309, 4.946741, 
    4.942723, 4.93059, 4.913219, 4.894607, 4.879008, 4.86998, 4.869713,
  // height(13,28, 0-49)
    5.055897, 5.024127, 4.992451, 4.961824, 4.933147, 4.907266, 4.884938, 
    4.866787, 4.853227, 4.844376, 4.839968, 4.839299, 4.841219, 4.844214, 
    4.846556, 0, 4.986444, 4.989986, 4.991482, 4.988878, 4.980467, 4.956567, 
    4.927253, 4.891089, 4.850602, 4.80798, 4.766706, 4.730566, 4.703684, 
    4.687934, 4.686851, 4.689076, 4.701419, 4.722225, 4.749526, 4.781257, 
    4.815298, 4.849463, 4.8815, 4.909118, 4.930127, 4.942695, 4.945752, 
    4.939439, 4.925432, 4.906913, 4.88804, 4.873039, 4.865275, 4.866679,
  // height(13,29, 0-49)
    5.057277, 5.025501, 4.993886, 4.963425, 4.935068, 4.909718, 4.888201, 
    4.871215, 4.859243, 4.852449, 4.850572, 4.852848, 4.858019, 4.864477, 
    4.870577, 0, 4.960837, 4.965211, 4.967146, 4.96498, 4.957272, 4.937307, 
    4.911318, 4.878489, 4.841214, 4.801627, 4.763185, 4.72964, 4.705064, 
    4.691149, 4.690714, 4.694875, 4.708726, 4.730634, 4.758652, 4.790708, 
    4.824646, 4.858231, 4.889145, 4.915062, 4.933808, 4.943669, 4.943821, 
    4.934777, 4.918635, 4.898928, 4.87997, 4.865904, 4.859822, 4.863319,
  // height(13,30, 0-49)
    5.059418, 5.028654, 4.997622, 4.96715, 4.938057, 4.911136, 4.887138, 
    4.866747, 4.850553, 4.839038, 4.832601, 4.831628, 4.836618, 4.848354, 
    4.867994, 4.90837, 4.928143, 4.951606, 4.967244, 4.973113, 4.968354, 
    4.949694, 4.92203, 4.886323, 4.846043, 4.804104, 4.764419, 4.730797, 
    4.707057, 4.694342, 4.694369, 4.700532, 4.715995, 4.739077, 4.76782, 
    4.800131, 4.833815, 4.866575, 4.896039, 4.919852, 4.935893, 4.942627, 
    4.93956, 4.927652, 4.909478, 4.888913, 4.870369, 4.857808, 4.853965, 
    4.860042,
  // height(13,31, 0-49)
    5.060282, 5.029759, 4.999126, 4.96925, 4.940992, 4.915175, 4.892564, 
    4.873836, 4.859542, 4.850095, 4.845772, 4.846765, 4.85328, 4.865714, 
    4.884841, 4.905748, 4.911053, 4.932447, 4.945031, 4.948086, 4.941575, 
    4.923994, 4.898461, 4.866093, 4.830063, 4.792876, 4.758057, 4.729052, 
    4.709362, 4.699802, 4.701348, 4.710032, 4.727447, 4.751931, 4.781534, 
    4.814127, 4.847456, 4.879147, 4.906764, 4.927947, 4.940672, 4.94366, 
    4.936833, 4.921684, 4.90129, 4.879853, 4.861801, 4.850834, 4.849262, 
    4.857854,
  // height(13,32, 0-49)
    5.060558, 5.030423, 5.000259, 4.970952, 4.943376, 4.918372, 4.896713, 
    4.879066, 4.865955, 4.857725, 4.854555, 4.856493, 4.863556, 4.875896, 
    4.894008, 4.900531, 4.896977, 4.915523, 4.924882, 4.9252, 4.916963, 
    4.900275, 4.876549, 4.847143, 4.815058, 4.782508, 4.752657, 4.728541, 
    4.713242, 4.707185, 4.710644, 4.721965, 4.741295, 4.766997, 4.797129, 
    4.829546, 4.861939, 4.891879, 4.916902, 4.9347, 4.943443, 4.94221, 
    4.931443, 4.913217, 4.891095, 4.869491, 4.85271, 4.844056, 4.845331, 
    4.856855,
  // height(13,33, 0-49)
    5.059862, 5.03015, 5.000467, 4.971692, 4.944696, 4.920317, 4.899325, 
    4.882373, 4.869952, 4.862354, 4.859664, 4.861796, 4.868586, 4.879933, 
    4.896007, 4.893321, 4.885574, 4.900522, 4.906545, 4.904282, 4.894521, 
    4.878765, 4.856861, 4.8304, 4.802221, 4.774295, 4.749418, 4.730218, 
    4.719326, 4.716811, 4.722351, 4.736221, 4.757266, 4.783872, 4.814105, 
    4.845798, 4.876605, 4.904065, 4.925737, 4.939448, 4.943662, 4.93793, 
    4.923305, 4.902457, 4.879358, 4.858486, 4.843853, 4.838239, 4.842885, 
    4.857669,
  // height(13,34, 0-49)
    5.058055, 5.028715, 4.999457, 4.971143, 4.944623, 4.920722, 4.900189, 
    4.883659, 4.871587, 4.864218, 4.861553, 4.863379, 4.869329, 4.879015, 
    4.892175, 4.88469, 4.876192, 4.887134, 4.889908, 4.885369, 4.874451, 
    4.859777, 4.839851, 4.816452, 4.79222, 4.768898, 4.748909, 4.734482, 
    4.727811, 4.728682, 4.736307, 4.752478, 4.774912, 4.802001, 4.831811, 
    4.862161, 4.890678, 4.914915, 4.93252, 4.941554, 4.94089, 4.930667, 
    4.912594, 4.889904, 4.866834, 4.847734, 4.836153, 4.834247, 4.842685, 
    4.860934,
  // height(13,35, 0-49)
    5.055274, 5.02619, 4.997241, 4.969266, 4.943089, 4.919506, 4.899241, 
    4.882901, 4.870915, 4.863482, 4.860535, 4.861737, 4.866537, 4.874239, 
    4.884109, 4.875016, 4.868087, 4.875023, 4.874868, 4.868522, 4.85693, 
    4.843543, 4.825792, 4.805592, 4.785332, 4.766533, 4.751252, 4.741336, 
    4.738557, 4.742521, 4.752098, 4.770198, 4.793586, 4.820644, 4.849438, 
    4.87777, 4.90328, 4.923584, 4.936518, 4.940488, 4.934902, 4.920564, 
    4.899837, 4.876399, 4.854555, 4.838321, 4.830633, 4.832978, 4.845473, 
    4.86724,
  // height(13,36, 0-49)
    5.051935, 5.022963, 4.994163, 4.966357, 4.940342, 4.916883, 4.896673, 
    4.880292, 4.868145, 4.860397, 4.856926, 4.857306, 4.860819, 4.866513, 
    4.873233, 4.864482, 4.860516, 4.863798, 4.861239, 4.853672, 4.841947, 
    4.830064, 4.814686, 4.797793, 4.781472, 4.767046, 4.756203, 4.750443, 
    4.751133, 4.757798, 4.76908, 4.788637, 4.812456, 4.838905, 4.86604, 
    4.891673, 4.9135, 4.929286, 4.937158, 4.935996, 4.925839, 4.908185, 
    4.885969, 4.863123, 4.843789, 4.831448, 4.828336, 4.835277, 4.851907, 
    4.87708,
  // height(13,37, 0-49)
    5.048712, 5.019714, 4.990895, 4.963061, 4.936992, 4.91342, 4.893018, 
    4.876333, 4.863755, 4.855429, 4.851202, 4.850588, 4.852764, 4.856591, 
    4.860627, 4.853176, 4.852786, 4.853034, 4.848742, 4.840593, 4.829271, 
    4.819106, 4.806266, 4.79274, 4.780269, 4.769989, 4.763242, 4.761208, 
    4.764874, 4.773776, 4.78642, 4.806883, 4.830554, 4.855775, 4.880613, 
    4.902925, 4.920528, 4.931437, 4.934191, 4.928248, 4.914334, 4.894584, 
    4.87234, 4.851547, 4.83594, 4.828331, 4.830231, 4.841869, 4.862504, 
    4.890805,
  // height(13,38, 0-49)
    5.046463, 5.017363, 4.988382, 4.960333, 4.933984, 4.910048, 4.889175, 
    4.871894, 4.858581, 4.849375, 4.84412, 4.842312, 4.843084, 4.84521, 
    4.847122, 4.841239, 4.84439, 4.842373, 4.837064, 4.828948, 4.818515, 
    4.810253, 4.800081, 4.789934, 4.781161, 4.774736, 4.771679, 4.772884, 
    4.778982, 4.789603, 4.803183, 4.82395, 4.846866, 4.87026, 4.892232, 
    4.910744, 4.923823, 4.92984, 4.927855, 4.917969, 4.901567, 4.881282, 
    4.860622, 4.843279, 4.832405, 4.830073, 4.83712, 4.853296, 4.877594, 
    4.908586,
  // height(13,39, 0-49)
    5.046107, 5.016935, 4.987735, 4.959342, 4.932527, 4.907993, 4.886375, 
    4.86819, 4.853814, 4.843393, 4.836789, 4.833525, 4.832754, 4.833261, 
    4.833495, 4.82901, 4.835154, 4.83167, 4.826, 4.818432, 4.809279, 
    4.803062, 4.795628, 4.788808, 4.783522, 4.780604, 4.780778, 4.78469, 
    4.79264, 4.804419, 4.818454, 4.838909, 4.860484, 4.881526, 4.900217, 
    4.914691, 4.92329, 4.924838, 4.918981, 4.90646, 4.889201, 4.870115, 
    4.852602, 4.839882, 4.834409, 4.837548, 4.849568, 4.869874, 4.897309, 
    4.930414,
  // height(13,40, 0-49)
    5.048494, 5.019421, 4.990073, 4.961317, 4.933938, 4.90864, 4.886052, 
    4.866689, 4.850931, 4.838945, 4.830641, 4.8256, 4.823055, 4.82189, 
    4.82068, 4.817156, 4.825377, 4.821116, 4.815586, 4.808927, 4.801313, 
    4.797197, 4.792489, 4.788867, 4.786796, 4.786984, 4.789888, 4.795939, 
    4.805148, 4.817516, 4.831503, 4.85106, 4.870792, 4.889106, 4.904329, 
    4.914861, 4.919432, 4.917396, 4.908987, 4.895493, 4.879183, 4.862983, 
    4.84994, 4.842655, 4.842869, 4.851325, 4.86787, 4.891695, 4.921583, 
    4.956109,
  // height(13,41, 0-49)
    5.05427, 5.025635, 4.996369, 4.967378, 4.939467, 4.913352, 4.889659, 
    4.868913, 4.851506, 4.837645, 4.827295, 4.820136, 4.815523, 4.812502, 
    4.809849, 4.806692, 4.81588, 4.811314, 4.806209, 4.800623, 4.794641, 
    4.79257, 4.790468, 4.789821, 4.790624, 4.793467, 4.798572, 4.806185, 
    4.816072, 4.828482, 4.841944, 4.860108, 4.877642, 4.893072, 4.90494, 
    4.911988, 4.913404, 4.909066, 4.899735, 4.887073, 4.87345, 4.861562, 
    4.85393, 4.852476, 4.858293, 4.871628, 4.892047, 4.918634, 4.950186, 
    4.985343,
  // height(13,42, 0-49)
    5.063781, 5.036088, 5.007306, 4.978371, 4.950112, 4.923259, 4.898448, 
    4.876221, 4.856994, 4.841022, 4.828345, 4.818758, 4.811777, 4.806639, 
    4.802362, 4.798909, 4.80793, 4.803259, 4.798624, 4.794068, 4.789628, 
    4.789413, 4.789672, 4.791672, 4.794939, 4.799946, 4.806708, 4.815324, 
    4.825358, 4.837329, 4.84987, 4.866296, 4.881484, 4.894133, 4.903078, 
    4.907446, 4.906895, 4.90178, 4.893241, 4.883102, 4.873612, 4.867048, 
    4.865321, 4.869707, 4.880752, 4.898339, 4.921859, 4.950371, 4.982732, 
    5.017666,
  // height(13,43, 0-49)
    5.077024, 5.050926, 5.02318, 4.994742, 4.966463, 4.939089, 4.913278, 
    4.889596, 4.868496, 4.850291, 4.835114, 4.822883, 4.813281, 4.80576, 
    4.799586, 4.79519, 4.80303, 4.798201, 4.793865, 4.790109, 4.786953, 
    4.788271, 4.790523, 4.794739, 4.799999, 4.80666, 4.814556, 4.823662, 
    4.8334, 4.84456, 4.855913, 4.87045, 4.883365, 4.893603, 4.900323, 
    4.903059, 4.901888, 4.897532, 4.891333, 4.885078, 4.880715, 4.880008, 
    4.884263, 4.894188, 4.909894, 4.931011, 4.956826, 4.986413, 5.018707, 
    5.052526,
  // height(13,44, 0-49)
    5.09363, 5.069897, 5.04386, 5.016483, 4.988629, 4.96107, 4.934496, 
    4.909508, 4.886611, 4.866188, 4.848468, 4.833498, 4.82113, 4.811025, 
    4.802682, 4.796786, 4.802666, 4.797429, 4.793074, 4.789756, 4.787496, 
    4.789924, 4.7937, 4.79963, 4.806377, 4.814182, 4.822727, 4.831895, 
    4.841009, 4.85113, 4.861181, 4.873878, 4.884815, 4.893214, 4.898576, 
    4.900804, 4.900312, 4.898042, 4.895368, 4.893885, 4.895139, 4.900371, 
    4.910341, 4.925292, 4.945001, 4.968908, 4.996238, 5.026088, 5.057459, 
    5.089253,
  // height(13,45, 0-49)
    5.112896, 5.092362, 5.068785, 5.043111, 5.016217, 4.988903, 4.961903, 
    4.935873, 4.911382, 4.88889, 4.868727, 4.851068, 4.835922, 4.823139, 
    4.812431, 4.804618, 4.808037, 4.802051, 4.79729, 4.793986, 4.792167, 
    4.79523, 4.800014, 4.807119, 4.814841, 4.823317, 4.832101, 4.841004, 
    4.8493, 4.858297, 4.867085, 4.878168, 4.887572, 4.894811, 4.899705, 
    4.902462, 4.903721, 4.904501, 4.906074, 4.909746, 4.916643, 4.927522, 
    4.942692, 4.962025, 4.985044, 5.011038, 5.039169, 5.068532, 5.098169, 
    5.127051,
  // height(13,46, 0-49)
    5.133814, 5.117327, 5.096988, 5.073705, 5.048361, 5.021798, 4.994802, 
    4.968101, 4.942336, 4.918055, 4.895684, 4.87552, 4.857718, 4.842292, 
    4.829139, 4.81916, 4.819887, 4.812812, 4.807271, 4.803571, 4.801742, 
    4.80497, 4.81025, 4.818002, 4.826226, 4.834962, 4.843659, 4.852087, 
    4.859497, 4.867418, 4.875102, 4.884908, 4.893291, 4.900041, 4.905254, 
    4.909355, 4.913095, 4.917461, 4.923537, 4.932306, 4.944498, 4.960462, 
    4.980148, 5.003146, 5.028774, 5.056185, 5.084462, 5.112659, 5.139817, 
    5.164942,
  // height(13,47, 0-49)
    5.155118, 5.143477, 5.127144, 5.10696, 5.083807, 5.058568, 5.032099, 
    5.005201, 4.978597, 4.952922, 4.928703, 4.906341, 4.886123, 4.868207, 
    4.85265, 4.840416, 4.838448, 4.830011, 4.823393, 4.818952, 4.816723, 
    4.819705, 4.825018, 4.832941, 4.841257, 4.849924, 4.85831, 4.866159, 
    4.872729, 4.879717, 4.886525, 4.895436, 4.903288, 4.910117, 4.91623, 
    4.922192, 4.928778, 4.936869, 4.947312, 4.960783, 4.977658, 4.997964, 
    5.021375, 5.047264, 5.074781, 5.102951, 5.130748, 5.157147, 5.181139, 
    5.201734,
  // height(13,48, 0-49)
    5.17534, 5.169244, 5.157641, 5.141272, 5.120998, 5.09774, 5.072417, 
    5.045903, 5.019007, 4.992444, 4.966833, 4.942678, 4.920383, 4.900235, 
    4.882427, 4.867987, 4.863477, 4.85351, 4.845624, 4.840209, 4.837288, 
    4.839696, 4.844657, 4.852349, 4.860429, 4.868786, 4.876736, 4.884, 
    4.889857, 4.896114, 4.9023, 4.910675, 4.918396, 4.925701, 4.933056, 
    4.941097, 4.950563, 4.962187, 4.976577, 4.994122, 5.014909, 5.038708, 
    5.064978, 5.092928, 5.121566, 5.149796, 5.176466, 5.200438, 5.22062, 5.236,
  // height(13,49, 0-49)
    5.18919, 5.190837, 5.186273, 5.175988, 5.160712, 5.141308, 5.11869, 
    5.09377, 5.067405, 5.04039, 5.013444, 4.987204, 4.962228, 4.938995, 
    4.917903, 4.901022, 4.900822, 4.888001, 4.877112, 4.869137, 4.864331, 
    4.86836, 4.875689, 4.886596, 4.896372, 4.905116, 4.911828, 4.916348, 
    4.917615, 4.919777, 4.922395, 4.930235, 4.938002, 4.946137, 4.955254, 
    4.966011, 4.979034, 4.994824, 5.013668, 5.035591, 5.060346, 5.087408, 
    5.116018, 5.145223, 5.173903, 5.200845, 5.22479, 5.244488, 5.258783, 
    5.266685,
  // height(14,0, 0-49)
    5.229131, 5.206501, 5.178502, 5.14638, 5.111412, 5.074858, 5.037918, 
    5.001689, 4.967128, 4.935019, 4.905952, 4.880305, 4.858244, 4.839743, 
    4.824595, 4.812624, 4.804584, 4.797328, 4.792109, 4.788625, 4.78663, 
    4.786323, 4.787329, 4.789779, 4.793612, 4.798909, 4.805624, 4.813658, 
    4.822749, 4.832749, 4.84324, 4.854219, 4.865003, 4.875406, 4.885445, 
    4.89538, 4.905724, 4.917185, 4.930576, 4.94668, 4.966119, 4.989237, 
    5.016041, 5.046188, 5.079033, 5.113686, 5.149096, 5.184103, 5.21749, 
    5.247988,
  // height(14,1, 0-49)
    5.207026, 5.182279, 5.152763, 5.119683, 5.084245, 5.047626, 5.010942, 
    4.975212, 4.941328, 4.910021, 4.881835, 4.857101, 4.835941, 4.818269, 
    4.80382, 4.79253, 4.786399, 4.779195, 4.773937, 4.770339, 4.768142, 
    4.767947, 4.769014, 4.771609, 4.775563, 4.781028, 4.787959, 4.796264, 
    4.805616, 4.816019, 4.826934, 4.838686, 4.850087, 4.860837, 4.870841, 
    4.880264, 4.889561, 4.899436, 4.910755, 4.924414, 4.941188, 4.961601, 
    4.985838, 5.013726, 5.044766, 5.078192, 5.113054, 5.148269, 5.182673, 
    5.215027,
  // height(14,2, 0-49)
    5.183304, 5.15703, 5.12666, 5.093325, 5.058139, 5.022183, 4.986475, 
    4.951942, 4.919401, 4.889516, 4.862769, 4.839439, 4.819584, 4.803053, 
    4.789515, 4.779003, 4.774808, 4.767579, 4.762142, 4.758224, 4.755566, 
    4.755175, 4.755948, 4.758294, 4.761974, 4.767229, 4.774033, 4.782334, 
    4.791769, 4.802477, 4.813826, 4.826488, 4.838775, 4.850249, 4.860665, 
    4.870028, 4.878657, 4.887173, 4.896429, 4.907394, 4.921, 4.937978, 
    4.958755, 4.983394, 5.011603, 5.042788, 5.076122, 5.110613, 5.14515, 
    5.178529,
  // height(14,3, 0-49)
    5.159269, 5.132011, 5.101366, 5.068372, 5.034046, 4.999361, 4.965226, 
    4.932481, 4.901851, 4.873924, 4.849108, 4.82761, 4.809415, 4.794293, 
    4.781828, 4.772121, 4.769814, 4.762452, 4.756672, 4.752212, 4.748813, 
    4.747893, 4.747982, 4.749643, 4.752614, 4.757233, 4.763523, 4.771494, 
    4.780782, 4.791656, 4.803401, 4.817072, 4.830497, 4.84309, 4.854418, 
    4.864275, 4.872768, 4.880341, 4.887757, 4.896002, 4.906137, 4.919126, 
    4.935688, 4.956191, 4.980619, 5.008601, 5.039472, 5.072342, 5.106161, 
    5.139763,
  // height(14,4, 0-49)
    5.136073, 5.108289, 5.077836, 5.045656, 5.012658, 4.979708, 4.947617, 
    4.91712, 4.888855, 4.863318, 4.840836, 4.821526, 4.805284, 4.791785, 
    4.780509, 4.771574, 4.771007, 4.763416, 4.75714, 4.751925, 4.747519, 
    4.745743, 4.744758, 4.745288, 4.747094, 4.75062, 4.755964, 4.763226, 
    4.772083, 4.782914, 4.794947, 4.809652, 4.824399, 4.838461, 4.851204, 
    4.862165, 4.871171, 4.878408, 4.884452, 4.890225, 4.896865, 4.905565, 
    4.917366, 4.933001, 4.952807, 4.976699, 5.004219, 5.034612, 5.066907, 
    5.099984,
  // height(14,5, 0-49)
    5.114647, 5.08669, 5.056768, 5.025724, 4.994371, 4.96347, 4.933736, 
    4.905807, 4.880225, 4.857395, 4.837543, 4.82069, 4.806624, 4.794909, 
    4.784913, 4.776653, 4.77757, 4.769712, 4.76284, 4.756712, 4.751087, 
    4.748175, 4.745767, 4.744746, 4.744943, 4.746911, 4.750852, 4.756979, 
    4.765056, 4.775557, 4.787667, 4.803314, 4.819453, 4.835233, 4.849818, 
    4.862471, 4.872696, 4.88035, 4.885726, 4.889578, 4.893041, 4.89748, 
    4.90426, 4.914527, 4.929033, 4.948059, 4.97142, 4.998543, 5.028562, 
    5.060421,
  // height(14,6, 0-49)
    5.095639, 5.06775, 5.038558, 5.008825, 4.979269, 4.950567, 4.923344, 
    4.898149, 4.875429, 4.855488, 4.838451, 4.824225, 4.812485, 4.802677, 
    4.79404, 4.786319, 4.788359, 4.780312, 4.772842, 4.76574, 4.758781, 
    4.754543, 4.750437, 4.747506, 4.745694, 4.74566, 4.747729, 4.752261, 
    4.759154, 4.768952, 4.780826, 4.797183, 4.814626, 4.832209, 4.848913, 
    4.86374, 4.875854, 4.884737, 4.890322, 4.893084, 4.894041, 4.894635, 
    4.896505, 4.901212, 4.909982, 4.923539, 4.942053, 4.9652, 4.992265, 
    5.022275,
  // height(14,7, 0-49)
    5.079382, 5.051685, 5.023293, 4.994893, 4.967136, 4.940629, 4.915915, 
    4.893468, 4.873641, 4.856643, 4.842487, 4.830967, 4.821641, 4.813837, 
    4.806674, 4.799337, 4.802044, 4.794051, 4.786124, 4.778114, 4.769837, 
    4.764191, 4.758224, 4.753119, 4.748968, 4.746531, 4.746279, 4.748741, 
    4.754, 4.762649, 4.773867, 4.790557, 4.809045, 4.82832, 4.847221, 
    4.864514, 4.879047, 4.889917, 4.896648, 4.899345, 4.898779, 4.896335, 
    4.893821, 4.893167, 4.896089, 4.903821, 4.916978, 4.935566, 4.959084, 
    4.986681,
  // height(14,8, 0-49)
    5.065872, 5.038401, 5.01076, 4.983597, 4.95751, 4.933054, 4.910717, 
    4.890898, 4.87387, 4.859747, 4.848433, 4.839616, 4.832747, 4.827052, 
    4.821545, 4.814451, 4.817304, 4.809798, 4.801712, 4.793008, 4.783563, 
    4.776557, 4.76869, 4.761254, 4.754529, 4.749352, 4.746367, 4.746292, 
    4.749443, 4.756443, 4.766504, 4.783024, 4.80213, 4.822789, 4.843732, 
    4.863547, 4.880808, 4.894256, 4.903001, 4.906718, 4.905815, 4.901471, 
    4.895508, 4.890118, 4.887469, 4.889338, 4.896865, 4.91048, 4.92997, 
    4.954655,
  // height(14,9, 0-49)
    5.054821, 5.027532, 5.000518, 4.974404, 4.949765, 4.927123, 4.906926, 
    4.889516, 4.875094, 4.863682, 4.855093, 4.848915, 4.84452, 4.841063, 
    4.837492, 4.83054, 4.83301, 4.826586, 4.818791, 4.809748, 4.799422, 
    4.791223, 4.781535, 4.77173, 4.762289, 4.754117, 4.748044, 4.744996, 
    4.74556, 4.750387, 4.75874, 4.774489, 4.79366, 4.815218, 4.837843, 
    4.859991, 4.880027, 4.896397, 4.907828, 4.913559, 4.913555, 4.908646, 
    4.9005, 4.891405, 4.883876, 4.880214, 4.88213, 4.890561, 4.905677, 
    4.927028,
  // height(14,10, 0-49)
    5.04573, 5.018534, 4.991975, 4.96668, 4.943219, 4.922101, 4.903752, 
    4.888469, 4.876389, 4.867462, 4.861423, 4.857787, 4.855875, 4.854819, 
    4.85357, 4.846726, 4.848333, 4.843694, 4.836761, 4.827849, 4.817042, 
    4.807907, 4.796583, 4.784479, 4.772281, 4.760951, 4.751504, 4.745098, 
    4.742626, 4.744754, 4.750842, 4.765165, 4.783755, 4.805612, 4.829389, 
    4.853467, 4.876074, 4.895433, 4.909956, 4.918473, 4.920488, 4.916383, 
    4.907503, 4.896041, 4.8847, 4.876213, 4.872857, 4.876142, 4.886695, 
    4.904379,
  // height(14,11, 0-49)
    5.038, 5.010782, 4.984499, 4.959789, 4.937232, 4.917344, 4.900531, 
    4.887064, 4.877037, 4.870335, 4.866637, 4.86542, 4.865989, 4.867517, 
    4.869044, 4.862404, 4.862796, 4.860651, 4.855209, 4.846973, 4.836166, 
    4.826419, 4.813724, 4.799486, 4.784587, 4.770025, 4.757013, 4.746933, 
    4.741017, 4.73996, 4.74325, 4.755486, 4.772819, 4.794303, 4.818602, 
    4.844064, 4.868836, 4.890996, 4.908724, 4.92051, 4.925418, 4.923341, 
    4.915177, 4.902844, 4.889031, 4.87675, 4.86878, 4.867208, 4.873197, 
    4.886992,
  // height(14,12, 0-49)
    5.031034, 5.003688, 4.977518, 4.953181, 4.931284, 4.912348, 4.896778, 
    4.884824, 4.876548, 4.871799, 4.870219, 4.871272, 4.8743, 4.878574, 
    4.883319, 4.877185, 4.876233, 4.87719, 4.873849, 4.866863, 4.856576, 
    4.846573, 4.832829, 4.816703, 4.799254, 4.781491, 4.764815, 4.750834, 
    4.741136, 4.736468, 4.736497, 4.746009, 4.761425, 4.781863, 4.806017, 
    4.832239, 4.858638, 4.883218, 4.904005, 4.919235, 4.927595, 4.928498, 
    4.922335, 4.910599, 4.895769, 4.880947, 4.869279, 4.863392, 4.865007, 
    4.874826,
  // height(14,13, 0-49)
    5.024333, 4.99677, 4.970584, 4.946457, 4.925018, 4.906796, 4.892203, 
    4.881479, 4.874665, 4.87159, 4.871881, 4.875025, 4.880433, 4.887527, 
    4.895803, 4.890821, 4.888721, 4.893181, 4.89245, 4.887251, 4.878012, 
    4.868104, 4.853672, 4.835969, 4.816206, 4.795377, 4.775051, 4.757049, 
    4.743318, 4.734697, 4.731096, 4.73732, 4.750211, 4.768974, 4.792344, 
    4.818688, 4.846123, 4.872623, 4.896131, 4.91471, 4.926751, 4.931248, 
    4.928075, 4.918214, 4.903775, 4.887743, 4.873465, 4.864006, 4.861628, 
    4.867535,
  // height(14,14, 0-49)
    5.017553, 4.989715, 4.963422, 4.939384, 4.918242, 4.90054, 4.88669, 
    4.876932, 4.871295, 4.869604, 4.871495, 4.876493, 4.884107, 4.893934, 
    4.905785, 4.903114, 4.900491, 4.908577, 4.910793, 4.907833, 4.900127, 
    4.890634, 4.875879, 4.856959, 4.835193, 4.811535, 4.787686, 4.765656, 
    4.747746, 4.734937, 4.727468, 4.729933, 4.739788, 4.756329, 4.778342, 
    4.804221, 4.832108, 4.85998, 4.88575, 4.90738, 4.923053, 4.931413, 
    4.931864, 4.92485, 4.912005, 4.896032, 4.880286, 4.868128, 4.8623, 
    4.864512,
  // height(14,15, 0-49)
    5.010522, 4.982379, 4.955929, 4.931895, 4.910927, 4.893575, 4.880256, 
    4.871205, 4.866455, 4.865833, 4.869004, 4.875539, 4.885052, 4.897312, 
    4.912402, 4.913854, 4.911866, 4.923392, 4.928685, 4.928277, 4.922505, 
    4.913686, 4.898948, 4.879184, 4.855774, 4.829604, 4.802463, 4.776515, 
    4.754398, 4.737293, 4.725864, 4.724226, 4.730651, 4.744537, 4.764725, 
    4.789639, 4.817448, 4.846156, 4.873679, 4.897934, 4.916968, 4.929162, 
    4.933515, 4.929967, 4.919626, 4.90479, 4.888655, 4.874717, 4.866093, 
    4.864969,
  // height(14,16, 0-49)
    5.003232, 4.974789, 4.948159, 4.924067, 4.903166, 4.886005, 4.872997, 
    4.864381, 4.860195, 4.860283, 4.864339, 4.872, 4.882958, 4.897115, 
    4.91473, 4.922801, 4.923217, 4.937708, 4.946001, 4.948301, 4.94475, 
    4.936777, 4.92233, 4.902053, 4.877351, 4.849022, 4.818892, 4.789238, 
    4.76301, 4.74164, 4.726334, 4.720396, 4.723143, 4.734078, 4.752094, 
    4.775647, 4.802935, 4.831992, 4.860762, 4.887154, 4.909132, 4.924897, 
    4.93313, 4.933318, 4.926054, 4.91317, 4.897569, 4.882729, 4.872013, 
    4.868022,
  // height(14,17, 0-49)
    4.995819, 4.967114, 4.940305, 4.916105, 4.895159, 4.878008, 4.865059, 
    4.856553, 4.85254, 4.852895, 4.857356, 4.865614, 4.877438, 4.892803, 
    4.912023, 4.929695, 4.934912, 4.951701, 4.962767, 4.967796, 4.966612, 
    4.959546, 4.945543, 4.924974, 4.899243, 4.869065, 4.836262, 4.803187, 
    4.773059, 4.747612, 4.728692, 4.718437, 4.717418, 4.725255, 4.740889, 
    4.762807, 4.789228, 4.818224, 4.84777, 4.875792, 4.900223, 4.919144, 
    4.930996, 4.934896, 4.930968, 4.920557, 4.906198, 4.891222, 4.879112, 
    4.872787,
  // height(14,18, 0-49)
    4.988537, 4.959641, 4.932666, 4.9083, 4.887167, 4.869789, 4.856569, 
    4.847752, 4.843416, 4.843479, 4.847744, 4.855983, 4.868048, 4.88397, 
    4.904027, 4.934335, 4.947203, 4.965634, 4.979208, 4.98692, 4.988139, 
    4.981914, 4.968329, 4.947478, 4.920774, 4.888891, 4.85365, 4.81746, 
    4.783762, 4.754593, 4.73253, 4.71814, 4.713455, 4.718208, 4.731387, 
    4.75151, 4.776821, 4.805424, 4.835332, 4.864502, 4.890868, 4.912439, 
    4.927494, 4.934857, 4.934252, 4.926565, 4.913923, 4.899424, 4.88655, 
    4.878451,
  // height(14,19, 0-49)
    4.981731, 4.952747, 4.925626, 4.901007, 4.879478, 4.86154, 4.847589, 
    4.837891, 4.832567, 4.831611, 4.834948, 4.842501, 4.854297, 4.870481, 
    4.891221, 4.936656, 4.959976, 4.979749, 4.995747, 5.00617, 5.009804, 
    5.004245, 4.990828, 4.969369, 4.941361, 4.907585, 4.869937, 4.830897, 
    4.794071, 4.761743, 4.73723, 4.719127, 4.711077, 4.712924, 4.723711, 
    4.741991, 4.766041, 4.793996, 4.823914, 4.853789, 4.881576, 4.90526, 
    4.923007, 4.933437, 4.93594, 4.930997, 4.920331, 4.906754, 4.893658, 
    4.88432,
  // height(14,20, 0-49)
    4.975356, 4.946013, 4.918895, 4.894783, 4.874384, 4.858284, 4.846906, 
    4.840438, 4.838765, 4.841401, 4.847481, 4.8558, 4.864954, 4.87357, 
    4.880587, 0, 4.989855, 4.995119, 5.000073, 5.003455, 5.004048, 4.997201, 
    4.985688, 4.96794, 4.944427, 4.914887, 4.880343, 4.842763, 4.805717, 
    4.771926, 4.745841, 4.724278, 4.712812, 4.711535, 4.719627, 4.735713, 
    4.758105, 4.784973, 4.814407, 4.844437, 4.873043, 4.898208, 4.918039, 
    4.931002, 4.936229, 4.933856, 4.92523, 4.912845, 4.899946, 4.889857,
  // height(14,21, 0-49)
    4.970289, 4.941153, 4.914182, 4.890114, 4.869606, 4.853193, 4.841239, 
    4.833877, 4.830952, 4.831978, 4.836136, 4.842323, 4.849247, 4.85558, 
    4.860119, 0, 5.006929, 5.011988, 5.017016, 5.020457, 5.020889, 5.011185, 
    4.997466, 4.977767, 4.952747, 4.922137, 4.886837, 4.848618, 4.81087, 
    4.776311, 4.749987, 4.726534, 4.71325, 4.710298, 4.716912, 4.731764, 
    4.753213, 4.779468, 4.808661, 4.838869, 4.868112, 4.894393, 4.915797, 
    4.930689, 4.938019, 4.937646, 4.930596, 4.919082, 4.906178, 4.895215,
  // height(14,22, 0-49)
    4.96617, 4.937153, 4.910255, 4.886184, 4.865558, 4.848874, 4.83646, 
    4.828418, 4.824572, 4.824438, 4.827231, 4.831902, 4.837212, 4.841824, 
    4.844385, 0, 5.018405, 5.023205, 5.02841, 5.032224, 5.033048, 5.021325, 
    5.00638, 4.985718, 4.960042, 4.928993, 4.893322, 4.85464, 4.816243, 
    4.780902, 4.754295, 4.728978, 4.713942, 4.709406, 4.71464, 4.728346, 
    4.748909, 4.774562, 4.803468, 4.833735, 4.863416, 4.890533, 4.913163, 
    4.929612, 4.938688, 4.940041, 4.934431, 4.923813, 4.911096, 4.899575,
  // height(14,23, 0-49)
    4.96328, 4.934348, 4.907502, 4.883425, 4.862714, 4.845841, 4.833112, 
    4.824607, 4.820145, 4.819244, 4.821142, 4.824821, 4.829068, 4.832527, 
    4.833734, 0, 5.025937, 5.030453, 5.035746, 5.039857, 5.041064, 5.027761, 
    5.011934, 4.990608, 4.964503, 4.9332, 4.897349, 4.85845, 4.819719, 
    4.783957, 4.757343, 4.730652, 4.714336, 4.708647, 4.712873, 4.725742, 
    4.745659, 4.770877, 4.799579, 4.829896, 4.859901, 4.887634, 4.911168, 
    4.928766, 4.939146, 4.941798, 4.937283, 4.927362, 4.914799, 4.902847,
  // height(14,24, 0-49)
    4.961791, 4.932945, 4.906162, 4.882113, 4.861383, 4.844429, 4.831546, 
    4.822805, 4.81802, 4.816717, 4.818145, 4.821302, 4.824994, 4.827858, 
    4.828371, 0, 5.029955, 5.034287, 5.039621, 5.043921, 5.045398, 5.031094, 
    5.014718, 4.992973, 4.966591, 4.935138, 4.899226, 4.8603, 4.821521, 
    4.785698, 4.759323, 4.731932, 4.714949, 4.708636, 4.712295, 4.724666, 
    4.744171, 4.76908, 4.797589, 4.827847, 4.857946, 4.88594, 4.909908, 
    4.928101, 4.939186, 4.942573, 4.93871, 4.929234, 4.916815, 4.904671,
  // height(14,25, 0-49)
    4.961771, 4.933026, 4.906334, 4.882361, 4.86169, 4.844777, 4.831912, 
    4.823165, 4.818351, 4.816997, 4.818359, 4.821449, 4.825079, 4.827899, 
    4.828384, 0, 5.03003, 5.034381, 5.039783, 5.044186, 5.045787, 5.031203, 
    5.014672, 4.992793, 4.966319, 4.934835, 4.89897, 4.860161, 4.821557, 
    4.785944, 4.759897, 4.732482, 4.715449, 4.709057, 4.712609, 4.724858, 
    4.744236, 4.769025, 4.797433, 4.827615, 4.857674, 4.88567, 4.909687, 
    4.927975, 4.939195, 4.942734, 4.939016, 4.929639, 4.917246, 4.905041,
  // height(14,26, 0-49)
    4.963167, 4.93454, 4.907962, 4.884112, 4.863579, 4.846827, 4.834151, 
    4.825628, 4.821076, 4.820027, 4.821736, 4.825215, 4.829287, 4.832619, 
    4.833757, 0, 5.026039, 5.030636, 5.036156, 5.040594, 5.042174, 5.028095, 
    5.011848, 4.990179, 4.963848, 4.932496, 4.896807, 4.858271, 4.820046, 
    4.784883, 4.759194, 4.73243, 4.715955, 4.710011, 4.713904, 4.726387, 
    4.745905, 4.770749, 4.799131, 4.829207, 4.85908, 4.886809, 4.91048, 
    4.928358, 4.939132, 4.942234, 4.938139, 4.928508, 4.91602, 4.903892,
  // height(14,27, 0-49)
    4.965813, 4.937301, 4.910845, 4.887145, 4.866809, 4.850321, 4.837995, 
    4.829924, 4.825934, 4.825562, 4.828056, 4.832419, 4.837465, 4.841897, 
    4.844372, 0, 5.018102, 5.023104, 5.028753, 5.033145, 5.034584, 5.021748, 
    5.006234, 4.985136, 4.959219, 4.928194, 4.892848, 4.854764, 4.817146, 
    4.782689, 4.757411, 4.731923, 4.71657, 4.711563, 4.716202, 4.729245, 
    4.749143, 4.774192, 4.802603, 4.832528, 4.862057, 4.88924, 4.912171, 
    4.929139, 4.938899, 4.940991, 4.93603, 4.925817, 4.913135, 4.901226,
  // height(14,28, 0-49)
    4.969423, 4.940984, 4.914621, 4.891065, 4.870954, 4.854809, 4.842978, 
    4.835584, 4.832475, 4.833191, 4.836968, 4.842775, 4.849395, 4.855551, 
    4.860049, 0, 5.006672, 5.0121, 5.017801, 5.022041, 5.023263, 5.01228, 
    4.997938, 4.977812, 4.952632, 4.922198, 4.887433, 4.850056, 4.81334, 
    4.779905, 4.755203, 4.731562, 4.717834, 4.714186, 4.719908, 4.733754, 
    4.754178, 4.779477, 4.80786, 4.837467, 4.866374, 4.892624, 4.914323, 
    4.929817, 4.937974, 4.938513, 4.932271, 4.921261, 4.908408, 4.896985,
  // height(14,29, 0-49)
    4.973598, 4.945132, 4.91878, 4.895313, 4.875417, 4.859663, 4.848455, 
    4.841969, 4.840096, 4.842386, 4.848045, 4.855969, 4.864852, 4.873392, 
    4.88053, 0, 4.991336, 4.997087, 5.002714, 5.006726, 5.007765, 4.999115, 
    4.986455, 4.96784, 4.943899, 4.91449, 4.880672, 4.844324, 4.808808, 
    4.776659, 4.752664, 4.731198, 4.719398, 4.717382, 4.724414, 4.739241, 
    4.760315, 4.785926, 4.81427, 4.84347, 4.871576, 4.896624, 4.916734, 
    4.930334, 4.936449, 4.935032, 4.927205, 4.915243, 4.902236, 4.891462,
  // height(14,30, 0-49)
    4.978459, 4.950448, 4.924171, 4.90026, 4.879285, 4.861737, 4.848003, 
    4.838342, 4.832888, 4.831677, 4.83469, 4.841944, 4.853562, 4.869802, 
    4.890952, 4.937116, 4.960141, 4.981357, 4.999086, 5.011297, 5.016665, 
    5.010939, 4.99806, 4.977265, 4.949973, 4.916874, 4.879813, 4.841241, 
    4.804756, 4.772696, 4.748902, 4.729621, 4.719982, 4.719895, 4.728523, 
    4.744562, 4.766439, 4.792431, 4.820715, 4.84939, 4.876489, 4.900041, 
    4.918213, 4.929551, 4.93329, 4.929682, 4.920183, 4.907356, 4.894434, 
    4.88467,
  // height(14,31, 0-49)
    4.983125, 4.955338, 4.929348, 4.905835, 4.885411, 4.868597, 4.85578, 
    4.847207, 4.842966, 4.843014, 4.847225, 4.855464, 4.867691, 4.884041, 
    4.904872, 4.935839, 4.949141, 4.969279, 4.984799, 4.994443, 4.997485, 
    4.991339, 4.978379, 4.958244, 4.932343, 4.901263, 4.86675, 4.83112, 
    4.797772, 4.768725, 4.747015, 4.731064, 4.72435, 4.726704, 4.737257, 
    4.754694, 4.777433, 4.803735, 4.831755, 4.85956, 4.885167, 4.906618, 
    4.922161, 4.930507, 4.931175, 4.92478, 4.913159, 4.899173, 4.886178, 
    4.877337,
  // height(14,32, 0-49)
    4.987358, 4.959856, 4.934148, 4.91095, 4.890905, 4.874556, 4.862307, 
    4.854393, 4.850876, 4.851655, 4.85653, 4.865274, 4.877754, 4.894031, 
    4.914469, 4.932961, 4.939357, 4.958105, 4.971329, 4.978452, 4.979202, 
    4.972534, 4.959299, 4.939528, 4.914677, 4.885373, 4.853353, 4.820845, 
    4.790998, 4.765457, 4.746442, 4.73423, 4.730731, 4.735687, 4.748199, 
    4.766947, 4.790341, 4.816634, 4.843962, 4.870373, 4.893885, 4.912594, 
    4.924883, 4.929708, 4.926944, 4.917631, 4.904008, 4.889196, 4.876601, 
    4.869208,
  // height(14,33, 0-49)
    4.99063, 4.963439, 4.938015, 4.915095, 4.895347, 4.879332, 4.867464, 
    4.859974, 4.856893, 4.858074, 4.863241, 4.872085, 4.88437, 4.900063, 
    4.919447, 4.928698, 4.931004, 4.947732, 4.958413, 4.962972, 4.961474, 
    4.954248, 4.940749, 4.921361, 4.897592, 4.870147, 4.840767, 4.811585, 
    4.785475, 4.763719, 4.747799, 4.739508, 4.739332, 4.746913, 4.761318, 
    4.78121, 4.804995, 4.83091, 4.85707, 4.88152, 4.902306, 4.917626, 
    4.926063, 4.926908, 4.920468, 4.908258, 4.892908, 4.877741, 4.866107, 
    4.860717,
  // height(14,34, 0-49)
    4.992525, 4.96564, 4.940499, 4.917854, 4.898386, 4.882666, 4.871113, 
    4.863943, 4.86116, 4.862561, 4.867793, 4.876443, 4.888147, 4.902713, 
    4.920231, 4.923387, 4.923928, 4.937998, 4.945892, 4.947875, 4.944241, 
    4.936496, 4.92287, 4.90407, 4.881607, 4.856267, 4.829761, 4.804101, 
    4.781861, 4.764022, 4.751439, 4.747082, 4.750193, 4.760307, 4.776446, 
    4.797251, 4.821106, 4.846224, 4.870707, 4.892605, 4.910032, 4.921345, 
    4.92542, 4.921961, 4.911783, 4.896895, 4.880278, 4.865354, 4.855299, 
    4.852454,
  // height(14,35, 0-49)
    4.99278, 4.96617, 4.941314, 4.91896, 4.899793, 4.884388, 4.873153, 
    4.866287, 4.863753, 4.865289, 4.87046, 4.87873, 4.889587, 4.902627, 
    4.917654, 4.917314, 4.917788, 4.928729, 4.933709, 4.933207, 4.927653, 
    4.919489, 4.905965, 4.888046, 4.867195, 4.844253, 4.820849, 4.798853, 
    4.780519, 4.766601, 4.757459, 4.756906, 4.763144, 4.775598, 4.793231, 
    4.814648, 4.838199, 4.862067, 4.884343, 4.903111, 4.916597, 4.923395, 
    4.922756, 4.914888, 4.901155, 4.884047, 4.866805, 4.85282, 4.844973, 
    4.84515,
  // height(14,36, 0-49)
    4.991346, 4.964972, 4.940395, 4.918357, 4.899533, 4.884483, 4.873598, 
    4.867045, 4.864746, 4.866374, 4.871405, 4.879189, 4.889049, 4.900362, 
    4.912611, 4.910634, 4.912133, 4.919724, 4.921842, 4.919075, 4.911914, 
    4.903495, 4.890347, 4.873635, 4.854704, 4.834425, 4.814302, 4.79603, 
    4.781533, 4.77143, 4.765703, 4.768709, 4.777803, 4.792308, 4.811116, 
    4.832782, 4.855612, 4.877761, 4.897319, 4.912441, 4.921529, 4.923491, 
    4.918043, 4.905955, 4.889152, 4.870528, 4.853456, 4.841154, 4.836089, 
    4.839647,
  // height(14,37, 0-49)
    4.988453, 4.962273, 4.937971, 4.916267, 4.897817, 4.883152, 4.872628, 
    4.866377, 4.864271, 4.865924, 4.870734, 4.877946, 4.88674, 4.896296, 
    4.905811, 4.903345, 4.906444, 4.910737, 4.910229, 4.90555, 4.897175, 
    4.888714, 4.876239, 4.86105, 4.844311, 4.826896, 4.810146, 4.795563, 
    4.784745, 4.778251, 4.77579, 4.782004, 4.793592, 4.809768, 4.829356, 
    4.850853, 4.87252, 4.892492, 4.908888, 4.919978, 4.924416, 4.921508, 
    4.911499, 4.895743, 4.87667, 4.857455, 4.841446, 4.831538, 4.829711, 
    4.836845,
  // height(14,38, 0-49)
    4.984639, 4.958626, 4.934591, 4.913228, 4.895154, 4.880854, 4.870646, 
    4.86461, 4.862578, 4.864117, 4.868563, 4.875087, 4.882763, 4.890626, 
    4.897676, 4.89531, 4.900163, 4.901466, 4.898746, 4.892606, 4.88346, 
    4.875215, 4.863713, 4.850336, 4.836003, 4.821574, 4.808197, 4.797181, 
    4.789793, 4.786611, 4.787156, 4.796136, 4.809761, 4.82715, 4.84706, 
    4.867931, 4.887993, 4.905383, 4.918293, 4.92518, 4.925019, 4.917578, 
    4.903661, 4.885168, 4.864916, 4.846192, 4.832146, 4.825239, 4.826932, 
    4.837641,
  // height(14,39, 0-49)
    4.980752, 4.95491, 4.931138, 4.910096, 4.892348, 4.878327, 4.868291, 
    4.862281, 4.86009, 4.861258, 4.865097, 4.870739, 4.877207, 4.88346, 
    4.888396, 4.886341, 4.892785, 4.891613, 4.887215, 4.88012, 4.87067, 
    4.862928, 4.852697, 4.841382, 4.829606, 4.818201, 4.808114, 4.800452, 
    4.796173, 4.795929, 4.799117, 4.810341, 4.825474, 4.843554, 4.863278, 
    4.883053, 4.901103, 4.915614, 4.924913, 4.927712, 4.92337, 4.912158, 
    4.895406, 4.875451, 4.855321, 4.838219, 4.826949, 4.82348, 4.828774, 
    4.842854,
  // height(14,40, 0-49)
    4.977879, 4.952263, 4.928766, 4.908001, 4.890475, 4.876557, 4.866449, 
    4.860152, 4.857441, 4.857857, 4.860724, 4.86519, 4.87028, 4.874952, 
    4.878095, 4.876329, 4.883979, 4.880965, 4.875467, 4.867936, 4.858642, 
    4.851704, 4.843017, 4.833961, 4.824832, 4.816414, 4.809454, 4.804865, 
    4.80331, 4.805566, 4.810947, 4.823834, 4.839893, 4.8581, 4.87712, 
    4.895356, 4.911077, 4.92258, 4.928399, 4.927567, 4.919873, 4.906066, 
    4.88791, 4.868001, 4.849374, 4.834966, 4.827127, 4.827327, 4.836097, 
    4.853168,
  // height(14,41, 0-49)
    4.977243, 4.951975, 4.928784, 4.908237, 4.890777, 4.876709, 4.866188, 
    4.859186, 4.855484, 4.854657, 4.856086, 4.858981, 4.862435, 4.865462, 
    4.867022, 4.865379, 4.873715, 4.869505, 4.863459, 4.855964, 4.84724, 
    4.841386, 4.834473, 4.827814, 4.821355, 4.81582, 4.811758, 4.8099, 
    4.810643, 4.814913, 4.82198, 4.835919, 4.852301, 4.870073, 4.8879, 
    4.904237, 4.91746, 4.92605, 4.928823, 4.925181, 4.915336, 4.900439, 
    4.882529, 4.864255, 4.848449, 4.837637, 4.833674, 4.837571, 4.849523, 
    4.869064,
  // height(14,42, 0-49)
    4.980048, 4.955317, 4.932497, 4.912102, 4.894521, 4.880002, 4.868662, 
    4.860474, 4.855247, 4.852629, 4.852093, 4.852965, 4.854447, 4.855668, 
    4.855711, 4.853931, 4.862373, 4.857519, 4.851374, 4.844295, 4.836475, 
    4.831925, 4.826941, 4.822737, 4.818897, 4.816074, 4.814629, 4.815122, 
    4.817711, 4.823489, 4.831711, 4.846095, 4.862226, 4.879052, 4.895293, 
    4.909513, 4.92027, 4.926304, 4.926771, 4.921447, 4.910919, 4.896608, 
    4.88063, 4.865476, 4.85361, 4.847065, 4.847208, 4.854662, 4.869378, 
    4.89079,
  // height(14,43, 0-49)
    4.987293, 4.963366, 4.941016, 4.920723, 4.902826, 4.887541, 4.874972, 
    4.865113, 4.857836, 4.852889, 4.849873, 4.848258, 4.847405, 4.846586, 
    4.845038, 4.842797, 4.850761, 4.845643, 4.839696, 4.833277, 4.826568, 
    4.82345, 4.820451, 4.818665, 4.817314, 4.816969, 4.817812, 4.820253, 
    4.824242, 4.831039, 4.839899, 4.854184, 4.869569, 4.885051, 4.89946, 
    4.911537, 4.920093, 4.924184, 4.923324, 4.917646, 4.908003, 4.895916, 
    4.88339, 4.872587, 4.865491, 4.863626, 4.867915, 4.878666, 4.895671, 
    4.918324,
  // height(14,44, 0-49)
    4.999643, 4.97684, 4.955107, 4.934894, 4.916515, 4.900183, 4.886018, 
    4.874065, 4.864291, 4.85656, 4.850628, 4.846134, 4.842605, 4.839487, 
    4.83618, 4.833108, 4.840065, 4.83484, 4.82921, 4.823539, 4.818005, 
    4.81632, 4.815243, 4.815725, 4.816647, 4.818492, 4.821272, 4.825261, 
    4.830235, 4.837609, 4.846658, 4.8604, 4.874674, 4.888574, 4.901094, 
    4.911215, 4.918052, 4.921008, 4.91994, 4.915264, 4.907966, 4.899511, 
    4.891633, 4.886055, 4.884239, 4.887223, 4.895544, 4.909267, 4.928077, 
    4.951357,
  // height(14,45, 0-49)
    5.017312, 4.996, 4.97507, 4.95496, 4.935992, 4.918405, 4.902376, 4.88803, 
    4.875444, 4.864624, 4.855481, 4.847826, 4.841365, 4.835716, 4.83044, 
    4.826169, 4.831665, 4.826299, 4.820926, 4.815934, 4.811489, 4.81111, 
    4.811764, 4.814254, 4.81716, 4.820862, 4.825219, 4.830384, 4.835991, 
    4.843586, 4.852475, 4.865373, 4.878339, 4.890605, 4.901376, 4.909918, 
    4.915675, 4.918389, 4.918215, 4.915745, 4.911979, 4.908191, 4.905741, 
    4.90587, 4.909535, 4.917328, 4.92946, 4.945801, 4.965949, 4.989285,
  // height(14,46, 0-49)
    5.040022, 5.0206, 5.000702, 4.98078, 4.9612, 4.942265, 4.924236, 
    4.907354, 4.891817, 4.877773, 4.865296, 4.854357, 4.84483, 4.83649, 
    4.829052, 4.823248, 4.82694, 4.821243, 4.81594, 4.811431, 4.807864, 
    4.808546, 4.810627, 4.814773, 4.819308, 4.82451, 4.8301, 4.836121, 
    4.842098, 4.849669, 4.858179, 4.870093, 4.881728, 4.892483, 4.901812, 
    4.909278, 4.914648, 4.917972, 4.919623, 4.920277, 4.920839, 4.922309, 
    4.92564, 4.931595, 4.94067, 4.953065, 4.968709, 4.987298, 5.008345, 
    5.031216,
  // height(14,47, 0-49)
    5.067022, 5.049904, 5.031317, 5.011751, 4.991643, 4.971396, 4.951393, 
    4.931998, 4.913552, 4.896341, 4.880581, 4.866395, 4.853802, 4.842718, 
    4.832986, 4.825392, 4.827056, 4.820758, 4.815261, 4.810961, 4.807976, 
    4.809393, 4.812525, 4.817905, 4.823682, 4.830026, 4.836539, 4.843167, 
    4.849349, 4.856772, 4.86482, 4.875768, 4.8862, 4.89571, 4.904, 4.910928, 
    4.916553, 4.921173, 4.925306, 4.929629, 4.934891, 4.941786, 4.950864, 
    4.962459, 4.976653, 4.993308, 5.012097, 5.032546, 5.05407, 5.075994,
  // height(14,48, 0-49)
    5.097138, 5.082759, 5.065822, 5.046871, 5.026447, 5.005077, 4.983285, 
    4.961578, 4.940433, 4.920274, 4.901444, 4.884194, 4.868665, 4.854891, 
    4.842824, 4.833281, 4.832807, 4.825633, 4.819666, 4.81528, 4.812549, 
    4.814342, 4.818109, 4.824279, 4.830903, 4.838052, 4.845232, 4.852296, 
    4.858621, 4.86589, 4.873518, 4.883643, 4.893113, 4.901714, 4.90939, 
    4.916262, 4.922637, 4.928999, 4.935947, 4.944109, 4.954046, 4.966163, 
    4.980648, 4.997454, 5.016309, 5.036768, 5.058268, 5.080154, 5.101726, 
    5.122242,
  // height(14,49, 0-49)
    5.131782, 5.121768, 5.107812, 5.090503, 5.070491, 5.048445, 5.025044, 
    5.000954, 4.976798, 4.953141, 4.93047, 4.909184, 4.889575, 4.87183, 
    4.856054, 4.844022, 4.848143, 4.838534, 4.83033, 4.824347, 4.820787, 
    4.825149, 4.832235, 4.842608, 4.852149, 4.861037, 4.868387, 4.874065, 
    4.877024, 4.881012, 4.885324, 4.894529, 4.902976, 4.910685, 4.917894, 
    4.925021, 4.93263, 4.941376, 4.951897, 4.964715, 4.980152, 4.99826, 
    5.018826, 5.04138, 5.065258, 5.08966, 5.113735, 5.1366, 5.15739, 5.175267,
  // height(15,0, 0-49)
    5.116331, 5.087602, 5.057508, 5.02688, 4.99647, 4.966957, 4.938937, 
    4.912934, 4.889373, 4.86856, 4.850661, 4.835689, 4.823497, 4.813806, 
    4.806232, 4.800476, 4.797285, 4.793497, 4.79044, 4.787902, 4.785748, 
    4.784293, 4.783263, 4.78291, 4.783345, 4.784853, 4.787655, 4.791958, 
    4.797826, 4.805394, 4.814459, 4.825126, 4.83667, 4.848646, 4.860583, 
    4.872067, 4.882796, 4.892663, 4.901782, 4.910505, 4.919398, 4.929152, 
    4.940503, 4.954107, 4.970463, 4.989839, 5.012252, 5.037459, 5.064975, 
    5.094105,
  // height(15,1, 0-49)
    5.096625, 5.067094, 5.036662, 5.006133, 4.976219, 4.94755, 4.920673, 
    4.896048, 4.874031, 4.854852, 4.838602, 4.825209, 4.81445, 4.805967, 
    4.799304, 4.794245, 4.792803, 4.788857, 4.785463, 4.782435, 4.779634, 
    4.777761, 4.776192, 4.775315, 4.77516, 4.776093, 4.778361, 4.782217, 
    4.787709, 4.795141, 4.804237, 4.815469, 4.827672, 4.840302, 4.852779, 
    4.864544, 4.87516, 4.884389, 4.892262, 4.899111, 4.905552, 4.912408, 
    4.920602, 4.931015, 4.944372, 4.961137, 4.981477, 5.005255, 5.032047, 
    5.061183,
  // height(15,2, 0-49)
    5.078791, 5.048922, 5.018562, 4.988491, 4.95939, 4.931859, 4.906399, 
    4.883417, 4.863198, 4.845896, 4.831511, 4.819883, 4.810696, 4.803508, 
    4.797784, 4.793371, 4.793595, 4.789402, 4.78556, 4.781904, 4.778296, 
    4.775818, 4.773477, 4.771796, 4.770742, 4.770769, 4.772155, 4.775218, 
    4.780015, 4.787013, 4.795884, 4.807501, 4.820284, 4.833621, 4.846819, 
    4.859183, 4.870113, 4.879212, 4.886373, 4.891838, 4.89621, 4.900389, 
    4.905457, 4.912516, 4.922533, 4.936205, 4.953891, 4.975585, 5.000948, 
    5.029352,
  // height(15,3, 0-49)
    5.06324, 5.033447, 5.003518, 4.974208, 4.946181, 4.920012, 4.896168, 
    4.875008, 4.856752, 4.841472, 4.829074, 4.819304, 4.811752, 4.805884, 
    4.801088, 4.797221, 4.798965, 4.794469, 4.790111, 4.78574, 4.781212, 
    4.777983, 4.774674, 4.771935, 4.769695, 4.768483, 4.768632, 4.770534, 
    4.774281, 4.780493, 4.788819, 4.800562, 4.81377, 4.827785, 4.841828, 
    4.855076, 4.866765, 4.876311, 4.883421, 4.888182, 4.891104, 4.893085, 
    4.895307, 4.899062, 4.905564, 4.915772, 4.93028, 4.949261, 4.972499, 
    4.999438,
  // height(15,4, 0-49)
    5.050073, 5.020701, 4.9915, 4.963202, 4.936454, 4.911811, 4.889717, 
    4.87048, 4.854262, 4.841056, 4.830678, 4.822776, 4.81685, 4.812282, 
    4.808378, 4.804924, 4.807982, 4.803201, 4.798327, 4.79323, 4.787751, 
    4.783697, 4.779289, 4.77529, 4.771614, 4.768863, 4.767426, 4.767785, 
    4.770104, 4.775139, 4.782532, 4.794057, 4.807438, 4.822003, 4.836916, 
    4.851248, 4.864085, 4.874649, 4.88243, 4.887299, 4.88959, 4.890103, 
    4.890029, 4.890785, 4.89381, 4.900341, 4.911246, 4.92694, 4.947388, 
    4.972149,
  // height(15,5, 0-49)
    5.039103, 5.010417, 4.982175, 4.95508, 4.929761, 4.906757, 4.886483, 
    4.869208, 4.855032, 4.843874, 4.835467, 4.829376, 4.825019, 4.821709, 
    4.818674, 4.815492, 4.819603, 4.814657, 4.809369, 4.803624, 4.797256, 
    4.792387, 4.786834, 4.781446, 4.776152, 4.771607, 4.768267, 4.766716, 
    4.767217, 4.770647, 4.77667, 4.787555, 4.800759, 4.81563, 4.831312, 
    4.846801, 4.861059, 4.873127, 4.882268, 4.888099, 4.8907, 4.89067, 
    4.889099, 4.887434, 4.887277, 4.890124, 4.89716, 4.909099, 4.926156, 
    4.948071,
  // height(15,6, 0-49)
    5.029912, 5.00209, 4.974963, 4.949202, 4.925413, 4.904112, 4.885684, 
    4.870354, 4.85817, 4.848981, 4.84245, 4.838074, 4.835212, 4.833121, 
    4.830979, 4.827941, 4.832795, 4.827935, 4.822438, 4.816226, 4.809129, 
    4.803551, 4.796894, 4.790074, 4.783056, 4.776528, 4.771018, 4.767218, 
    4.765527, 4.766914, 4.771096, 4.780854, 4.793445, 4.80827, 4.824483, 
    4.841054, 4.856845, 4.870752, 4.88182, 4.889394, 4.893252, 4.893704, 
    4.891622, 4.888361, 4.885583, 4.885003, 4.888118, 4.895999, 4.909183, 
    4.927671,
  // height(15,7, 0-49)
    5.021935, 4.99507, 4.96914, 4.944782, 4.922575, 4.902999, 4.886406, 
    4.872977, 4.862704, 4.855379, 4.850611, 4.847847, 4.846417, 4.845552, 
    4.844402, 4.841412, 4.846661, 4.84226, 4.836864, 4.83046, 4.822882, 
    4.816778, 4.809143, 4.800937, 4.792175, 4.783555, 4.775673, 4.769339, 
    4.765112, 4.764037, 4.765896, 4.774005, 4.785484, 4.799817, 4.816212, 
    4.833632, 4.850895, 4.866778, 4.880141, 4.89007, 4.896023, 4.897958, 
    4.896429, 4.892569, 4.887981, 4.884502, 4.88391, 4.887653, 4.896658, 
    4.911267,
  // height(15,8, 0-49)
    5.014567, 4.988669, 4.963949, 4.941008, 4.920386, 4.902526, 4.887734, 
    4.876143, 4.867693, 4.862128, 4.859016, 4.857789, 4.857767, 4.858192, 
    4.858227, 4.855232, 4.860509, 4.857036, 4.852131, 4.845875, 4.838133, 
    4.83175, 4.82334, 4.813871, 4.803432, 4.792694, 4.782328, 4.773249, 
    4.766201, 4.762278, 4.76136, 4.767284, 4.777114, 4.790453, 4.806582, 
    4.824496, 4.842996, 4.860787, 4.876583, 4.889243, 4.897914, 4.902189, 
    4.902226, 4.898835, 4.893422, 4.887823, 4.884019, 4.883815, 4.888562, 
    4.899018,
  // height(15,9, 0-49)
    5.007263, 4.982272, 4.958714, 4.937149, 4.918076, 4.901892, 4.888849, 
    4.879029, 4.872319, 4.868426, 4.866897, 4.867163, 4.868573, 4.870416, 
    4.871912, 4.868925, 4.873866, 4.87183, 4.867853, 4.862131, 4.854586, 
    4.848204, 4.83927, 4.828737, 4.816766, 4.803984, 4.791113, 4.779171, 
    4.76909, 4.762001, 4.7579, 4.761126, 4.768773, 4.780583, 4.795938, 
    4.813896, 4.833264, 4.85271, 4.870847, 4.886352, 4.898101, 4.905329, 
    4.907785, 4.905872, 4.900687, 4.893928, 4.887661, 4.883976, 4.884649, 
    4.890883,
  // height(15,10, 0-49)
    4.999604, 4.975416, 4.952922, 4.932649, 4.915052, 4.900475, 4.889113, 
    4.880991, 4.875949, 4.873662, 4.873672, 4.875424, 4.878328, 4.881759, 
    4.885052, 4.882169, 4.886457, 4.886337, 4.883721, 4.878932, 4.87196, 
    4.865866, 4.856699, 4.845355, 4.832079, 4.817416, 4.802129, 4.787311, 
    4.774088, 4.7636, 4.755988, 4.756044, 4.760993, 4.770745, 4.784802, 
    4.802295, 4.822069, 4.84278, 4.862974, 4.881195, 4.896103, 4.906617, 
    4.912094, 4.912504, 4.908549, 4.901665, 4.893864, 4.887411, 4.884446, 
    4.886625,
  // height(15,11, 0-49)
    4.991342, 4.967822, 4.946262, 4.927166, 4.910937, 4.897869, 4.8881, 
    4.881597, 4.878156, 4.877424, 4.878942, 4.882198, 4.886673, 4.891865, 
    4.897288, 4.89474, 4.898158, 4.900331, 4.899464, 4.895978, 4.889944, 
    4.88441, 4.875308, 4.863452, 4.849164, 4.832879, 4.815373, 4.797784, 
    4.781417, 4.767402, 4.756055, 4.752538, 4.754327, 4.761522, 4.773763, 
    4.790272, 4.809944, 4.831436, 4.853266, 4.873887, 4.891792, 4.905651, 
    4.914472, 4.917807, 4.915928, 4.909914, 4.901585, 4.893248, 4.8873, 
    4.885808,
  // height(15,12, 0-49)
    4.982402, 4.959404, 4.938636, 4.920569, 4.905574, 4.893891, 4.885602, 
    4.880623, 4.878705, 4.879471, 4.882472, 4.887239, 4.893341, 4.900425, 
    4.908225, 4.906451, 4.908953, 4.913633, 4.914804, 4.91294, 4.908176, 
    4.903432, 4.894686, 4.88264, 4.867683, 4.850114, 4.830691, 4.810552, 
    4.791155, 4.773605, 4.758424, 4.751015, 4.749251, 4.753448, 4.763399, 
    4.778428, 4.797483, 4.819242, 4.842208, 4.86478, 4.885344, 4.90237, 
    4.914593, 4.92119, 4.922007, 4.917713, 4.90983, 4.900563, 4.892437, 
    4.887838,
  // height(15,13, 0-49)
    4.972854, 4.950241, 4.930109, 4.912913, 4.898992, 4.888544, 4.881598, 
    4.87802, 4.877524, 4.879713, 4.884143, 4.890391, 4.89812, 4.907125, 
    4.917382, 4.917123, 4.918903, 4.926107, 4.929477, 4.929471, 4.926257, 
    4.922477, 4.914348, 4.90243, 4.887171, 4.868714, 4.847758, 4.825398, 
    4.803198, 4.782228, 4.763248, 4.751732, 4.746114, 4.746946, 4.7542, 
    4.767303, 4.785262, 4.806781, 4.830365, 4.854382, 4.877144, 4.897, 
    4.912463, 4.922406, 4.926286, 4.924352, 4.917756, 4.908478, 4.899033, 
    4.892014,
  // height(15,14, 0-49)
    4.96287, 4.940514, 4.920871, 4.904384, 4.891365, 4.881975, 4.876204, 
    4.873875, 4.874665, 4.878159, 4.883919, 4.89156, 4.900823, 4.911641, 
    4.924194, 4.926576, 4.928138, 4.937673, 4.943261, 4.945259, 4.943804, 
    4.941094, 4.933791, 4.922291, 4.907089, 4.888156, 4.866101, 4.841918, 
    4.817236, 4.793077, 4.770475, 4.754752, 4.745088, 4.742292, 4.746523, 
    4.757329, 4.773777, 4.7946, 4.818307, 4.843254, 4.867715, 4.889956, 
    4.908341, 4.921505, 4.928574, 4.929399, 4.924733, 4.916243, 4.906309, 
    4.897605,
  // height(15,15, 0-49)
    4.952686, 4.930484, 4.911194, 4.895252, 4.88295, 4.874424, 4.869629, 
    4.868354, 4.870248, 4.874878, 4.881808, 4.890677, 4.901279, 4.913642, 
    4.92807, 4.93463, 4.936832, 4.948342, 4.95604, 4.960089, 4.960528, 
    4.958922, 4.952585, 4.941731, 4.926888, 4.907864, 4.885134, 4.85956, 
    4.832775, 4.80575, 4.779841, 4.759933, 4.746149, 4.739574, 4.740567, 
    4.748801, 4.763408, 4.783151, 4.806544, 4.831944, 4.857608, 4.881755, 
    4.90265, 4.918758, 4.928937, 4.932689, 4.930367, 4.923283, 4.913586, 
    4.903914,
  // height(15,16, 0-49)
    4.942564, 4.920435, 4.90138, 4.885822, 4.874048, 4.866168, 4.862118, 
    4.86166, 4.864422, 4.869958, 4.877826, 4.887679, 4.899335, 4.912846, 
    4.92854, 4.941131, 4.945195, 4.958213, 4.967833, 4.973904, 4.976303, 
    4.975766, 4.970457, 4.960384, 4.946107, 4.927279, 4.904236, 4.877665, 
    4.849168, 4.819665, 4.790876, 4.766929, 4.749082, 4.738706, 4.736363, 
    4.741861, 4.7544, 4.77277, 4.795497, 4.820938, 4.847348, 4.872924, 
    4.89588, 4.91456, 4.92762, 4.934264, 4.934485, 4.929224, 4.920336, 
    4.910336,
  // height(15,17, 0-49)
    4.932777, 4.910663, 4.891735, 4.876411, 4.864961, 4.857486, 4.853906, 
    4.853971, 4.857299, 4.863437, 4.871946, 4.88248, 4.894852, 4.909085, 
    4.925418, 4.945959, 4.953385, 4.967457, 4.978798, 4.986842, 4.991218, 
    4.991667, 4.987359, 4.978087, 4.964433, 4.945938, 4.922795, 4.895525, 
    4.865663, 4.834091, 4.80294, 4.77522, 4.753508, 4.739446, 4.733802, 
    4.736515, 4.746866, 4.76367, 4.785466, 4.810616, 4.837379, 4.863954, 
    4.888523, 4.909357, 4.924963, 4.934315, 4.937086, 4.933866, 4.926193, 
    4.916392,
  // height(15,18, 0-49)
    4.923589, 4.901454, 4.882562, 4.867312, 4.855964, 4.848607, 4.845161, 
    4.845378, 4.848886, 4.855247, 4.864042, 4.874938, 4.887739, 4.902402, 
    4.918972, 4.949069, 4.961415, 4.976269, 4.989225, 4.999232, 5.005604, 
    5.006928, 5.003522, 4.994929, 4.981759, 4.963496, 4.940249, 4.9124, 
    4.881422, 4.848179, 4.815248, 4.784146, 4.758912, 4.741425, 4.732646, 
    4.732654, 4.740804, 4.755947, 4.776639, 4.801248, 4.828047, 4.855239, 
    4.881002, 4.903563, 4.921335, 4.933104, 4.938289, 4.93716, 4.930946, 
    4.921741,
  // height(15,19, 0-49)
    4.915263, 4.893085, 4.874133, 4.858778, 4.847258, 4.839663, 4.83592, 
    4.835809, 4.838999, 4.845114, 4.853805, 4.864809, 4.877959, 4.89312, 
    4.910018, 4.950513, 4.968981, 4.984726, 4.999439, 5.011564, 5.02004, 
    5.022157, 5.019508, 5.011316, 4.998226, 4.979774, 4.956087, 4.927523, 
    4.895533, 4.860983, 4.826902, 4.792949, 4.764691, 4.744195, 4.732588, 
    4.730083, 4.736119, 4.749599, 4.769093, 4.792991, 4.819576, 4.847066, 
    4.873648, 4.897533, 4.917068, 4.93091, 4.938273, 4.939157, 4.934505, 
    4.926172,
  // height(15,20, 0-49)
    4.908185, 4.886056, 4.867468, 4.852916, 4.84274, 4.837077, 4.835821, 
    4.838592, 4.844738, 4.853366, 4.863411, 4.873747, 4.883327, 4.89133, 
    4.897302, 0, 4.994577, 4.999668, 5.005548, 5.011305, 5.016126, 5.015633, 
    5.013115, 5.006968, 4.997258, 4.982792, 4.962961, 4.937488, 4.907465, 
    4.873701, 4.839848, 4.803802, 4.772908, 4.749545, 4.735105, 4.72999, 
    4.733762, 4.745383, 4.763453, 4.786373, 4.812434, 4.839869, 4.866875, 
    4.891658, 4.912527, 4.928051, 4.937283, 4.939999, 4.936891, 4.929584,
  // height(15,21, 0-49)
    4.90235, 4.880386, 4.861916, 4.847402, 4.837146, 4.831253, 4.829581, 
    4.831733, 4.837054, 4.844685, 4.853627, 4.862837, 4.871323, 4.878238, 
    4.882979, 0, 5.004196, 5.009486, 5.015777, 5.021951, 5.027033, 5.024549, 
    5.020569, 5.013208, 5.002763, 4.988084, 4.968498, 4.943565, 4.914167, 
    4.880956, 4.847917, 4.810899, 4.778774, 4.753971, 4.737977, 4.73131, 
    4.733636, 4.743992, 4.761029, 4.783178, 4.80876, 4.836029, 4.863201, 
    4.888492, 4.910194, 4.926821, 4.937312, 4.941274, 4.939192, 4.932497,
  // height(15,22, 0-49)
    4.897773, 4.875886, 4.857458, 4.842922, 4.832562, 4.826463, 4.824469, 
    4.826171, 4.830924, 4.837883, 4.846084, 4.854511, 4.862186, 4.868207, 
    4.871812, 0, 5.010537, 5.015932, 5.022656, 5.029411, 5.035066, 5.0311, 
    5.026239, 5.01824, 5.007516, 4.992895, 4.973616, 4.949099, 4.920087, 
    4.887161, 4.854692, 4.816629, 4.78334, 4.757275, 4.739974, 4.732033, 
    4.73318, 4.742507, 4.758702, 4.78022, 4.805398, 4.83251, 4.859784, 
    4.885447, 4.907785, 4.925273, 4.936773, 4.941762, 4.940569, 4.934464,
  // height(15,23, 0-49)
    4.894632, 4.872791, 4.854372, 4.839801, 4.829348, 4.823086, 4.820855, 
    4.822244, 4.826617, 4.833141, 4.840868, 4.848798, 4.855937, 4.861334, 
    4.864092, 0, 5.014832, 5.020237, 5.02725, 5.034447, 5.040577, 5.035399, 
    5.029847, 5.021343, 5.010375, 4.995757, 4.976672, 4.952449, 4.923741, 
    4.891075, 4.859142, 4.82031, 4.786209, 4.75929, 4.741114, 4.732311, 
    4.73266, 4.741292, 4.75692, 4.778018, 4.802937, 4.829955, 4.857316, 
    4.883248, 4.906034, 4.924124, 4.93632, 4.94202, 4.941433, 4.935718,
  // height(15,24, 0-49)
    4.89303, 4.871227, 4.852822, 4.83823, 4.827715, 4.821345, 4.818963, 
    4.820161, 4.824309, 4.830588, 4.838061, 4.845731, 4.8526, 4.857682, 4.86, 
    0, 5.017446, 5.022851, 5.03004, 5.037525, 5.043984, 5.038036, 5.032043, 
    5.023195, 5.012022, 4.997339, 4.978312, 4.954233, 4.925709, 4.893244, 
    4.861749, 4.822506, 4.787988, 4.760626, 4.741983, 4.732702, 4.732585, 
    4.740788, 4.756044, 4.776845, 4.801548, 4.828448, 4.855792, 4.881816, 
    4.904807, 4.9232, 4.935774, 4.941876, 4.941653, 4.936192,
  // height(15,25, 0-49)
    4.892978, 4.871228, 4.852853, 4.838268, 4.827735, 4.821324, 4.818879, 
    4.820003, 4.824073, 4.830282, 4.8377, 4.84534, 4.852205, 4.857303, 
    4.859646, 0, 5.017977, 5.023447, 5.030755, 5.038391, 5.045011, 5.03886, 
    5.032743, 5.023767, 5.012475, 4.997696, 4.978612, 4.954521, 4.926036, 
    4.893661, 4.862384, 4.823091, 4.788538, 4.761134, 4.742421, 4.733041, 
    4.732802, 4.74087, 4.755989, 4.776659, 4.801252, 4.828063, 4.855346, 
    4.881342, 4.904335, 4.922764, 4.935397, 4.941571, 4.941417, 4.935998,
  // height(15,26, 0-49)
    4.894406, 4.87272, 4.854392, 4.839842, 4.829338, 4.822953, 4.820543, 
    4.82172, 4.82587, 4.832198, 4.839781, 4.84764, 4.854785, 4.860251, 
    4.863098, 0, 5.016332, 5.021949, 5.029336, 5.036996, 5.043603, 5.037862, 
    5.031976, 5.023129, 5.011848, 4.996982, 4.977752, 4.953513, 4.924929, 
    4.892527, 4.861219, 4.822248, 4.78804, 4.760976, 4.742573, 4.733451, 
    4.733408, 4.741605, 4.756795, 4.777483, 4.802044, 4.828778, 4.855942, 
    4.881776, 4.904565, 4.922753, 4.935126, 4.941044, 4.940664, 4.935086,
  // height(15,27, 0-49)
    4.89715, 4.875522, 4.857244, 4.842745, 4.83231, 4.826026, 4.823761, 
    4.825141, 4.829566, 4.836245, 4.84426, 4.852632, 4.860379, 4.866575, 
    4.870389, 0, 5.012642, 5.018445, 5.025831, 5.033369, 5.039788, 5.035005, 
    5.029674, 5.021203, 5.01006, 4.995123, 4.97568, 4.951184, 4.922391, 
    4.889878, 4.858337, 4.820057, 4.786572, 4.760231, 4.74251, 4.733994, 
    4.734449, 4.743031, 4.758483, 4.779317, 4.80391, 4.830564, 4.857533, 
    4.883053, 4.905414, 4.923075, 4.934859, 4.940183, 4.939286, 4.933345,
  // height(15,28, 0-49)
    4.900956, 4.87935, 4.861095, 4.846647, 4.83631, 4.830202, 4.828211, 
    4.829986, 4.834939, 4.842281, 4.851081, 4.860333, 4.869051, 4.876345, 
    4.881514, 0, 5.007342, 5.013274, 5.020514, 5.02774, 5.033801, 5.030379, 
    5.02587, 5.017995, 5.00712, 4.992149, 4.972463, 4.947652, 4.918607, 
    4.885978, 4.854132, 4.816909, 4.784528, 4.759285, 4.742601, 4.735004, 
    4.736219, 4.745374, 4.761208, 4.782232, 4.806831, 4.833304, 4.85991, 
    4.884882, 4.906523, 4.923325, 4.934174, 4.938588, 4.936932, 4.93051,
  // height(15,29, 0-49)
    4.905488, 4.883822, 4.865526, 4.851095, 4.840873, 4.835017, 4.833459, 
    4.83588, 4.841707, 4.850139, 4.860193, 4.870795, 4.8809, 4.889626, 
    4.896388, 0, 5.000063, 5.005975, 5.012874, 5.019604, 5.025175, 5.023331, 
    5.019852, 5.012797, 5.002379, 4.987502, 4.967638, 4.942543, 4.913272, 
    4.880569, 4.848407, 4.812506, 4.781537, 4.757733, 4.742431, 4.736076, 
    4.738331, 4.748291, 4.764679, 4.786003, 4.810646, 4.836909, 4.86304, 
    4.887277, 4.907935, 4.923557, 4.933121, 4.936285, 4.933587, 4.926498,
  // height(15,30, 0-49)
    4.910488, 4.888827, 4.870213, 4.855021, 4.843503, 4.83578, 4.831827, 
    4.831496, 4.834548, 4.840704, 4.849711, 4.861379, 4.875586, 4.892223, 
    4.911034, 4.954827, 4.973868, 4.991736, 5.008694, 5.022947, 5.033298, 
    5.035358, 5.033057, 5.025144, 5.012241, 4.993824, 4.97003, 4.941264, 
    4.909084, 4.874454, 4.840883, 4.805935, 4.77645, 4.754404, 4.74091, 
    4.73623, 4.739908, 4.750978, 4.768137, 4.789886, 4.814612, 4.84061, 
    4.866129, 4.889415, 4.908816, 4.922949, 4.930926, 4.932596, 4.928713, 
    4.920949,
  // height(15,31, 0-49)
    4.915942, 4.89447, 4.876083, 4.861194, 4.850078, 4.842865, 4.83952, 
    4.839871, 4.843635, 4.850474, 4.860056, 4.872119, 4.886497, 4.903143, 
    4.922074, 4.95497, 4.968733, 4.986028, 5.00144, 5.013679, 5.021948, 
    5.023351, 5.020294, 5.011942, 4.998954, 4.980783, 4.957542, 4.929637, 
    4.898599, 4.865321, 4.832775, 4.800514, 4.773793, 4.754419, 4.743352, 
    4.740744, 4.746068, 4.758324, 4.776205, 4.798216, 4.822738, 4.848071, 
    4.872464, 4.894181, 4.911629, 4.923537, 4.929198, 4.928702, 4.923073, 
    4.914211,
  // height(15,32, 0-49)
    4.921215, 4.899942, 4.881758, 4.8671, 4.856259, 4.849372, 4.846404, 
    4.847165, 4.851349, 4.858582, 4.868499, 4.880802, 4.895323, 4.912056, 
    4.93118, 4.954336, 4.96384, 4.98057, 4.994486, 5.004793, 5.011045, 
    5.011725, 5.007792, 4.99875, 4.985291, 4.966941, 4.943911, 4.916705, 
    4.886889, 4.855299, 4.824359, 4.795338, 4.771907, 4.755643, 4.747331, 
    4.746997, 4.754054, 4.767476, 4.785954, 4.808, 4.832004, 4.856267, 
    4.879059, 4.898688, 4.913652, 4.922843, 4.925797, 4.9229, 4.91548, 
    4.905674,
  // height(15,33, 0-49)
    4.92593, 4.904881, 4.886914, 4.872478, 4.861875, 4.855245, 4.852547, 
    4.853583, 4.858017, 4.865453, 4.875493, 4.887812, 4.902227, 4.91875, 
    4.937635, 4.952839, 4.959489, 4.975294, 4.98753, 4.995835, 5.000043, 
    4.999904, 4.99502, 4.985198, 4.971148, 4.952522, 4.929667, 4.903242, 
    4.874849, 4.845289, 4.816482, 4.7911, 4.771321, 4.758461, 4.753111, 
    4.755168, 4.763979, 4.778497, 4.797407, 4.819228, 4.842355, 4.865105, 
    4.885779, 4.902761, 4.914688, 4.920676, 4.920567, 4.915102, 4.905936, 
    4.895429,
  // height(15,34, 0-49)
    4.929762, 4.908973, 4.891263, 4.877086, 4.866748, 4.860384, 4.857946, 
    4.859209, 4.863815, 4.871333, 4.881327, 4.893431, 4.907422, 4.923276, 
    4.941233, 4.950496, 4.955647, 4.969988, 4.980257, 4.986433, 4.988561, 
    4.987503, 4.981656, 4.971096, 4.956528, 4.937751, 4.915259, 4.889861, 
    4.86318, 4.836005, 4.809812, 4.788346, 4.772446, 4.763155, 4.760866, 
    4.765345, 4.775867, 4.791358, 4.810493, 4.831789, 4.853648, 4.874407, 
    4.892422, 4.906191, 4.914549, 4.916904, 4.913468, 4.905375, 4.89462, 
    4.883753,
  // height(15,35, 0-49)
    4.932462, 4.911976, 4.894581, 4.880731, 4.870724, 4.864684, 4.862538, 
    4.864038, 4.868792, 4.87632, 4.886137, 4.897826, 4.911088, 4.925822, 
    4.942156, 4.947344, 4.952077, 4.964399, 4.972419, 4.976362, 4.976421, 
    4.974379, 4.967628, 4.95648, 4.941605, 4.922957, 4.901151, 4.877123, 
    4.852477, 4.828023, 4.80485, 4.787461, 4.77554, 4.769867, 4.77063, 
    4.777473, 4.789596, 4.805881, 4.824989, 4.845424, 4.865595, 4.883875, 
    4.898703, 4.908737, 4.913075, 4.911485, 4.904602, 4.893983, 4.881938, 
    4.87114,
  // height(15,36, 0-49)
    4.933903, 4.91376, 4.896746, 4.883297, 4.873699, 4.86805, 4.866251, 
    4.868015, 4.872907, 4.880397, 4.889943, 4.901053, 4.91335, 4.926611, 
    4.940794, 4.943399, 4.948446, 4.958294, 4.963863, 4.965548, 4.963623, 
    4.960588, 4.953065, 4.941565, 4.926686, 4.908533, 4.887803, 4.865521, 
    4.843225, 4.821772, 4.801928, 4.788659, 4.780696, 4.778567, 4.782275, 
    4.791337, 4.804873, 4.821717, 4.840497, 4.85971, 4.87777, 4.893103, 
    4.904272, 4.910153, 4.91017, 4.904511, 4.894277, 4.881431, 4.868542, 
    4.858325,
  // height(15,37, 0-49)
    4.934103, 4.914344, 4.897767, 4.884783, 4.875652, 4.870442, 4.86902, 
    4.871055, 4.876065, 4.883467, 4.892656, 4.903069, 4.914239, 4.925816, 
    4.937567, 4.938635, 4.944391, 4.951484, 4.954533, 4.954038, 4.950295, 
    4.946325, 4.938226, 4.926672, 4.912144, 4.894886, 4.875633, 4.855452, 
    4.83577, 4.817514, 4.801187, 4.791965, 4.787823, 4.789057, 4.795502, 
    4.806548, 4.821237, 4.838345, 4.856464, 4.874076, 4.889618, 4.9016, 
    4.908755, 4.910237, 4.905857, 4.896271, 4.883037, 4.868485, 4.855347, 
    4.846265,
  // height(15,38, 0-49)
    4.933275, 4.913924, 4.897812, 4.885321, 4.876671, 4.871897, 4.870824, 
    4.873085, 4.878146, 4.88538, 4.894122, 4.903744, 4.913695, 4.923514, 
    4.932799, 4.932977, 4.93955, 4.943816, 4.944435, 4.941947, 4.936632, 
    4.93186, 4.923436, 4.912159, 4.898354, 4.882379, 4.864967, 4.847182, 
    4.8303, 4.815341, 4.802587, 4.797229, 4.79666, 4.800972, 4.809848, 
    4.822561, 4.83807, 4.855095, 4.872189, 4.887829, 4.900504, 4.908844, 
    4.911808, 4.908888, 4.900332, 4.88727, 4.871682, 4.85616, 4.843473, 
    4.836088,
  // height(15,39, 0-49)
    4.931844, 4.912904, 4.897245, 4.885211, 4.876986, 4.87256, 4.871725, 
    4.874079, 4.879056, 4.885987, 4.894164, 4.902904, 4.911595, 4.919686, 
    4.926654, 4.926291, 4.933585, 4.935168, 4.933599, 4.929408, 4.922832, 
    4.91746, 4.909001, 4.898345, 4.885618, 4.871275, 4.856004, 4.840826, 
    4.826837, 4.815162, 4.805911, 4.804132, 4.80679, 4.813807, 4.824722, 
    4.838705, 4.85464, 4.871191, 4.88689, 4.900232, 4.909787, 4.914362, 
    4.913201, 4.906186, 4.894016, 4.878262, 4.861233, 4.845648, 4.834178, 
    4.828999,
  // height(15,40, 0-49)
    4.930457, 4.911899, 4.896629, 4.884946, 4.876993, 4.872725, 4.87191, 
    4.874125, 4.878788, 4.885204, 4.892647, 4.900396, 4.907799, 4.914251, 
    4.919162, 4.918425, 4.926207, 4.925446, 4.92205, 4.916519, 4.909047, 
    4.903338, 4.895158, 4.885455, 4.874131, 4.861706, 4.848792, 4.836337, 
    4.825235, 4.816731, 4.810798, 4.812224, 4.817683, 4.826947, 4.839435, 
    4.854232, 4.870153, 4.885829, 4.899788, 4.910583, 4.91692, 4.917839, 
    4.912915, 4.902449, 4.887573, 4.870214, 4.852869, 4.838229, 4.828725, 
    4.826172,
  // height(15,41, 0-49)
    4.929952, 4.911724, 4.896721, 4.885202, 4.877274, 4.872872, 4.871749, 
    4.873485, 4.877499, 4.883104, 4.889571, 4.896175, 4.902244, 4.907153, 
    4.910297, 4.909247, 4.917224, 4.914587, 4.909807, 4.903347, 4.895372, 
    4.889627, 4.882048, 4.873604, 4.863957, 4.853662, 4.843232, 4.833522, 
    4.825214, 4.819678, 4.816773, 4.820962, 4.828731, 4.839725, 4.853273, 
    4.868386, 4.883842, 4.898261, 4.910213, 4.918354, 4.921581, 4.919222, 
    4.911222, 4.898285, 4.881907, 4.864242, 4.847815, 4.835123, 4.828254, 
    4.828617,
  // height(15,42, 0-49)
    4.931294, 4.913325, 4.898424, 4.886817, 4.878589, 4.873669, 4.871818, 
    4.872636, 4.875574, 4.879983, 4.885159, 4.890398, 4.895037, 4.898464, 
    4.900094, 4.898733, 4.906603, 4.902615, 4.896917, 4.88995, 4.881868, 
    4.876405, 4.86973, 4.862811, 4.855051, 4.847018, 4.839118, 4.832088, 
    4.826405, 4.823557, 4.823317, 4.829775, 4.83932, 4.851501, 4.865571, 
    4.880503, 4.89507, 4.907923, 4.917725, 4.923294, 4.923772, 4.918811, 
    4.908726, 4.894571, 4.878089, 4.861507, 4.847205, 4.837363, 4.833653, 
    4.837076,
  // height(15,43, 0-49)
    4.935475, 4.917697, 4.902711, 4.890727, 4.881828, 4.875952, 4.872892, 
    4.872292, 4.873665, 4.876423, 4.879921, 4.883506, 4.886554, 4.888489, 
    4.888772, 4.887052, 4.894532, 4.889695, 4.883519, 4.876438, 4.868618, 
    4.863738, 4.85823, 4.853035, 4.847303, 4.841592, 4.836183, 4.831695, 
    4.828406, 4.827918, 4.829926, 4.83814, 4.84892, 4.86174, 4.875812, 
    4.89011, 4.90344, 4.914546, 4.922236, 4.925542, 4.923896, 4.917282, 
    4.906342, 4.892384, 4.877251, 4.863077, 4.851962, 4.845681, 4.845468, 
    4.851949,
  // height(15,44, 0-49)
    4.943389, 4.925753, 4.910508, 4.897867, 4.887924, 4.880651, 4.875891, 
    4.873359, 4.872651, 4.87327, 4.874662, 4.876251, 4.877479, 4.87783, 
    4.876827, 4.87465, 4.881481, 4.876204, 4.869909, 4.863044, 4.855793, 
    4.851745, 4.847598, 4.844251, 4.840609, 4.837198, 4.834173, 4.832032, 
    4.830871, 4.832383, 4.836201, 4.845671, 4.857166, 4.870117, 4.883736, 
    4.897036, 4.908914, 4.918256, 4.924076, 4.925666, 4.922758, 4.91564, 
    4.905199, 4.892863, 4.880429, 4.869793, 4.862683, 4.860432, 4.863861, 
    4.873267,
  // height(15,45, 0-49)
    4.955724, 4.938224, 4.922591, 4.909056, 4.897744, 4.88868, 4.881776, 
    4.876834, 4.873561, 4.871572, 4.870428, 4.86966, 4.868797, 4.867399, 
    4.865062, 4.862271, 4.868221, 4.862769, 4.856599, 4.850181, 4.843715, 
    4.840663, 4.837982, 4.836504, 4.834927, 4.833717, 4.832911, 4.832884, 
    4.833569, 4.836724, 4.841933, 4.852195, 4.863946, 4.876606, 4.889421, 
    4.901495, 4.911865, 4.919618, 4.924015, 4.924632, 4.921483, 4.915091, 
    4.906478, 4.897058, 4.888436, 4.882178, 4.879595, 4.881592, 4.888622, 
    4.900716,
  // height(15,46, 0-49)
    4.972857, 4.955551, 4.939471, 4.924886, 4.911969, 4.900812, 4.891409, 
    4.883674, 4.877432, 4.872438, 4.868383, 4.864922, 4.861692, 4.858339, 
    4.854538, 4.850924, 4.855777, 4.850251, 4.844319, 4.838459, 4.832879, 
    4.830882, 4.82966, 4.82997, 4.830338, 4.831164, 4.832362, 4.834197, 
    4.836456, 4.840928, 4.847151, 4.857822, 4.869471, 4.881536, 4.893338, 
    4.904113, 4.913095, 4.919608, 4.923187, 4.923685, 4.921351, 4.916856, 
    4.911235, 4.905757, 4.901744, 4.900376, 4.902549, 4.908782, 4.91922, 
    4.933684,
  // height(15,47, 0-49)
    4.994822, 4.977833, 4.961337, 4.945648, 4.931002, 4.917567, 4.905441, 
    4.894656, 4.885172, 4.87689, 4.869647, 4.863233, 4.857401, 4.851891, 
    4.846448, 4.841775, 4.845335, 4.839686, 4.833971, 4.828657, 4.82394, 
    4.822939, 4.823054, 4.824963, 4.827073, 4.829704, 4.832666, 4.836111, 
    4.839708, 4.845225, 4.85217, 4.862968, 4.874279, 4.885587, 4.896322, 
    4.905891, 4.913754, 4.9195, 4.922939, 4.92417, 4.923613, 4.921988, 
    4.920238, 4.919398, 4.920445, 4.924166, 4.931067, 4.941337, 4.954875, 
    4.971336,
  // height(15,48, 0-49)
    5.021287, 5.004817, 4.988027, 4.971284, 4.954903, 4.939142, 4.92421, 
    4.910266, 4.897417, 4.885714, 4.875143, 4.865629, 4.857044, 4.849217, 
    4.841962, 4.835991, 4.838085, 4.832155, 4.826528, 4.821638, 4.817649, 
    4.817477, 4.818703, 4.821928, 4.825503, 4.829668, 4.834137, 4.838961, 
    4.843709, 4.850078, 4.857544, 4.868315, 4.879192, 4.88973, 4.899494, 
    4.908081, 4.915195, 4.920693, 4.92464, 4.927336, 4.929301, 4.931226, 
    4.933884, 4.938024, 4.944261, 4.953, 4.964405, 4.978386, 4.994637, 5.01268,
  // height(15,49, 0-49)
    5.058356, 5.043217, 5.026606, 5.00895, 4.990648, 4.972076, 4.953585, 
    4.935503, 4.918123, 4.901687, 4.886375, 4.872292, 4.859453, 4.847805, 
    4.837231, 4.829314, 4.83676, 4.82897, 4.82178, 4.815975, 4.811789, 
    4.814678, 4.819662, 4.827548, 4.834721, 4.8415, 4.847211, 4.851875, 
    4.854626, 4.859023, 4.86429, 4.875, 4.885332, 4.89494, 4.903584, 
    4.911133, 4.917612, 4.923219, 4.928326, 4.933444, 4.939155, 4.946041, 
    4.9546, 4.965176, 4.977912, 4.992743, 5.009426, 5.027546, 5.046576, 
    5.065892,
  // height(16,0, 0-49)
    5.010379, 4.983305, 4.957535, 4.933589, 4.911873, 4.89267, 4.876139, 
    4.862313, 4.851107, 4.842322, 4.835676, 4.830809, 4.827321, 4.824801, 
    4.82285, 4.821224, 4.82087, 4.8188, 4.816489, 4.813863, 4.810887, 
    4.80795, 4.804797, 4.801712, 4.798837, 4.796524, 4.795112, 4.794984, 
    4.796442, 4.799865, 4.805302, 4.813079, 4.822648, 4.833603, 4.845372, 
    4.857257, 4.868512, 4.878438, 4.88649, 4.892384, 4.896164, 4.898243, 
    4.899375, 4.90057, 4.90296, 4.907646, 4.915551, 4.92732, 4.943265, 
    4.963357,
  // height(16,1, 0-49)
    4.998121, 4.971027, 4.945522, 4.922115, 4.901196, 4.88303, 4.86775, 
    4.855347, 4.845687, 4.838506, 4.833449, 4.830081, 4.827929, 4.826505, 
    4.825345, 4.824247, 4.825438, 4.823134, 4.820419, 4.817234, 4.813533, 
    4.810053, 4.806176, 4.802295, 4.798471, 4.795121, 4.792607, 4.79137, 
    4.791726, 4.794225, 4.798886, 4.806432, 4.81596, 4.827044, 4.839068, 
    4.851271, 4.86282, 4.87292, 4.880921, 4.886435, 4.889426, 4.890259, 
    4.889693, 4.888795, 4.888814, 4.891007, 4.896475, 4.906033, 4.920139, 
    4.938877,
  // height(16,2, 0-49)
    4.988944, 4.96211, 4.937086, 4.914367, 4.894336, 4.877245, 4.863204, 
    4.852176, 4.84398, 4.838302, 4.834718, 4.832727, 4.831792, 4.831364, 
    4.830914, 4.830249, 4.832897, 4.830378, 4.827298, 4.8236, 4.819216, 
    4.815224, 4.810616, 4.805884, 4.801012, 4.796468, 4.792636, 4.790017, 
    4.788951, 4.790158, 4.793639, 4.800545, 4.809657, 4.82056, 4.832631, 
    4.845079, 4.857021, 4.867584, 4.876018, 4.881814, 4.884809, 4.885249, 
    4.883801, 4.88151, 4.879666, 4.879637, 4.882692, 4.889841, 4.901728, 
    4.918592,
  // height(16,3, 0-49)
    4.98254, 4.95621, 4.931844, 4.90993, 4.890845, 4.874831, 4.861982, 
    4.852237, 4.845376, 4.841043, 4.838762, 4.837986, 4.838121, 4.838571, 
    4.838752, 4.838411, 4.842396, 4.83975, 4.836403, 4.832302, 4.827349, 
    4.822939, 4.817657, 4.812073, 4.806106, 4.800255, 4.794926, 4.790676, 
    4.787887, 4.787426, 4.789301, 4.795124, 4.80339, 4.813739, 4.82558, 
    4.838131, 4.850492, 4.86174, 4.871041, 4.877756, 4.88156, 4.882516, 
    4.881122, 4.878296, 4.87528, 4.873495, 4.874341, 4.879025, 4.888411, 
    4.902944,
  // height(16,4, 0-49)
    4.978348, 4.952726, 4.929165, 4.908149, 4.890049, 4.875096, 4.863371, 
    4.854793, 4.849114, 4.845946, 4.844783, 4.845037, 4.846092, 4.847313, 
    4.848078, 4.847959, 4.853121, 4.85051, 4.847063, 4.842731, 4.837382, 
    4.832712, 4.826875, 4.8205, 4.813451, 4.806242, 4.799288, 4.793202, 
    4.788418, 4.785934, 4.785778, 4.790048, 4.797011, 4.806389, 4.817661, 
    4.830092, 4.842803, 4.854854, 4.865345, 4.873514, 4.878854, 4.881207, 
    4.880831, 4.878424, 4.875085, 4.872192, 4.871225, 4.873564, 4.880309, 
    4.89215,
  // height(16,5, 0-49)
    4.975636, 4.950883, 4.928251, 4.908212, 4.891126, 4.877218, 4.866553, 
    4.859032, 4.85439, 4.852214, 4.851986, 4.853107, 4.85495, 4.856871, 
    4.858217, 4.858232, 4.864367, 4.862026, 4.858702, 4.854363, 4.848849, 
    4.844121, 4.837903, 4.830859, 4.822809, 4.814256, 4.805618, 4.797554, 
    4.790562, 4.785738, 4.78315, 4.785407, 4.790595, 4.798553, 4.808867, 
    4.820886, 4.833784, 4.84663, 4.858483, 4.868478, 4.87593, 4.880437, 
    4.881971, 4.880943, 4.878209, 4.875005, 4.872805, 4.87311, 4.877246, 
    4.886169,
  // height(16,6, 0-49)
    4.97359, 4.949832, 4.92823, 4.909238, 4.893208, 4.880342, 4.870695, 
    4.864148, 4.860424, 4.859102, 4.859666, 4.861528, 4.864074, 4.866668, 
    4.868656, 4.868736, 4.875587, 4.873809, 4.870874, 4.866787, 4.861371, 
    4.856816, 4.85043, 4.842885, 4.83398, 4.824172, 4.81387, 4.803766, 
    4.794423, 4.787009, 4.781643, 4.781456, 4.784411, 4.790498, 4.799439, 
    4.810699, 4.823528, 4.837036, 4.850263, 4.862264, 4.872192, 4.87941, 
    4.883584, 4.884794, 4.883579, 4.880935, 4.878224, 4.876989, 4.878732, 
    4.884682,
  // height(16,7, 0-49)
    4.971429, 4.948754, 4.928265, 4.910394, 4.895467, 4.883669, 4.87503, 
    4.869415, 4.866539, 4.865985, 4.867253, 4.869784, 4.872997, 4.876294, 
    4.879041, 4.879138, 4.8864, 4.885508, 4.883248, 4.879677, 4.874628, 
    4.870487, 4.864169, 4.856335, 4.846771, 4.835867, 4.824009, 4.811897, 
    4.800161, 4.789993, 4.781582, 4.778574, 4.778876, 4.782658, 4.789808, 
    4.799926, 4.812365, 4.826291, 4.840752, 4.85474, 4.86728, 4.877518, 
    4.884831, 4.888952, 4.890053, 4.888813, 4.886382, 4.88424, 4.883992, 
    4.887099,
  // height(16,8, 0-49)
    4.9685, 4.946961, 4.927648, 4.910966, 4.897206, 4.886523, 4.878919, 
    4.874241, 4.872197, 4.872381, 4.874321, 4.877502, 4.881399, 4.885472, 
    4.889145, 4.889234, 4.896564, 4.896873, 4.895561, 4.892765, 4.888341, 
    4.884839, 4.878826, 4.870933, 4.860958, 4.849187, 4.835968, 4.82198, 
    4.807916, 4.794942, 4.783319, 4.777194, 4.774482, 4.775564, 4.780519, 
    4.789104, 4.800787, 4.814806, 4.83023, 4.846014, 4.861082, 4.874398, 
    4.885083, 4.892534, 4.896551, 4.897444, 4.896061, 4.893718, 4.892021, 
    4.892599,
  // height(16,9, 0-49)
    4.964339, 4.943954, 4.92586, 4.910425, 4.897897, 4.888393, 4.88188, 
    4.878181, 4.876997, 4.87794, 4.88057, 4.88443, 4.889064, 4.894015, 
    4.898808, 4.898908, 4.90595, 4.907724, 4.907599, 4.905803, 4.90224, 
    4.89956, 4.894073, 4.886361, 4.876246, 4.863895, 4.849592, 4.833972, 
    4.817759, 4.802047, 4.787168, 4.777723, 4.771718, 4.769764, 4.772158, 
    4.778826, 4.789371, 4.803106, 4.81913, 4.836383, 4.853708, 4.869932, 
    4.883956, 4.894887, 4.902172, 4.905732, 4.906059, 4.904214, 4.901698, 
    4.900219,
  // height(16,10, 0-49)
    4.958708, 4.939458, 4.922597, 4.908445, 4.897206, 4.888947, 4.88359, 
    4.880938, 4.880676, 4.882433, 4.885808, 4.890401, 4.895841, 4.901774, 
    4.907865, 4.908079, 4.914513, 4.917924, 4.919169, 4.918551, 4.916037, 
    4.914315, 4.909543, 4.902239, 4.892272, 4.879665, 4.864626, 4.847709, 
    4.829641, 4.811388, 4.793344, 4.780487, 4.770998, 4.76575, 4.765265, 
    4.769666, 4.77869, 4.791737, 4.807944, 4.826241, 4.845419, 4.864198, 
    4.881311, 4.895623, 4.906263, 4.912791, 4.915321, 4.914591, 4.911907, 
    4.908954,
  // height(16,11, 0-49)
    4.951579, 4.933411, 4.917763, 4.904904, 4.894985, 4.88802, 4.883884, 
    4.882345, 4.883079, 4.88572, 4.889904, 4.895293, 4.901602, 4.9086, 
    4.916114, 4.916668, 4.922263, 4.927371, 4.930091, 4.930777, 4.929453, 
    4.928766, 4.924852, 4.918157, 4.908612, 4.89609, 4.88071, 4.862903, 
    4.84337, 4.822893, 4.801913, 4.785665, 4.77261, 4.763888, 4.760275, 
    4.762101, 4.769247, 4.781209, 4.797158, 4.816027, 4.836568, 4.857426, 
    4.877209, 4.894594, 4.908454, 4.918019, 4.923042, 4.923909, 4.92166, 
    4.917865,
  // height(16,12, 0-49)
    4.94311, 4.925941, 4.911447, 4.899851, 4.89125, 4.885598, 4.882725, 
    4.882352, 4.884141, 4.887729, 4.892781, 4.899015, 4.906228, 4.914317, 
    4.923285, 4.924597, 4.929274, 4.936002, 4.940219, 4.942276, 4.942241, 
    4.942596, 4.939634, 4.933708, 4.924829, 4.912722, 4.897404, 4.879156, 
    4.858614, 4.836325, 4.812768, 4.793261, 4.776662, 4.764382, 4.757468, 
    4.756468, 4.761423, 4.771923, 4.787184, 4.80614, 4.827521, 4.849919, 
    4.871853, 4.891866, 4.908628, 4.921103, 4.928713, 4.931497, 4.930191, 
    4.926173,
  // height(16,13, 0-49)
    4.933587, 4.917305, 4.903876, 4.893475, 4.886146, 4.881787, 4.880175, 
    4.88099, 4.883869, 4.888443, 4.894396, 4.901491, 4.909599, 4.918728, 
    4.929043, 4.931781, 4.935657, 4.943816, 4.94947, 4.952912, 4.954217, 
    4.955572, 4.953596, 4.948547, 4.940525, 4.92912, 4.914241, 4.895998, 
    4.874925, 4.8513, 4.825628, 4.803096, 4.783074, 4.767251, 4.756944, 
    4.752938, 4.755445, 4.764153, 4.778327, 4.796912, 4.81862, 4.842006, 
    4.865535, 4.887653, 4.906889, 4.921998, 4.932122, 4.936985, 4.937004, 
    4.933322,
  // height(16,14, 0-49)
    4.923371, 4.90785, 4.895366, 4.886055, 4.879909, 4.876776, 4.87638, 
    4.87836, 4.882319, 4.887879, 4.894729, 4.902659, 4.9116, 4.921633, 
    4.933037, 4.938135, 4.941565, 4.95087, 4.957839, 4.962636, 4.965298, 
    4.967563, 4.966561, 4.962437, 4.955395, 4.944908, 4.93078, 4.912937, 
    4.891786, 4.867318, 4.84006, 4.814806, 4.791577, 4.772316, 4.758617, 
    4.751506, 4.751376, 4.758027, 4.770776, 4.788579, 4.810141, 4.833998, 
    4.858574, 4.882263, 4.903494, 4.920869, 4.933316, 4.940278, 4.941876, 
    4.938986,
  // height(16,15, 0-49)
    4.912854, 4.897959, 4.88628, 4.877921, 4.87283, 4.870809, 4.871537, 
    4.874606, 4.87959, 4.886088, 4.893784, 4.90248, 4.912133, 4.922858, 
    4.93496, 4.94358, 4.947157, 4.957278, 4.965407, 4.971506, 4.97552, 
    4.978578, 4.978491, 4.975286, 4.969269, 4.959824, 4.946657, 4.929514, 
    4.908661, 4.883808, 4.855515, 4.827887, 4.801735, 4.779232, 4.762231, 
    4.752002, 4.749129, 4.753531, 4.764589, 4.781275, 4.80229, 4.826159, 
    4.851291, 4.876046, 4.898795, 4.918036, 4.932535, 4.941511, 4.944815, 
    4.943059,
  // height(16,16, 0-49)
    4.902413, 4.888007, 4.876982, 4.869414, 4.865215, 4.864151, 4.865855, 
    4.869885, 4.87578, 4.883116, 4.891562, 4.900916, 4.911123, 4.922285, 
    4.934649, 4.948032, 4.952551, 4.96318, 4.972324, 4.979673, 4.985033, 
    4.98876, 4.989505, 4.98716, 4.982129, 4.973736, 4.961613, 4.945337, 
    4.92504, 4.900175, 4.871372, 4.841729, 4.81299, 4.787511, 4.767387, 
    4.75412, 4.748487, 4.750541, 4.759723, 4.775039, 4.795194, 4.818704, 
    4.843974, 4.86935, 4.893178, 4.913892, 4.930142, 4.940972, 4.946005, 
    4.945608,
  // height(16,17, 0-49)
    4.892386, 4.878341, 4.867813, 4.860855, 4.857354, 4.857041, 4.859523, 
    4.864323, 4.870955, 4.878976, 4.88804, 4.897923, 4.908541, 4.919922, 
    4.932185, 4.951418, 4.957764, 4.968699, 4.978784, 4.987378, 4.994099, 
    4.998383, 4.999869, 4.998282, 4.994113, 4.986661, 4.975505, 4.960099, 
    4.940459, 4.915834, 4.886974, 4.855661, 4.824695, 4.796576, 4.773589, 
    4.757456, 4.749144, 4.748833, 4.756054, 4.769843, 4.78891, 4.811782, 
    4.836864, 4.862501, 4.88703, 4.908854, 4.926551, 4.939031, 4.945736, 
    4.946805,
  // height(16,18, 0-49)
    4.883057, 4.86925, 4.859056, 4.852509, 4.849472, 4.849656, 4.852646, 
    4.857956, 4.865088, 4.873597, 4.88313, 4.893447, 4.904416, 4.91596, 
    4.927983, 4.95368, 4.962641, 4.973895, 4.984979, 4.994907, 5.003065, 
    5.007842, 5.009997, 5.009035, 5.005515, 4.998745, 4.988299, 4.973565, 
    4.954499, 4.930216, 4.901648, 4.868981, 4.836173, 4.805798, 4.780288, 
    4.761552, 4.750729, 4.748141, 4.753402, 4.76559, 4.783442, 4.805486, 
    4.83014, 4.855759, 4.880685, 4.903311, 4.922166, 4.936076, 4.944336, 
    4.946891,
  // height(16,19, 0-49)
    4.874649, 4.860956, 4.850918, 4.844546, 4.841686, 4.842038, 4.845186, 
    4.850657, 4.857982, 4.866745, 4.876626, 4.887396, 4.898871, 4.910821, 
    4.922827, 4.954803, 4.966801, 4.978681, 4.991045, 5.002561, 5.012359, 
    5.017647, 5.020454, 5.019977, 5.016799, 5.010279, 5.000051, 4.985547, 
    4.966752, 4.942739, 4.9147, 4.880971, 4.846727, 4.814543, 4.786932, 
    4.765944, 4.752872, 4.748176, 4.751559, 4.76216, 4.778742, 4.799853, 
    4.823924, 4.849325, 4.874414, 4.897583, 4.917346, 4.932465, 4.942127, 
    4.946119,
  // height(16,20, 0-49)
    4.867816, 4.854584, 4.845321, 4.840126, 4.838893, 4.841312, 4.846864, 
    4.85486, 4.864492, 4.874896, 4.885221, 4.894706, 4.902756, 4.909014, 
    4.913389, 0, 4.987489, 4.991956, 4.99765, 5.003873, 5.010102, 5.012218, 
    5.01397, 5.014071, 5.012827, 5.009157, 5.002196, 4.990902, 4.974914, 
    4.953116, 4.927007, 4.893116, 4.858006, 4.824359, 4.79484, 4.771689, 
    4.756392, 4.749557, 4.751001, 4.759923, 4.775121, 4.79516, 4.818483, 
    4.843477, 4.868512, 4.891992, 4.912422, 4.928527, 4.93941, 4.944731,
  // height(16,21, 0-49)
    4.861976, 4.848943, 4.839874, 4.834837, 4.833697, 4.836112, 4.841539, 
    4.849289, 4.858567, 4.868547, 4.878441, 4.887538, 4.895265, 4.901219, 
    4.905196, 0, 4.992397, 4.997305, 5.003582, 5.010384, 5.017054, 5.017688, 
    5.018337, 5.017498, 5.015707, 5.011953, 5.005382, 4.994881, 4.979984, 
    4.959462, 4.935041, 4.90137, 4.866254, 4.832252, 4.801982, 4.777731, 
    4.761089, 4.752796, 4.752783, 4.760341, 4.774326, 4.793342, 4.815856, 
    4.840277, 4.864996, 4.888429, 4.909086, 4.925674, 4.937243, 4.943362,
  // height(16,22, 0-49)
    4.857375, 4.844437, 4.83546, 4.830493, 4.82939, 4.83179, 4.837147, 
    4.844765, 4.853857, 4.863614, 4.873266, 4.882125, 4.889603, 4.895244, 
    4.898731, 0, 4.995681, 5.000916, 5.007755, 5.015225, 5.022527, 5.022017, 
    5.021948, 5.020552, 5.018504, 5.014805, 5.008574, 4.99863, 4.984444, 
    4.964725, 4.941484, 4.907679, 4.872356, 4.837974, 4.807092, 4.781999, 
    4.764341, 4.754937, 4.753801, 4.760295, 4.773324, 4.791523, 4.813382, 
    4.837328, 4.86177, 4.885137, 4.905946, 4.922899, 4.935011, 4.941789,
  // height(16,23, 0-49)
    4.854089, 4.841188, 4.83224, 4.82729, 4.82618, 4.828554, 4.833859, 
    4.841405, 4.850407, 4.860065, 4.869614, 4.878358, 4.885695, 4.891115, 
    4.894202, 0, 4.998227, 5.003655, 5.010888, 5.018858, 5.026659, 5.025187, 
    5.024527, 5.02266, 5.020362, 5.016635, 5.010581, 5.000975, 4.98724, 
    4.968055, 4.945672, 4.911668, 4.876164, 4.841541, 4.810292, 4.784687, 
    4.76639, 4.756265, 4.754383, 4.760154, 4.772521, 4.790148, 4.811541, 
    4.835138, 4.85936, 4.882646, 4.903519, 4.920674, 4.933112, 4.940302,
  // height(16,24, 0-49)
    4.852131, 4.839238, 4.830288, 4.825319, 4.824179, 4.826513, 4.831777, 
    4.839285, 4.848259, 4.8579, 4.867444, 4.876188, 4.88351, 4.888863, 
    4.891764, 0, 5.000336, 5.005877, 5.013352, 5.021645, 5.029784, 5.027698, 
    5.026659, 5.024476, 5.021976, 5.018165, 5.01214, 5.002656, 4.989122, 
    4.970199, 4.948319, 4.914134, 4.878489, 4.843718, 4.812261, 4.786366, 
    4.767694, 4.757131, 4.754774, 4.760069, 4.771986, 4.789208, 4.810258, 
    4.833585, 4.857615, 4.880801, 4.901666, 4.918907, 4.931514, 4.938937,
  // height(16,25, 0-49)
    4.85146, 4.838564, 4.829591, 4.824589, 4.823408, 4.825703, 4.830941, 
    4.838443, 4.847441, 4.857141, 4.866776, 4.875635, 4.883084, 4.888557, 
    4.891555, 0, 5.001617, 5.00724, 5.014842, 5.023288, 5.03158, 5.02933, 
    5.02819, 5.025898, 5.02329, 5.019381, 5.01327, 5.003716, 4.990139, 
    4.971201, 4.949409, 4.915092, 4.87936, 4.844524, 4.813005, 4.787022, 
    4.768224, 4.757499, 4.754951, 4.760036, 4.771738, 4.788752, 4.809611, 
    4.83277, 4.856662, 4.879742, 4.900535, 4.917737, 4.930336, 4.937777,
  // height(16,26, 0-49)
    4.851977, 4.839075, 4.830077, 4.825035, 4.82382, 4.826095, 4.831341, 
    4.838893, 4.847992, 4.857843, 4.867679, 4.876782, 4.884514, 4.890315, 
    4.893711, 0, 5.001983, 5.007671, 5.015292, 5.023718, 5.031972, 5.030043, 
    5.029104, 5.026941, 5.024355, 5.020361, 5.014077, 5.004286, 4.990434, 
    4.971213, 4.949087, 4.914718, 4.878968, 4.844158, 4.812709, 4.786823, 
    4.768129, 4.757494, 4.755009, 4.760123, 4.771822, 4.788801, 4.809599, 
    4.832676, 4.856466, 4.87942, 4.900066, 4.917099, 4.929512, 4.936756,
  // height(16,27, 0-49)
    4.853549, 4.84063, 4.831599, 4.826528, 4.825302, 4.827601, 4.832926, 
    4.840624, 4.849943, 4.860089, 4.870278, 4.879788, 4.887972, 4.894296, 
    4.898354, 0, 5.001553, 5.007257, 5.014753, 5.022965, 5.030978, 5.02979, 
    5.029314, 5.027491, 5.025039, 5.020969, 5.014422, 5.00423, 4.989888, 
    4.970133, 4.947292, 4.912957, 4.877278, 4.842611, 4.811395, 4.785818, 
    4.767478, 4.757198, 4.755036, 4.760416, 4.772312, 4.789418, 4.810269, 
    4.833325, 4.857021, 4.879806, 4.900201, 4.916908, 4.928932, 4.935752,
  // height(16,28, 0-49)
    4.855995, 4.843037, 4.833967, 4.828879, 4.827681, 4.830082, 4.835604, 
    4.843608, 4.853339, 4.863991, 4.874754, 4.884873, 4.89369, 4.900697, 
    4.905574, 0, 5.000744, 5.006339, 5.013515, 5.021286, 5.028846, 5.028683, 
    5.02886, 5.027533, 5.025298, 5.021149, 5.014251, 5.003506, 4.988485, 
    4.967993, 4.944139, 4.909925, 4.874425, 4.840048, 4.809262, 4.78423, 
    4.766501, 4.756835, 4.75523, 4.761073, 4.773315, 4.790642, 4.811593, 
    4.834626, 4.858176, 4.88069, 4.900694, 4.916894, 4.928325, 4.934512,
  // height(16,29, 0-49)
    4.859104, 4.846059, 4.836926, 4.831833, 4.830725, 4.833347, 4.839246, 
    4.847798, 4.858232, 4.869702, 4.881335, 4.892307, 4.901924, 4.909692, 
    4.91538, 0, 4.999225, 5.004516, 5.011139, 5.018236, 5.025145, 5.026101, 
    5.027013, 5.026284, 5.024335, 5.02012, 5.012819, 5.001411, 4.985559, 
    4.964156, 4.939056, 4.904996, 4.869781, 4.835892, 4.805812, 4.781667, 
    4.764914, 4.756218, 4.755496, 4.762076, 4.774881, 4.792583, 4.813718, 
    4.836743, 4.86009, 4.882205, 4.90162, 4.917064, 4.927612, 4.93287,
  // height(16,30, 0-49)
    4.862476, 4.849107, 4.839384, 4.833349, 4.830894, 4.831782, 4.835658, 
    4.842111, 4.850717, 4.861089, 4.872904, 4.885905, 4.899866, 4.914509, 
    4.92938, 4.966947, 4.978901, 4.992922, 5.007429, 5.020907, 5.032383, 
    5.037577, 5.040587, 5.040208, 5.037008, 5.03027, 5.019615, 5.004519, 
    4.98509, 4.960538, 4.932539, 4.897691, 4.862357, 4.828973, 4.799906, 
    4.777106, 4.761838, 4.754601, 4.75519, 4.762854, 4.776481, 4.794729, 
    4.81613, 4.839152, 4.862225, 4.883802, 4.902434, 4.91689, 4.926324, 
    4.930448,
  // height(16,31, 0-49)
    4.866781, 4.853611, 4.844128, 4.83839, 4.836299, 4.837609, 4.84195, 
    4.848881, 4.857934, 4.868675, 4.880737, 4.893844, 4.9078, 4.922468, 
    4.937697, 4.967824, 4.977847, 4.991458, 5.004806, 5.016727, 5.02653, 
    5.031267, 5.033574, 5.032618, 5.028995, 5.021968, 5.011114, 4.995862, 
    4.976276, 4.951561, 4.923069, 4.889333, 4.855425, 4.823767, 4.796635, 
    4.775844, 4.762507, 4.756995, 4.759011, 4.767756, 4.782095, 4.800686, 
    4.822061, 4.844687, 4.867003, 4.887477, 4.904691, 4.917486, 4.925124, 
    4.927476,
  // height(16,32, 0-49)
    4.871303, 4.858335, 4.849073, 4.843582, 4.841766, 4.843366, 4.848002, 
    4.855215, 4.864517, 4.875458, 4.887661, 4.900854, 4.91489, 4.929732, 
    4.945438, 4.968321, 4.976445, 4.989829, 5.002178, 5.012691, 5.02094, 
    5.025236, 5.026824, 5.025161, 5.020825, 5.013091, 5.001563, 4.985727, 
    4.965698, 4.940761, 4.912001, 4.879725, 4.847709, 4.81828, 4.793566, 
    4.775197, 4.764112, 4.760547, 4.764117, 4.773983, 4.788996, 4.807811, 
    4.82897, 4.850946, 4.872193, 4.891208, 4.906636, 4.917415, 4.922964, 
    4.92335,
  // height(16,33, 0-49)
    4.875925, 4.863193, 4.854173, 4.84893, 4.847354, 4.84918, 4.854009, 
    4.861369, 4.870765, 4.881741, 4.893917, 4.907042, 4.921004, 4.935845, 
    4.951768, 4.968263, 4.974986, 4.988035, 4.999339, 5.008449, 5.015163, 
    5.01895, 5.019767, 5.017297, 5.012066, 5.003394, 4.99095, 4.974339, 
    4.95378, 4.928711, 4.900013, 4.869541, 4.839824, 4.813044, 4.791133, 
    4.775503, 4.766909, 4.765444, 4.770644, 4.78163, 4.797239, 4.816132, 
    4.836852, 4.857888, 4.877718, 4.894889, 4.908136, 4.916543, 4.919724, 
    4.917984,
  // height(16,34, 0-49)
    4.880545, 4.868095, 4.859358, 4.854384, 4.85305, 4.855068, 4.860024, 
    4.867435, 4.876794, 4.887642, 4.899608, 4.912449, 4.926073, 4.940565, 
    4.956202, 4.967526, 4.973517, 4.985917, 4.996002, 5.003626, 5.008771, 
    5.011938, 5.011914, 5.00858, 5.002374, 4.992685, 4.979272, 4.961896, 
    4.940898, 4.915932, 4.887727, 4.859404, 4.832354, 4.80857, 4.789754, 
    4.777088, 4.771133, 4.771847, 4.778687, 4.790736, 4.806821, 4.825599, 
    4.845624, 4.865399, 4.883441, 4.89837, 4.909048, 4.914743, 4.915324, 
    4.911375,
  // height(16,35, 0-49)
    4.885081, 4.87296, 4.864542, 4.85986, 4.858766, 4.86095, 4.865981, 
    4.873355, 4.882562, 4.893137, 4.904713, 4.917045, 4.930042, 4.943787, 
    4.95856, 4.96601, 4.971895, 4.98324, 4.991876, 4.997907, 5.001445, 
    5.003863, 5.002946, 4.998738, 4.991569, 4.980916, 4.966636, 4.948666, 
    4.927465, 4.902946, 4.87573, 4.849896, 4.825834, 4.805314, 4.78979, 
    4.780211, 4.776949, 4.779835, 4.788252, 4.801247, 4.817632, 4.836062, 
    4.855099, 4.87327, 4.889144, 4.901443, 4.909194, 4.911911, 4.909752, 
    4.903614,
  // height(16,36, 0-49)
    4.889462, 4.877706, 4.869629, 4.86524, 4.864367, 4.866679, 4.871722, 
    4.878978, 4.887927, 4.898099, 4.909123, 4.920747, 4.932858, 4.9455, 
    4.958887, 4.963627, 4.969875, 4.979753, 4.986724, 4.99107, 4.992982, 
    4.994537, 4.992704, 4.987673, 4.979637, 4.968187, 4.95327, 4.935, 
    4.913944, 4.890288, 4.86458, 4.841549, 4.820729, 4.803648, 4.791512, 
    4.78504, 4.784429, 4.789392, 4.799244, 4.812998, 4.82945, 4.847256, 
    4.864984, 4.881196, 4.894536, 4.903861, 4.908413, 4.907989, 4.90308, 
    4.894912,
  // height(16,37, 0-49)
    4.893633, 4.882252, 4.874506, 4.870379, 4.869679, 4.872052, 4.877029, 
    4.88408, 4.892673, 4.902333, 4.912676, 4.923434, 4.934464, 4.94574, 
    4.957366, 4.960308, 4.967186, 4.975255, 4.980393, 4.983005, 4.983312, 
    4.983918, 4.981193, 4.975446, 4.966719, 4.954725, 4.939501, 4.921314, 
    4.900814, 4.878473, 4.854766, 4.834799, 4.817393, 4.803834, 4.79508, 
    4.791636, 4.793539, 4.800397, 4.811465, 4.825723, 4.841955, 4.858814, 
    4.87489, 4.888796, 4.899277, 4.905368, 4.906568, 4.902996, 4.895502, 
    4.885627,
  // height(16,38, 0-49)
    4.897552, 4.886523, 4.879058, 4.875122, 4.874506, 4.876844, 4.881657, 
    4.888404, 4.896548, 4.905604, 4.915175, 4.924968, 4.934794, 4.944555, 
    4.954224, 4.956, 4.963574, 4.969604, 4.972828, 4.973719, 4.972487, 
    4.972108, 4.968562, 4.962262, 4.953082, 4.940866, 4.925722, 4.908052, 
    4.888546, 4.867952, 4.846678, 4.82996, 4.816054, 4.805999, 4.800521, 
    4.799932, 4.804125, 4.812616, 4.824606, 4.83905, 4.854722, 4.870285, 
    4.884364, 4.895648, 4.903024, 4.905744, 4.903603, 4.897072, 4.887355, 
    4.876265,
  // height(16,39, 0-49)
    4.901218, 4.89047, 4.88319, 4.879328, 4.878665, 4.880836, 4.885359, 
    4.891698, 4.899304, 4.907685, 4.916423, 4.925197, 4.933774, 4.94198, 
    4.94967, 4.950666, 4.958837, 4.962734, 4.964062, 4.96331, 4.960653, 
    4.959311, 4.955066, 4.948422, 4.939073, 4.926993, 4.912344, 4.89563, 
    4.877538, 4.859074, 4.840569, 4.827199, 4.81678, 4.810116, 4.807721, 
    4.809731, 4.815915, 4.825707, 4.838266, 4.852526, 4.867264, 4.881167, 
    4.892925, 4.901339, 4.905478, 4.904854, 4.89959, 4.890512, 4.879136, 
    4.86748,
  // height(16,40, 0-49)
    4.904684, 4.894101, 4.886861, 4.882905, 4.882024, 4.883858, 4.887946, 
    4.893749, 4.900727, 4.90837, 4.916239, 4.923985, 4.931323, 4.938021, 
    4.943837, 4.94427, 4.952819, 4.954637, 4.954183, 4.951932, 4.948014, 
    4.94579, 4.941018, 4.934273, 4.925064, 4.913489, 4.89974, 4.884389, 
    4.868077, 4.852043, 4.83653, 4.826512, 4.819475, 4.816006, 4.816424, 
    4.820711, 4.828525, 4.839235, 4.851963, 4.865639, 4.879057, 4.89096, 
    4.900132, 4.905531, 4.906458, 4.902721, 4.89478, 4.883789, 4.871507, 
    4.860053,
  // height(16,41, 0-49)
    4.908092, 4.897519, 4.89013, 4.885876, 4.884562, 4.88586, 4.889328, 
    4.894451, 4.90069, 4.907524, 4.914495, 4.921216, 4.927366, 4.932658, 
    4.93679, 4.93676, 4.945415, 4.945338, 4.943303, 4.939752, 4.934779, 
    4.93182, 4.926731, 4.920149, 4.911396, 4.900678, 4.888195, 4.874551, 
    4.86031, 4.846904, 4.834485, 4.827735, 4.823891, 4.823347, 4.826247, 
    4.832436, 4.841479, 4.852689, 4.86517, 4.87786, 4.889602, 4.899222, 
    4.905647, 4.908044, 4.905981, 4.899584, 4.889641, 4.877569, 4.865269, 
    4.854838,
  // height(16,42, 0-49)
    4.911717, 4.900965, 4.893209, 4.888418, 4.886428, 4.886953, 4.889586, 
    4.893843, 4.899196, 4.905123, 4.911144, 4.91684, 4.921854, 4.925863, 
    4.928534, 4.928086, 4.936563, 4.934877, 4.931522, 4.926918, 4.92114, 
    4.917643, 4.912477, 4.906325, 4.89833, 4.888782, 4.877871, 4.866199, 
    4.854226, 4.843546, 4.834213, 4.830557, 4.829648, 4.831701, 4.836706, 
    4.84439, 4.854242, 4.865532, 4.877361, 4.888703, 4.898479, 4.905645, 
    4.909317, 4.908913, 4.904303, 4.895933, 4.88486, 4.872675, 4.861303, 
    4.852696,
  // height(16,43, 0-49)
    4.915979, 4.904849, 4.896491, 4.890907, 4.887977, 4.887463, 4.889009, 
    4.892169, 4.896441, 4.901309, 4.90628, 4.910909, 4.914815, 4.91765, 
    4.919073, 4.918221, 4.926271, 4.923316, 4.918942, 4.91356, 4.907251, 
    4.903452, 4.898461, 4.892997, 4.886028, 4.877912, 4.868806, 4.859283, 
    4.849682, 4.841722, 4.835365, 4.834563, 4.836274, 4.840557, 4.847266, 
    4.856031, 4.866275, 4.877251, 4.888074, 4.897788, 4.905428, 4.910126, 
    4.911233, 4.908454, 4.901965, 4.892494, 4.881298, 4.870026, 4.860497, 
    4.854419,
  // height(16,44, 0-49)
    4.921442, 4.909743, 4.900558, 4.893926, 4.889781, 4.887942, 4.888114, 
    4.889902, 4.892839, 4.89643, 4.900186, 4.903648, 4.906418, 4.90814, 
    4.908477, 4.907215, 4.914638, 4.910761, 4.905677, 4.899805, 4.89325, 
    4.8894, 4.884832, 4.880281, 4.874562, 4.868074, 4.860928, 4.853642, 
    4.846432, 4.841105, 4.837529, 4.839285, 4.843264, 4.849389, 4.857398, 
    4.866843, 4.877102, 4.887429, 4.896988, 4.90492, 4.910418, 4.912833, 
    4.911785, 4.907272, 4.89976, 4.890192, 4.879921, 4.87054, 4.863652, 
    4.860648,
  // height(16,45, 0-49)
    4.928774, 4.916354, 4.906143, 4.89823, 4.892606, 4.889152, 4.887639, 
    4.887737, 4.889032, 4.891066, 4.893369, 4.895489, 4.897025, 4.897626, 
    4.89697, 4.895264, 4.901911, 4.897421, 4.891912, 4.885824, 4.879295, 
    4.875637, 4.871709, 4.868249, 4.863946, 4.85921, 4.854095, 4.849058, 
    4.844183, 4.84133, 4.840287, 4.844272, 4.850154, 4.857734, 4.866662, 
    4.876428, 4.886393, 4.895836, 4.903998, 4.910158, 4.913705, 4.914233, 
    4.911644, 4.906223, 4.898661, 4.890035, 4.881682, 4.875031, 4.871395, 
    4.871812,
  // height(16,46, 0-49)
    4.93868, 4.925437, 4.914054, 4.904667, 4.897326, 4.891982, 4.888477, 
    4.886553, 4.885867, 4.886013, 4.886566, 4.887105, 4.88724, 4.886635, 
    4.884993, 4.88277, 4.888525, 4.883657, 4.877955, 4.871884, 4.865617, 
    4.862357, 4.859235, 4.856978, 4.854181, 4.851244, 4.848159, 4.845309, 
    4.842661, 4.842082, 4.843284, 4.849162, 4.856587, 4.865265, 4.874779, 
    4.88458, 4.894042, 4.902493, 4.909286, 4.913868, 4.915846, 4.915076, 
    4.911729, 4.906325, 4.899712, 4.892994, 4.887399, 4.884111, 4.884117, 
    4.888099,
  // height(16,47, 0-49)
    4.951799, 4.937706, 4.925067, 4.914071, 4.904827, 4.897355, 4.891575, 
    4.887312, 4.884302, 4.88222, 4.880702, 4.879376, 4.87789, 4.875928, 
    4.873226, 4.870365, 4.875134, 4.870023, 4.864284, 4.858397, 4.852556, 
    4.849838, 4.847615, 4.846592, 4.845309, 4.844142, 4.843019, 4.842241, 
    4.841671, 4.843141, 4.846299, 4.853746, 4.862389, 4.871863, 4.881702, 
    4.891355, 4.900224, 4.907723, 4.913341, 4.916712, 4.917672, 4.916331, 
    4.913086, 4.908631, 4.903881, 4.899878, 4.897662, 4.89813, 4.901938, 
    4.909441,
  // height(16,48, 0-49)
    4.968619, 4.953721, 4.939814, 4.927141, 4.915872, 4.906098, 4.897817, 
    4.890945, 4.885314, 4.880691, 4.876794, 4.873322, 4.869973, 4.866468, 
    4.862566, 4.858901, 4.862593, 4.857264, 4.85155, 4.845926, 4.840598, 
    4.838478, 4.837162, 4.837315, 4.837472, 4.837968, 4.838675, 4.839813, 
    4.841158, 4.844455, 4.849295, 4.858031, 4.867624, 4.877662, 4.887666, 
    4.897097, 4.905418, 4.912148, 4.916932, 4.919597, 4.920197, 4.91906, 
    4.916761, 4.914085, 4.911936, 4.911226, 4.912759, 4.917141, 4.92471, 
    4.935537,
  // height(16,49, 0-49)
    4.997341, 4.981748, 4.96641, 4.95162, 4.937616, 4.924573, 4.9126, 
    4.901742, 4.89198, 4.883229, 4.875348, 4.868152, 4.861418, 4.854907, 
    4.848384, 4.843278, 4.852906, 4.845834, 4.83861, 4.832042, 4.8264, 
    4.827126, 4.82929, 4.833854, 4.837558, 4.840845, 4.843235, 4.844953, 
    4.845376, 4.847987, 4.852074, 4.862319, 4.872993, 4.88364, 4.893794, 
    4.902972, 4.910752, 4.916822, 4.921046, 4.923507, 4.924527, 4.92465, 
    4.9246, 4.925184, 4.927189, 4.931278, 4.93792, 4.947337, 4.959503, 
    4.974175,
  // height(17,0, 0-49)
    4.932086, 4.910845, 4.892358, 4.876889, 4.864563, 4.855368, 4.849143, 
    4.845583, 4.844279, 4.84473, 4.846404, 4.84877, 4.851345, 4.853716, 
    4.855547, 4.85666, 4.858193, 4.857396, 4.855773, 4.853347, 4.850139, 
    4.846555, 4.84232, 4.837674, 4.832701, 4.827689, 4.822936, 4.818818, 
    4.815685, 4.813998, 4.813952, 4.81605, 4.819995, 4.825649, 4.832704, 
    4.840699, 4.849057, 4.857137, 4.864295, 4.869975, 4.873768, 4.8755, 
    4.875279, 4.87353, 4.870981, 4.868604, 4.867512, 4.868828, 4.873548, 
    4.882422,
  // height(17,1, 0-49)
    4.927293, 4.906449, 4.888511, 4.873724, 4.862199, 4.853904, 4.848652, 
    4.846119, 4.845862, 4.847353, 4.850029, 4.853331, 4.856744, 4.859819, 
    4.862175, 4.863629, 4.866576, 4.865678, 4.863865, 4.861151, 4.857523, 
    4.853695, 4.849001, 4.843752, 4.837935, 4.831862, 4.825829, 4.820256, 
    4.815511, 4.812222, 4.810579, 4.811505, 4.814435, 4.819283, 4.825787, 
    4.83351, 4.841879, 4.850229, 4.85787, 4.864164, 4.868599, 4.870879, 
    4.870985, 4.869229, 4.866257, 4.863015, 4.860652, 4.860381, 4.863338, 
    4.87043,
  // height(17,2, 0-49)
    4.925047, 4.904743, 4.887443, 4.873371, 4.862625, 4.855145, 4.85073, 
    4.849032, 4.849593, 4.851871, 4.855292, 4.859291, 4.863336, 4.866961, 
    4.86975, 4.871462, 4.875763, 4.874875, 4.873009, 4.870171, 4.866305, 
    4.862421, 4.857438, 4.851728, 4.845177, 4.838098, 4.830777, 4.823665, 
    4.817146, 4.812004, 4.80843, 4.807797, 4.809296, 4.812929, 4.81851, 
    4.825661, 4.833847, 4.842411, 4.850638, 4.857832, 4.863382, 4.866856, 
    4.868075, 4.867185, 4.864679, 4.861393, 4.858432, 4.857043, 4.85846, 
    4.863751,
  // height(17,3, 0-49)
    4.924704, 4.905055, 4.888456, 4.875116, 4.865107, 4.858351, 4.854629, 
    4.85358, 4.85474, 4.85757, 4.861506, 4.865989, 4.870497, 4.874556, 
    4.877724, 4.879621, 4.88518, 4.884454, 4.882708, 4.879936, 4.876042, 
    4.872316, 4.867249, 4.861258, 4.854124, 4.846151, 4.837596, 4.828926, 
    4.820539, 4.813347, 4.807551, 4.805, 4.804668, 4.806671, 4.810932, 
    4.817171, 4.824917, 4.833555, 4.842372, 4.850632, 4.85764, 4.862832, 
    4.865854, 4.866643, 4.865483, 4.863023, 4.860238, 4.858329, 4.858582, 
    4.862187,
  // height(17,4, 0-49)
    4.925554, 4.906652, 4.890803, 4.878195, 4.868879, 4.862763, 4.859605, 
    4.859044, 4.860619, 4.863809, 4.868073, 4.87288, 4.877728, 4.882148, 
    4.885689, 4.887709, 4.894379, 4.894003, 4.892564, 4.890065, 4.886366, 
    4.88302, 4.878093, 4.872019, 4.8645, 4.855797, 4.846127, 4.835956, 
    4.825689, 4.816328, 4.808094, 4.803315, 4.800786, 4.800761, 4.803308, 
    4.808267, 4.815266, 4.823757, 4.833058, 4.842415, 4.85107, 4.858335, 
    4.863684, 4.866829, 4.867804, 4.867007, 4.865207, 4.863475, 4.863067, 
    4.865251,
  // height(17,5, 0-49)
    4.926895, 4.908814, 4.893754, 4.881882, 4.873228, 4.86768, 4.86499, 
    4.864796, 4.866652, 4.870066, 4.874532, 4.879558, 4.884674, 4.889433, 
    4.893384, 4.89547, 4.903042, 4.903224, 4.902287, 4.900254, 4.896966, 
    4.894212, 4.889642, 4.883701, 4.87602, 4.866802, 4.856206, 4.844675, 
    4.832611, 4.821059, 4.810258, 4.803021, 4.79799, 4.795586, 4.796041, 
    4.799346, 4.805257, 4.813318, 4.822897, 4.833249, 4.843571, 4.853073, 
    4.861067, 4.867047, 4.870778, 4.872372, 4.872322, 4.871489, 4.871013, 
    4.872166,
  // height(17,6, 0-49)
    4.928093, 4.910898, 4.896666, 4.885541, 4.877535, 4.872518, 4.870237, 
    4.870338, 4.872396, 4.875957, 4.880558, 4.885754, 4.891115, 4.89623, 
    4.900664, 4.902766, 4.910966, 4.911911, 4.911652, 4.910261, 4.907574, 
    4.905591, 4.901582, 4.895983, 4.888383, 4.878903, 4.867634, 4.85497, 
    4.841294, 4.827643, 4.814258, 4.804423, 4.796666, 4.791592, 4.789618, 
    4.790914, 4.795382, 4.802684, 4.812258, 4.823384, 4.835237, 4.84695, 
    4.857692, 4.866757, 4.873649, 4.878177, 4.88052, 4.881258, 4.881336, 
    4.881945,
  // height(17,7, 0-49)
    4.928635, 4.912382, 4.89902, 4.888669, 4.88132, 4.87683, 4.874942, 
    4.875315, 4.877554, 4.88124, 4.88596, 4.891318, 4.896939, 4.902454, 
    4.907468, 4.909537, 4.918041, 4.919922, 4.920493, 4.919884, 4.91795, 
    4.916876, 4.913595, 4.908529, 4.901253, 4.891789, 4.880151, 4.866659, 
    4.851659, 4.836112, 4.820251, 4.80779, 4.797184, 4.789228, 4.78455, 
    4.783514, 4.786196, 4.792386, 4.801616, 4.813207, 4.826326, 4.840052, 
    4.853444, 4.865614, 4.875832, 4.883608, 4.8888, 4.891662, 4.892874, 
    4.893465,
  // height(17,8, 0-49)
    4.928143, 4.912886, 4.900441, 4.890904, 4.884245, 4.880311, 4.878841, 
    4.87951, 4.88195, 4.885783, 4.890644, 4.89619, 4.902103, 4.908071, 
    4.913764, 4.915773, 4.92422, 4.927168, 4.928677, 4.928949, 4.927879, 
    4.927794, 4.925365, 4.920992, 4.914267, 4.905104, 4.893435, 4.879482, 
    4.863534, 4.846408, 4.828302, 4.813304, 4.799834, 4.788882, 4.781299, 
    4.777662, 4.778239, 4.782969, 4.791487, 4.803172, 4.817198, 4.83261, 
    4.848373, 4.863461, 4.876935, 4.88804, 4.896313, 4.901678, 4.904503, 
    4.905589,
  // height(17,9, 0-49)
    4.926387, 4.91217, 4.900692, 4.892024, 4.88611, 4.882786, 4.881791, 
    4.882813, 4.88551, 4.889541, 4.894586, 4.900361, 4.906602, 4.913068, 
    4.919524, 4.921489, 4.929521, 4.933596, 4.936105, 4.937315, 4.937177, 
    4.938101, 4.936598, 4.933035, 4.927056, 4.918464, 4.90711, 4.893102, 
    4.876647, 4.85835, 4.838352, 4.821018, 4.804783, 4.790828, 4.780226, 
    4.773788, 4.771987, 4.774931, 4.782368, 4.793742, 4.808257, 4.824928, 
    4.84266, 4.860311, 4.876772, 4.891061, 4.902427, 4.910475, 4.915247, 
    4.917273,
  // height(17,10, 0-49)
    4.923273, 4.910128, 4.899665, 4.891922, 4.886822, 4.884184, 4.883743, 
    4.885196, 4.888224, 4.892519, 4.897807, 4.903848, 4.910443, 4.917434, 
    4.924696, 4.92671, 4.934017, 4.939202, 4.942721, 4.944888, 4.945706, 
    4.947608, 4.947049, 4.944363, 4.939278, 4.931495, 4.920787, 4.907132, 
    4.890639, 4.871647, 4.850207, 4.83084, 4.812048, 4.795187, 4.781552, 
    4.772192, 4.767801, 4.768667, 4.774671, 4.785334, 4.799887, 4.817338, 
    4.836549, 4.856289, 4.875316, 4.892464, 4.906739, 4.917458, 4.924351, 
    4.92766,
  // height(17,11, 0-49)
    4.918819, 4.906762, 4.897353, 4.890594, 4.886381, 4.884509, 4.884711, 
    4.886684, 4.890129, 4.89476, 4.90034, 4.906679, 4.913639, 4.921144, 
    4.929193, 4.931473, 4.937835, 4.944029, 4.948521, 4.951626, 4.953395, 
    4.95619, 4.956545, 4.954758, 4.950663, 4.943872, 4.934094, 4.921172, 
    4.905105, 4.885919, 4.863553, 4.842531, 4.821484, 4.801915, 4.785327, 
    4.773007, 4.765884, 4.764438, 4.768693, 4.778259, 4.792406, 4.810146, 
    4.830305, 4.851591, 4.872667, 4.89222, 4.909069, 4.922284, 4.931321, 
    4.936136,
  // height(17,12, 0-49)
    4.913151, 4.902174, 4.89384, 4.888111, 4.884847, 4.883822, 4.884756, 
    4.887339, 4.891278, 4.896312, 4.90223, 4.908882, 4.91619, 4.924158, 
    4.932895, 4.935816, 4.941145, 4.948177, 4.953555, 4.957557, 4.960253, 
    4.96382, 4.965019, 4.964102, 4.961035, 4.955356, 4.946728, 4.934856, 
    4.919626, 4.900735, 4.877989, 4.855725, 4.832791, 4.810797, 4.791426, 
    4.776199, 4.766277, 4.762349, 4.764593, 4.772719, 4.786045, 4.803592, 
    4.82417, 4.846443, 4.869005, 4.890441, 4.90943, 4.924849, 4.935921, 
    4.942349,
  // height(17,13, 0-49)
    4.906466, 4.896542, 4.889278, 4.884605, 4.882339, 4.882226, 4.883963, 
    4.887234, 4.891738, 4.897228, 4.903514, 4.91048, 4.918095, 4.926425, 
    4.93566, 4.939777, 4.944144, 4.951789, 4.95794, 4.962779, 4.966364, 
    4.970561, 4.972504, 4.972393, 4.970335, 4.96582, 4.958477, 4.947888, 
    4.933827, 4.915659, 4.893061, 4.869974, 4.845552, 4.821473, 4.799566, 
    4.781562, 4.768855, 4.762346, 4.762383, 4.768782, 4.78092, 4.797838, 
    4.818337, 4.841057, 4.864547, 4.887329, 4.907979, 4.925239, 4.938151, 
    4.946199,
  // height(17,14, 0-49)
    4.899024, 4.89009, 4.883871, 4.880249, 4.879004, 4.879846, 4.882438, 
    4.886447, 4.891568, 4.897552, 4.90422, 4.911483, 4.919337, 4.927886, 
    4.937351, 4.943377, 4.947018, 4.955034, 4.961828, 4.967443, 4.971882, 
    4.976558, 4.979132, 4.979733, 4.97862, 4.975255, 4.969245, 4.960069, 
    4.947399, 4.930287, 4.908312, 4.884778, 4.859268, 4.833473, 4.809331, 
    4.788751, 4.773347, 4.764234, 4.761935, 4.766388, 4.777039, 4.792955, 
    4.812939, 4.835619, 4.859524, 4.883137, 4.904978, 4.923697, 4.9382, 
    4.947796,
  // height(17,15, 0-49)
    4.891112, 4.883087, 4.877852, 4.875248, 4.875012, 4.876813, 4.880279, 
    4.885053, 4.890813, 4.897305, 4.904356, 4.911882, 4.919893, 4.928493, 
    4.93788, 4.946609, 4.949912, 4.958069, 4.965397, 4.97174, 4.97701, 
    4.982026, 4.985116, 4.986323, 4.986053, 4.983757, 4.979042, 4.971297, 
    4.960118, 4.944283, 4.923313, 4.899639, 4.873401, 4.84626, 4.820212, 
    4.797309, 4.779364, 4.767699, 4.763014, 4.76538, 4.774317, 4.788934, 
    4.808044, 4.830278, 4.854156, 4.87815, 4.900752, 4.920557, 4.936386, 
    4.947409,
  // height(17,16, 0-49)
    4.883029, 4.875806, 4.871468, 4.869812, 4.870532, 4.873254, 4.877571, 
    4.883094, 4.889482, 4.896476, 4.903892, 4.911646, 4.919736, 4.928235, 
    4.937255, 4.949426, 4.952873, 4.96102, 4.968817, 4.975876, 4.981983, 
    4.987225, 4.990734, 4.992444, 4.992887, 4.991526, 4.987975, 4.981569, 
    4.971848, 4.957378, 4.937684, 4.914083, 4.887414, 4.859268, 4.831649, 
    4.806712, 4.786437, 4.772339, 4.765296, 4.765512, 4.772596, 4.785703, 
    4.803671, 4.825141, 4.84864, 4.872643, 4.89564, 4.916207, 4.933103, 
    4.945402,
  // height(17,17, 0-49)
    4.875055, 4.868514, 4.864955, 4.864135, 4.86571, 4.869261, 4.87435, 
    4.880558, 4.88753, 4.89499, 4.902754, 4.910722, 4.918859, 4.927171, 
    4.935653, 4.951737, 4.955822, 4.963933, 4.972224, 4.980051, 4.987048, 
    4.992446, 4.996313, 4.998434, 4.999444, 4.99883, 4.99623, 4.990953, 
    4.982525, 4.969369, 4.951089, 4.927674, 4.900793, 4.871935, 4.843071, 
    4.816412, 4.794065, 4.777717, 4.768412, 4.766494, 4.771667, 4.783143, 
    4.799794, 4.820279, 4.843141, 4.866875, 4.889984, 4.911039, 4.928771, 
    4.942188,
  // height(17,18, 0-49)
    4.867438, 4.861432, 4.858498, 4.858359, 4.860627, 4.864854, 4.870573, 
    4.87735, 4.884819, 4.892704, 4.900818, 4.909043, 4.917301, 4.925497, 
    4.93346, 4.953443, 4.958536, 4.966762, 4.975693, 4.984436, 4.992451, 
    4.997995, 5.002215, 5.004687, 5.006111, 5.006001, 5.004041, 4.999564, 
    4.992125, 4.980086, 4.963223, 4.940009, 4.913056, 4.88373, 4.853928, 
    4.825867, 4.801744, 4.783382, 4.771981, 4.768018, 4.771304, 4.781112, 
    4.796357, 4.815728, 4.83779, 4.861065, 4.884079, 4.905415, 4.923792, 
    4.938173,
  // height(17,19, 0-49)
    4.860362, 4.854715, 4.852209, 4.85253, 4.855262, 4.859932, 4.866065, 
    4.87323, 4.881079, 4.889356, 4.89789, 4.906549, 4.915184, 4.923564, 
    4.931289, 4.954461, 4.960647, 4.969331, 4.979218, 4.989158, 4.998429, 
    5.004205, 5.008854, 5.011667, 5.013352, 5.01345, 5.011711, 5.007554, 
    5.000636, 4.989366, 4.973771, 4.950686, 4.92374, 4.894152, 4.863704, 
    4.834578, 4.809007, 4.788918, 4.775646, 4.769795, 4.771284, 4.77946, 
    4.793291, 4.811497, 4.83268, 4.855388, 4.878173, 4.899641, 4.918513, 
    4.933718,
  // height(17,20, 0-49)
    4.854655, 4.849918, 4.84861, 4.850455, 4.855026, 4.861779, 4.870096, 
    4.879328, 4.888843, 4.898059, 4.906477, 4.913717, 4.919533, 4.923843, 
    4.926725, 0, 4.976701, 4.980468, 4.985542, 4.99134, 4.997496, 5.000072, 
    5.003079, 5.005518, 5.008004, 5.009818, 5.010391, 5.008807, 5.004483, 
    4.995662, 4.982596, 4.960472, 4.934066, 4.904542, 4.873656, 4.843603, 
    4.816685, 4.794946, 4.779853, 4.772143, 4.771838, 4.778371, 4.790754, 
    4.807751, 4.827991, 4.850053, 4.872515, 4.894001, 4.913239, 4.929135,
  // height(17,21, 0-49)
    4.849359, 4.844958, 4.844018, 4.846222, 4.851108, 4.858102, 4.866564, 
    4.875849, 4.885345, 4.89451, 4.90289, 4.910137, 4.916014, 4.920402, 
    4.923314, 0, 4.978804, 4.983113, 4.98882, 4.995245, 5.001908, 5.003341, 
    5.005481, 5.007151, 5.009163, 5.010862, 5.011708, 5.010763, 5.007414, 
    4.999859, 4.988595, 4.967202, 4.941577, 4.912706, 4.882171, 4.852049, 
    4.824604, 4.801916, 4.785548, 4.776368, 4.774518, 4.77953, 4.790494, 
    4.806223, 4.825388, 4.846598, 4.868461, 4.889622, 4.908823, 4.924966,
  // height(17,22, 0-49)
    4.84491, 4.840719, 4.840024, 4.842488, 4.847629, 4.854852, 4.863504, 
    4.872935, 4.882536, 4.891777, 4.900223, 4.907533, 4.913461, 4.917856, 
    4.920673, 0, 4.980448, 4.985187, 4.991485, 4.998569, 5.005846, 5.006361, 
    5.007894, 5.009054, 5.010793, 5.012468, 5.013533, 5.01302, 5.010294, 
    5.003533, 4.9935, 4.972336, 4.947056, 4.918531, 4.888209, 4.858057, 
    4.830273, 4.806931, 4.789643, 4.779356, 4.776308, 4.780115, 4.789931, 
    4.804622, 4.822892, 4.843383, 4.864727, 4.885594, 4.904738, 4.921063,
  // height(17,23, 0-49)
    4.841343, 4.837268, 4.836722, 4.839362, 4.844692, 4.852111, 4.860959, 
    4.870574, 4.880348, 4.889748, 4.898341, 4.905778, 4.911798, 4.916217, 
    4.918941, 0, 4.982242, 4.987259, 4.993968, 5.001531, 5.009266, 5.00898, 
    5.009981, 5.010692, 5.012161, 5.013753, 5.014909, 5.014637, 5.012286, 
    5.006017, 4.996813, 4.975653, 4.950515, 4.922195, 4.892049, 4.861947, 
    4.834018, 4.810307, 4.792441, 4.781416, 4.77753, 4.780464, 4.789426, 
    4.803322, 4.820889, 4.840794, 4.86169, 4.882262, 4.901279, 4.917653,
  // height(17,24, 0-49)
    4.838642, 4.834622, 4.834155, 4.836901, 4.842365, 4.849943, 4.858972, 
    4.868788, 4.878774, 4.888392, 4.897195, 4.904826, 4.911006, 4.915524, 
    4.918251, 0, 4.984415, 4.98959, 4.996536, 5.004384, 5.012406, 5.011586, 
    5.012234, 5.012639, 5.013902, 5.015387, 5.016535, 5.016338, 5.014139, 
    5.008089, 4.999325, 4.978053, 4.952898, 4.924624, 4.894527, 4.864416, 
    4.836373, 4.812413, 4.794162, 4.782639, 4.778178, 4.7805, 4.788852, 
    4.80217, 4.819218, 4.838678, 4.859221, 4.879544, 4.898427, 4.914783,
  // height(17,25, 0-49)
    4.836769, 4.832759, 4.832325, 4.83513, 4.840688, 4.8484, 4.857604, 
    4.867634, 4.877865, 4.887749, 4.896824, 4.904718, 4.911138, 4.915858, 
    4.918736, 0, 4.986551, 4.991792, 4.998822, 5.006766, 5.014881, 5.013883, 
    5.014416, 5.014708, 5.015873, 5.017272, 5.018345, 5.018085, 5.015834, 
    5.009744, 5.001011, 4.979569, 4.954289, 4.925926, 4.895759, 4.865575, 
    4.83743, 4.813322, 4.794866, 4.783079, 4.778309, 4.780292, 4.788291, 
    4.801262, 4.817979, 4.837139, 4.85742, 4.877531, 4.89625, 4.912501,
  // height(17,26, 0-49)
    4.835672, 4.83165, 4.831218, 4.834058, 4.839693, 4.847535, 4.856926, 
    4.867199, 4.877722, 4.887929, 4.897342, 4.905571, 4.912312, 4.917341, 
    4.920526, 0, 4.988527, 4.993752, 5.000716, 5.008561, 5.016568, 5.015782, 
    5.016457, 5.016857, 5.018059, 5.019417, 5.020375, 5.019933, 5.017445, 
    5.011068, 5.001957, 4.980327, 4.954838, 4.92627, 4.895921, 4.865594, 
    4.837351, 4.813177, 4.794672, 4.782838, 4.778008, 4.779906, 4.787796, 
    4.800632, 4.817194, 4.836185, 4.856286, 4.876206, 4.894732, 4.910787,
  // height(17,27, 0-49)
    4.835305, 4.831254, 4.830816, 4.833688, 4.83941, 4.847407, 4.857031, 
    4.86761, 4.878496, 4.889104, 4.898934, 4.907572, 4.914705, 4.920119, 
    4.923718, 0, 4.990418, 4.995515, 5.002238, 5.00977, 5.01746, 5.017213, 
    5.018252, 5.01895, 5.020303, 5.021653, 5.022446, 5.021699, 5.018786, 
    5.011879, 5.002003, 4.980161, 4.954391, 4.925523, 4.894915, 4.864421, 
    4.836125, 4.812012, 4.793656, 4.782018, 4.777392, 4.779467, 4.787487, 
    4.800394, 4.816962, 4.835893, 4.855869, 4.875599, 4.893869, 4.909608,
  // height(17,28, 0-49)
    4.835628, 4.831538, 4.831094, 4.834014, 4.839862, 4.848079, 4.85802, 
    4.869009, 4.880377, 4.891504, 4.90185, 4.910967, 4.91853, 4.924347, 
    4.928369, 0, 4.992599, 4.997404, 5.003668, 5.010651, 5.017807, 5.018314, 
    5.019859, 5.020988, 5.022568, 5.023917, 5.02448, 5.023301, 5.019778, 
    5.01211, 5.00112, 4.979014, 4.952876, 4.923621, 4.892708, 4.862062, 
    4.833807, 4.809922, 4.791938, 4.780753, 4.776589, 4.779086, 4.787449, 
    4.8006, 4.817302, 4.836254, 4.856133, 4.875648, 4.893589, 4.908889,
  // height(17,29, 0-49)
    4.836607, 4.832465, 4.832018, 4.835017, 4.841056, 4.849597, 4.859998, 
    4.871566, 4.883592, 4.8954, 4.906381, 4.916035, 4.924014, 4.930147, 
    4.934448, 0, 4.994762, 4.999057, 5.004619, 5.010811, 5.01722, 5.01852, 
    5.020604, 5.022212, 5.02405, 5.025388, 5.025658, 5.023925, 5.019612, 
    5.010951, 4.998516, 4.976011, 4.949397, 4.919718, 4.888555, 4.857924, 
    4.829979, 4.806665, 4.789436, 4.779088, 4.77575, 4.778986, 4.787952, 
    4.80154, 4.818505, 4.837532, 4.857296, 4.876508, 4.89396, 4.908601,
  // height(17,30, 0-49)
    4.837832, 4.833149, 4.831962, 4.833973, 4.838768, 4.84586, 4.854743, 
    4.86493, 4.875998, 4.887613, 4.899509, 4.911485, 4.923332, 4.93478, 
    4.945404, 4.975517, 4.979926, 4.9902, 5.001615, 5.01291, 5.023316, 
    5.028723, 5.033325, 5.036073, 5.037669, 5.037555, 5.035443, 5.030748, 
    5.023216, 5.011344, 4.995587, 4.971336, 4.943355, 4.912786, 4.881282, 
    4.850867, 4.823629, 4.801392, 4.785451, 4.776451, 4.77439, 4.778745, 
    4.788615, 4.802867, 4.820241, 4.839418, 4.859073, 4.87792, 4.894762, 
    4.908581,
  // height(17,31, 0-49)
    4.840512, 4.836057, 4.835127, 4.837435, 4.842564, 4.85002, 4.85927, 
    4.869801, 4.881155, 4.892956, 4.904926, 4.916868, 4.928643, 4.940125, 
    4.951134, 4.976396, 4.981072, 4.990958, 5.001443, 5.011515, 5.020609, 
    5.025819, 5.029953, 5.032291, 5.033554, 5.033181, 5.03083, 5.025838, 
    5.017842, 5.005279, 4.988306, 4.964038, 4.936157, 4.905926, 4.875092, 
    4.845701, 4.81979, 4.799075, 4.784719, 4.777233, 4.77651, 4.781954, 
    4.792624, 4.80736, 4.824892, 4.843892, 4.863036, 4.881039, 4.896733, 
    4.90915,
  // height(17,32, 0-49)
    4.84394, 4.839687, 4.838961, 4.84147, 4.8468, 4.854445, 4.863869, 
    4.874544, 4.886004, 4.897867, 4.909857, 4.921802, 4.933619, 4.9453, 
    4.956847, 4.976905, 4.981479, 4.991234, 5.00101, 5.010061, 5.018018, 
    5.023118, 5.026866, 5.028792, 5.02958, 5.028664, 5.025671, 5.019921, 
    5.011018, 4.997434, 4.979104, 4.954812, 4.927166, 4.897542, 4.867736, 
    4.839773, 4.815597, 4.796778, 4.784322, 4.7786, 4.779403, 4.786065, 
    4.797607, 4.812852, 4.830517, 4.849267, 4.867775, 4.88477, 4.899115, 
    4.909908,
  // height(17,33, 0-49)
    4.848188, 4.844136, 4.843581, 4.846228, 4.851653, 4.859349, 4.868777, 
    4.879411, 4.890791, 4.902544, 4.914413, 4.926251, 4.938032, 4.949833, 
    4.961806, 4.976944, 4.981427, 4.991122, 5.000261, 5.008378, 5.015282, 
    5.02028, 5.023657, 5.025142, 5.025333, 5.023657, 5.019734, 5.012911, 
    5.002809, 4.988014, 4.968327, 4.944061, 4.916827, 4.88808, 4.859641, 
    4.83347, 4.811376, 4.794761, 4.784458, 4.780696, 4.783165, 4.791138, 
    4.803601, 4.819355, 4.837107, 4.855516, 4.87325, 4.889057, 4.901842, 
    4.910791,
  // height(17,34, 0-49)
    4.853289, 4.849438, 4.849027, 4.851749, 4.857172, 4.864788, 4.874062, 
    4.88448, 4.895594, 4.907053, 4.91862, 4.930174, 4.941731, 4.953428, 
    4.965522, 4.976438, 4.981064, 4.990592, 4.999053, 5.006239, 5.012118, 
    5.01695, 5.019924, 5.020919, 5.020409, 5.017825, 5.01279, 5.004707, 
    4.993249, 4.9772, 4.956297, 4.932189, 4.905595, 4.878024, 4.85128, 
    4.827223, 4.8075, 4.793324, 4.785354, 4.783679, 4.787896, 4.797219, 
    4.810601, 4.826828, 4.844588, 4.862535, 4.879337, 4.893764, 4.904784, 
    4.911689,
  // height(17,35, 0-49)
    4.859222, 4.855562, 4.855252, 4.857974, 4.863289, 4.870693, 4.879658, 
    4.889689, 4.900362, 4.911344, 4.922421, 4.933497, 4.944608, 4.955915, 
    4.967728, 4.975316, 4.980386, 4.989532, 4.997201, 5.003416, 5.00826, 
    5.012824, 5.015333, 5.015789, 5.014503, 5.010921, 5.004682, 4.995273, 
    4.982435, 4.965222, 4.943371, 4.919636, 4.893962, 4.867884, 4.843148, 
    4.82148, 4.804347, 4.792766, 4.787225, 4.787683, 4.793653, 4.804296, 
    4.81854, 4.835147, 4.852794, 4.870125, 4.885816, 4.898671, 4.907736, 
    4.912441,
  // height(17,36, 0-49)
    4.865902, 4.862398, 4.862123, 4.86475, 4.869839, 4.876892, 4.885399, 
    4.894885, 4.904952, 4.915292, 4.925711, 4.936127, 4.946576, 4.957216, 
    4.968345, 4.973502, 4.979285, 4.987776, 4.994511, 4.999691, 5.003481, 
    5.007654, 5.009626, 5.009497, 5.007393, 5.002791, 4.995346, 4.984653, 
    4.97054, 4.952381, 4.929957, 4.90688, 4.882451, 4.858187, 4.835741, 
    4.816682, 4.802279, 4.793364, 4.790259, 4.792812, 4.800456, 4.812315, 
    4.827287, 4.844121, 4.861478, 4.877997, 4.892375, 4.903469, 4.910425, 
    4.912837,
  // height(17,37, 0-49)
    4.873171, 4.869758, 4.869428, 4.871847, 4.876582, 4.883149, 4.891055, 
    4.899855, 4.909174, 4.918733, 4.928355, 4.93796, 4.947573, 4.957314, 
    4.967422, 4.970922, 4.977585, 4.98515, 4.990809, 4.994896, 4.997612, 
    5.001259, 5.002623, 5.001882, 4.998955, 4.993373, 4.984812, 4.972988, 
    4.957819, 4.939039, 4.916505, 4.894428, 4.871589, 4.849447, 4.829532, 
    4.813232, 4.801623, 4.795353, 4.794603, 4.799121, 4.808279, 4.821166, 
    4.836657, 4.853489, 4.870317, 4.885788, 4.898634, 4.907787, 4.91253, 
    4.912643,
  // height(17,38, 0-49)
    4.880799, 4.877385, 4.876884, 4.878968, 4.88322, 4.889169, 4.896352, 
    4.904349, 4.912816, 4.921493, 4.930215, 4.938902, 4.947552, 4.956231, 
    4.965086, 4.967517, 4.975098, 4.981501, 4.985966, 4.988914, 4.990543, 
    4.993541, 4.994239, 4.992883, 4.989176, 4.982718, 4.973215, 4.960507, 
    4.944603, 4.925617, 4.903484, 4.88278, 4.861875, 4.842131, 4.824929, 
    4.811468, 4.802634, 4.798907, 4.800348, 4.806618, 4.817043, 4.830686, 
    4.846407, 4.862938, 4.878937, 4.893082, 4.904164, 4.911223, 4.913716, 
    4.911637,
  // height(17,39, 0-49)
    4.8885, 4.884964, 4.884163, 4.885783, 4.889422, 4.894643, 4.901007, 
    4.908122, 4.915665, 4.923398, 4.931163, 4.938869, 4.946483, 4.95401, 
    4.961489, 4.963247, 4.971654, 4.976719, 4.979917, 4.981703, 4.982242, 
    4.984488, 4.984486, 4.982543, 4.978146, 4.970976, 4.960778, 4.947517, 
    4.931282, 4.912557, 4.891349, 4.872391, 4.853734, 4.836616, 4.822244, 
    4.811627, 4.805473, 4.804114, 4.807503, 4.815238, 4.826606, 4.840658, 
    4.856246, 4.87211, 4.886935, 4.899451, 4.908543, 4.913409, 4.913702, 
    4.909656,
  // height(17,40, 0-49)
    4.895968, 4.892166, 4.890924, 4.891946, 4.894863, 4.899263, 4.90474, 
    4.910928, 4.917522, 4.924296, 4.931087, 4.937795, 4.944351, 4.950702, 
    4.956784, 4.958094, 4.967124, 4.970757, 4.972659, 4.973285, 4.972751, 
    4.974173, 4.973469, 4.971002, 4.966048, 4.958385, 4.947799, 4.934374, 
    4.918255, 4.900277, 4.880496, 4.863629, 4.847486, 4.833153, 4.821659, 
    4.813825, 4.810189, 4.810955, 4.815989, 4.824837, 4.836764, 4.850812, 
    4.865849, 4.880637, 4.893913, 4.904496, 4.911415, 4.914057, 4.912313, 
    4.906664,
  // height(17,41, 0-49)
    4.902921, 4.898695, 4.89686, 4.897158, 4.899249, 4.902759, 4.907311, 
    4.91256, 4.918214, 4.924046, 4.929891, 4.935626, 4.941149, 4.946351, 
    4.951089, 4.952054, 4.96143, 4.963621, 4.964247, 4.963741, 4.962173, 
    4.962739, 4.96137, 4.958476, 4.95314, 4.945245, 4.934614, 4.921438, 
    4.905893, 4.88913, 4.871221, 4.856738, 4.843309, 4.831854, 4.823215, 
    4.818036, 4.816703, 4.819304, 4.825633, 4.835196, 4.847248, 4.860843, 
    4.874875, 4.888161, 4.899525, 4.907917, 4.912551, 4.913051, 4.909559, 
    4.9028,
  // height(17,42, 0-49)
    4.909159, 4.904336, 4.901761, 4.901208, 4.902383, 4.904947, 4.90855, 
    4.912868, 4.917612, 4.922549, 4.9275, 4.932313, 4.936859, 4.940983, 
    4.944482, 4.945125, 4.954541, 4.955351, 4.954765, 4.953189, 4.95065, 
    4.950379, 4.948419, 4.945224, 4.939711, 4.931865, 4.921547, 4.909028, 
    4.894497, 4.879364, 4.863691, 4.851813, 4.841222, 4.832664, 4.826799, 
    4.8241, 4.824811, 4.828923, 4.836165, 4.846019, 4.857746, 4.870423, 
    4.883003, 4.894386, 4.903529, 4.90956, 4.911921, 4.910494, 4.905684, 
    4.898421,
  // height(17,43, 0-49)
    4.914628, 4.909033, 4.905563, 4.904037, 4.904203, 4.905764, 4.908397, 
    4.91179, 4.915656, 4.919752, 4.923867, 4.927831, 4.931473, 4.934608, 
    4.936998, 4.937302, 4.946457, 4.946009, 4.944318, 4.94176, 4.938349, 
    4.937307, 4.934862, 4.93152, 4.926051, 4.91854, 4.908878, 4.897394, 
    4.884263, 4.871099, 4.857931, 4.848797, 4.84109, 4.835384, 4.832156, 
    4.83172, 4.834194, 4.839475, 4.847241, 4.856964, 4.867921, 4.879242, 
    4.889966, 4.899126, 4.905847, 4.909483, 4.909735, 4.906756, 4.901185, 
    4.894104,
  // height(17,44, 0-49)
    4.919461, 4.912925, 4.908408, 4.905779, 4.904836, 4.90532, 4.90694, 
    4.909394, 4.912395, 4.915678, 4.919009, 4.92218, 4.924991, 4.92723, 
    4.928645, 4.928577, 4.937214, 4.935669, 4.933005, 4.929586, 4.925431, 
    4.923725, 4.920937, 4.917611, 4.91241, 4.905505, 4.896807, 4.88668, 
    4.875265, 4.864319, 4.85382, 4.847488, 4.84264, 4.839678, 4.838911, 
    4.8405, 4.844442, 4.850554, 4.858476, 4.867672, 4.877462, 4.887057, 
    4.895621, 4.902356, 4.906611, 4.907991, 4.906475, 4.902468, 4.896797, 
    4.890616,
  // height(17,45, 0-49)
    4.924008, 4.916375, 4.910664, 4.906796, 4.904622, 4.903929, 4.904456, 
    4.905918, 4.908018, 4.910478, 4.913033, 4.91544, 4.91747, 4.918889, 
    4.919441, 4.918964, 4.926886, 4.924419, 4.920935, 4.916797, 4.912052, 
    4.909824, 4.906849, 4.903707, 4.898986, 4.892923, 4.885447, 4.876929, 
    4.86746, 4.858889, 4.851131, 4.847575, 4.845493, 4.84512, 4.846608, 
    4.849974, 4.855102, 4.861737, 4.869482, 4.877822, 4.886137, 4.893749, 
    4.899987, 4.904269, 4.906194, 4.90565, 4.902875, 4.898486, 4.893424, 
    4.888831,
  // height(17,46, 0-49)
    4.928825, 4.919962, 4.912918, 4.90767, 4.904126, 4.902122, 4.90143, 
    4.901784, 4.902892, 4.904456, 4.906185, 4.907807, 4.909061, 4.909698, 
    4.909465, 4.908536, 4.915604, 4.912388, 4.908238, 4.903537, 4.898368, 
    4.895784, 4.892784, 4.88998, 4.885921, 4.880892, 4.874827, 4.868092, 
    4.860718, 4.854588, 4.849548, 4.848677, 4.849215, 4.851243, 4.854764, 
    4.859663, 4.865725, 4.87262, 4.879941, 4.887194, 4.89385, 4.899375, 
    4.903301, 4.905291, 4.905223, 4.903256, 4.899861, 4.895799, 4.892039, 
    4.889628,
  // height(17,47, 0-49)
    4.934628, 4.924436, 4.915936, 4.909171, 4.904103, 4.900622, 4.898542, 
    4.897622, 4.897577, 4.898103, 4.89889, 4.899638, 4.900064, 4.899903, 
    4.898912, 4.897471, 4.903601, 4.899779, 4.895105, 4.889996, 4.884573, 
    4.881795, 4.878922, 4.876583, 4.873326, 4.869465, 4.864933, 4.860072, 
    4.85486, 4.851156, 4.848743, 4.850405, 4.853375, 4.857594, 4.862926, 
    4.869143, 4.875928, 4.882905, 4.889649, 4.895721, 4.900694, 4.904212, 
    4.906034, 4.906089, 4.904534, 4.901772, 4.898455, 4.895413, 4.893567, 
    4.893793,
  // height(17,48, 0-49)
    4.942206, 4.930628, 4.920584, 4.912177, 4.905432, 4.900293, 4.896624, 
    4.894217, 4.892807, 4.892093, 4.891754, 4.891472, 4.890954, 4.889923, 
    4.888144, 4.886106, 4.891249, 4.886915, 4.881835, 4.876449, 4.870919, 
    4.868098, 4.865475, 4.863686, 4.861314, 4.858688, 4.855734, 4.852766, 
    4.84971, 4.848352, 4.848417, 4.852421, 4.857611, 4.863803, 4.870745, 
    4.878098, 4.885471, 4.89244, 4.898585, 4.903532, 4.906981, 4.908762, 
    4.908873, 4.907512, 4.905091, 4.902219, 4.899659, 4.898243, 4.898774, 
    4.901918,
  // height(17,49, 0-49)
    4.959617, 4.946238, 4.934052, 4.923233, 4.913883, 4.906022, 4.89959, 
    4.894449, 4.890389, 4.887144, 4.884412, 4.881876, 4.879222, 4.876143, 
    4.872361, 4.869101, 4.880398, 4.874001, 4.866947, 4.860031, 4.853502, 
    4.852767, 4.852791, 4.85458, 4.855067, 4.854731, 4.853221, 4.850918, 
    4.847435, 4.846223, 4.846673, 4.853611, 4.861576, 4.870242, 4.879228, 
    4.888075, 4.896299, 4.903437, 4.909089, 4.912979, 4.914989, 4.915207, 
    4.913942, 4.911713, 4.909215, 4.907247, 4.906631, 4.908108, 4.91226, 
    4.919442,
  // height(18,0, 0-49)
    4.884809, 4.871144, 4.860725, 4.853534, 4.849423, 4.848121, 4.849251, 
    4.852354, 4.856926, 4.862458, 4.868456, 4.874484, 4.880164, 4.885192, 
    4.88933, 4.892411, 4.895638, 4.896484, 4.896322, 4.895182, 4.893073, 
    4.890365, 4.886718, 4.882278, 4.87701, 4.871042, 4.864499, 4.857598, 
    4.850573, 4.843819, 4.837571, 4.832456, 4.82845, 4.825788, 4.824625, 
    4.825011, 4.826875, 4.830015, 4.834108, 4.838731, 4.843399, 4.84762, 
    4.850959, 4.853108, 4.853957, 4.853652, 4.852622, 4.851551, 4.851324, 
    4.852911,
  // height(18,1, 0-49)
    4.884934, 4.871832, 4.862022, 4.855465, 4.85199, 4.851309, 4.853025, 
    4.856676, 4.861752, 4.867746, 4.874176, 4.880609, 4.886672, 4.892051, 
    4.896487, 4.899747, 4.904272, 4.905182, 4.905079, 4.903979, 4.901849, 
    4.899334, 4.895684, 4.891092, 4.885404, 4.878729, 4.871161, 4.862932, 
    4.854278, 4.845744, 4.837555, 4.830768, 4.825129, 4.820971, 4.818543, 
    4.817976, 4.819256, 4.822213, 4.826527, 4.831753, 4.837351, 4.842746, 
    4.847396, 4.850862, 4.852898, 4.853511, 4.853005, 4.851987, 4.851309, 
    4.851967,
  // height(18,2, 0-49)
    4.886409, 4.873914, 4.864717, 4.858756, 4.855839, 4.85566, 4.857812, 
    4.861832, 4.867219, 4.87348, 4.880151, 4.886819, 4.893123, 4.898752, 
    4.903427, 4.906798, 4.912543, 4.913613, 4.913682, 4.912762, 4.910775, 
    4.908639, 4.905188, 4.900646, 4.894743, 4.887562, 4.879149, 4.869736, 
    4.859549, 4.849249, 4.839058, 4.830468, 4.823002, 4.817106, 4.813138, 
    4.811329, 4.811743, 4.814265, 4.818604, 4.82431, 4.830813, 4.837478, 
    4.84367, 4.848833, 4.852573, 4.854734, 4.855453, 4.855189, 4.854686, 
    4.854899,
  // height(18,3, 0-49)
    4.888647, 4.876785, 4.868192, 4.862783, 4.86035, 4.860566, 4.863028, 
    4.867271, 4.872816, 4.879192, 4.885966, 4.892745, 4.899195, 4.905011, 
    4.909902, 4.913323, 4.920159, 4.921499, 4.921853, 4.921245, 4.919561, 
    4.917976, 4.914915, 4.910623, 4.904731, 4.897276, 4.888249, 4.877862, 
    4.866318, 4.854356, 4.842188, 4.831735, 4.822308, 4.814471, 4.808708, 
    4.805367, 4.804612, 4.806405, 4.810504, 4.816482, 4.823758, 4.831663, 
    4.839493, 4.846585, 4.852404, 4.856616, 4.859165, 4.860306, 4.860612, 
    4.860924,
  // height(18,4, 0-49)
    4.89114, 4.879928, 4.871926, 4.867028, 4.865009, 4.865537, 4.868205, 
    4.872565, 4.878159, 4.884547, 4.891326, 4.898142, 4.904681, 4.910653, 
    4.915773, 4.919184, 4.926921, 4.92865, 4.929398, 4.929215, 4.927966, 
    4.927078, 4.924573, 4.920717, 4.91506, 4.907583, 4.898214, 4.887125, 
    4.874485, 4.861058, 4.847029, 4.834742, 4.823296, 4.813377, 4.805604, 
    4.800458, 4.798227, 4.798971, 4.802519, 4.808488, 4.816317, 4.825317, 
    4.834739, 4.843832, 4.851933, 4.858536, 4.863369, 4.866457, 4.868152, 
    4.869117,
  // height(18,5, 0-49)
    4.893487, 4.882936, 4.875515, 4.871094, 4.869439, 4.870214, 4.873019, 
    4.877421, 4.882993, 4.889328, 4.89606, 4.90287, 4.909472, 4.915598, 
    4.920979, 4.924315, 4.932712, 4.934937, 4.936172, 4.936502, 4.935794, 
    4.935705, 4.933889, 4.930626, 4.925414, 4.918171, 4.908759, 4.897293, 
    4.883885, 4.869284, 4.853611, 4.839611, 4.826176, 4.814109, 4.80417, 
    4.796988, 4.792989, 4.792358, 4.795018, 4.800653, 4.808738, 4.818592, 
    4.829433, 4.840447, 4.85086, 4.860002, 4.867395, 4.872821, 4.876379, 
    4.878513,
  // height(18,6, 0-49)
    4.895404, 4.88553, 4.878681, 4.874718, 4.873394, 4.874374, 4.877271, 
    4.881673, 4.887185, 4.893434, 4.900091, 4.906876, 4.913533, 4.919827, 
    4.925513, 4.928716, 4.937472, 4.940289, 4.942079, 4.942984, 4.942886, 
    4.94365, 4.942612, 4.940061, 4.935476, 4.928711, 4.919563, 4.908076, 
    4.894294, 4.878877, 4.861876, 4.846375, 4.831077, 4.816886, 4.8047, 
    4.795306, 4.789286, 4.78697, 4.788401, 4.79335, 4.801349, 4.811738, 
    4.823725, 4.836451, 4.849043, 4.860695, 4.870737, 4.878716, 4.884475, 
    4.888203,
  // height(18,7, 0-49)
    4.896717, 4.887537, 4.881267, 4.877753, 4.876744, 4.877908, 4.880875, 
    4.885259, 4.890693, 4.896843, 4.903419, 4.910171, 4.916884, 4.92336, 
    4.929397, 4.932419, 4.941206, 4.944678, 4.947065, 4.948576, 4.949125, 
    4.950751, 4.950533, 4.948766, 4.944954, 4.938883, 4.930294, 4.919146, 
    4.905412, 4.889598, 4.871658, 4.854958, 4.838015, 4.821816, 4.807391, 
    4.795682, 4.787444, 4.783171, 4.783046, 4.786955, 4.794499, 4.80506, 
    4.81785, 4.831971, 4.846484, 4.860461, 4.873067, 4.88364, 4.891777, 
    4.897409,
  // height(18,8, 0-49)
    4.897334, 4.888876, 4.8832, 4.880144, 4.879449, 4.880795, 4.88383, 
    4.888193, 4.893551, 4.899602, 4.906095, 4.912813, 4.919581, 4.926244, 
    4.932665, 4.935491, 4.943973, 4.948122, 4.951126, 4.953247, 4.954448, 
    4.956897, 4.957495, 4.956541, 4.953597, 4.948393, 4.940624, 4.930164, 
    4.916898, 4.901135, 4.882703, 4.865164, 4.846878, 4.828883, 4.812316, 
    4.798274, 4.78769, 4.78124, 4.779273, 4.781801, 4.788523, 4.798871, 
    4.812071, 4.82721, 4.843288, 4.859285, 4.874232, 4.887288, 4.897826, 
    4.905539,
  // height(18,9, 0-49)
    4.897227, 4.889523, 4.884467, 4.881888, 4.881528, 4.883073, 4.886189, 
    4.890546, 4.895837, 4.901796, 4.908204, 4.914883, 4.921696, 4.928542, 
    4.935356, 4.938022, 4.945889, 4.950691, 4.9543, 4.957017, 4.958854, 
    4.962049, 4.963417, 4.963258, 4.96123, 4.957014, 4.950277, 4.940805, 
    4.928404, 4.913132, 4.894676, 4.876698, 4.85743, 4.837928, 4.819408, 
    4.803104, 4.790129, 4.78135, 4.777303, 4.778151, 4.783701, 4.793451, 
    4.806657, 4.822395, 4.839628, 4.857264, 4.874227, 4.889527, 4.902359, 
    4.912195,
  // height(18,10, 0-49)
    4.896404, 4.88949, 4.885093, 4.883026, 4.883033, 4.884808, 4.888037, 
    4.892411, 4.897654, 4.903532, 4.909855, 4.916485, 4.923323, 4.930325, 
    4.937502, 4.940127, 4.947123, 4.952506, 4.956683, 4.959964, 4.962405, 
    4.966238, 4.968298, 4.968881, 4.967768, 4.964606, 4.959049, 4.950807, 
    4.939605, 4.925227, 4.90721, 4.889191, 4.869336, 4.848673, 4.828465, 
    4.810056, 4.79473, 4.783552, 4.777253, 4.776168, 4.780232, 4.789024, 
    4.80184, 4.817754, 4.835709, 4.854557, 4.873146, 4.890373, 4.905285, 
    4.917168,
  // height(18,11, 0-49)
    4.894901, 4.888815, 4.885118, 4.88361, 4.884029, 4.886082, 4.889462, 
    4.893889, 4.899112, 4.904922, 4.911164, 4.917727, 4.924558, 4.931664, 
    4.939128, 4.941932, 4.947885, 4.95373, 4.958413, 4.962218, 4.965225, 
    4.969569, 4.972219, 4.97346, 4.973217, 4.971121, 4.966827, 4.95998, 
    4.950234, 4.937087, 4.91993, 4.90224, 4.882188, 4.860743, 4.839166, 
    4.818886, 4.801331, 4.787762, 4.779115, 4.775909, 4.778225, 4.785737, 
    4.797791, 4.813478, 4.831725, 4.851353, 4.87115, 4.889936, 4.906639, 
    4.920398,
  // height(18,12, 0-49)
    4.892765, 4.88754, 4.884587, 4.88369, 4.884581, 4.886966, 4.890554, 
    4.89508, 4.900316, 4.906077, 4.912237, 4.918715, 4.925493, 4.932621, 
    4.940238, 4.94356, 4.948406, 4.954556, 4.959667, 4.963951, 4.967489, 
    4.972205, 4.97533, 4.977124, 4.977676, 4.976608, 4.973598, 4.968228, 
    4.960105, 4.94844, 4.9325, 4.915447, 4.895557, 4.873702, 4.851109, 
    4.829243, 4.809653, 4.793781, 4.782765, 4.777319, 4.777685, 4.783647, 
    4.794613, 4.809704, 4.827843, 4.847833, 4.868425, 4.888381, 4.906549, 
    4.921947,
  // height(18,13, 0-49)
    4.890054, 4.885715, 4.88355, 4.883318, 4.884742, 4.887525, 4.891382, 
    4.89606, 4.901348, 4.907085, 4.913165, 4.919536, 4.926205, 4.93325, 
    4.940831, 4.945117, 4.948902, 4.955187, 4.960639, 4.96536, 4.969398, 
    4.97435, 4.977834, 4.980072, 4.981319, 4.981205, 4.979434, 4.975549, 
    4.969117, 4.959093, 4.944644, 4.928452, 4.909022, 4.887101, 4.86384, 
    4.840705, 4.81933, 4.801309, 4.787976, 4.780247, 4.778527, 4.782729, 
    4.792338, 4.806513, 4.824186, 4.844155, 4.865149, 4.885897, 4.905189, 
    4.921952,
  // height(18,14, 0-49)
    4.886841, 4.883399, 4.882051, 4.882535, 4.884551, 4.887797, 4.891985, 
    4.896872, 4.902257, 4.907996, 4.914003, 4.920245, 4.926744, 4.933584, 
    4.940909, 4.94667, 4.949551, 4.95581, 4.961526, 4.966652, 4.971175, 
    4.976239, 4.979972, 4.982547, 4.984378, 4.98511, 4.984487, 4.982019, 
    4.977257, 4.968933, 4.956161, 4.94096, 4.922206, 4.900504, 4.876897, 
    4.852814, 4.829932, 4.809971, 4.794442, 4.784451, 4.780582, 4.782882, 
    4.790926, 4.803923, 4.820827, 4.840441, 4.861489, 4.882676, 4.90276, 
    4.920603,
  // height(18,15, 0-49)
    4.883207, 4.880651, 4.880136, 4.881371, 4.884029, 4.887794, 4.892372, 
    4.897519, 4.903045, 4.908817, 4.914763, 4.920861, 4.927134, 4.93365, 
    4.940502, 4.948238, 4.950455, 4.956568, 4.962499, 4.96802, 4.973034, 
    4.978105, 4.982003, 4.984821, 4.987122, 4.988574, 4.988962, 4.987782, 
    4.984583, 4.977922, 4.966918, 4.952744, 4.934793, 4.913519, 4.889838, 
    4.865107, 4.84101, 4.819353, 4.801796, 4.789631, 4.783615, 4.783937, 
    4.790273, 4.801894, 4.817789, 4.836773, 4.857575, 4.878895, 4.899468, 
    4.918118,
  // height(18,16, 0-49)
    4.879242, 4.87754, 4.87785, 4.879844, 4.883172, 4.887492, 4.892501, 
    4.897952, 4.903658, 4.909498, 4.915406, 4.921362, 4.92738, 4.933488, 
    4.939705, 4.949776, 4.951613, 4.95754, 4.963687, 4.969635, 4.975175, 
    4.98018, 4.984186, 4.987179, 4.989842, 4.991875, 4.993103, 4.993021, 
    4.991203, 4.986084, 4.976843, 4.963641, 4.946527, 4.925811, 4.902266, 
    4.877148, 4.852115, 4.829021, 4.809649, 4.795449, 4.787349, 4.785682, 
    4.790234, 4.800347, 4.815056, 4.8332, 4.853517, 4.874714, 4.895517, 
    4.914725,
  // height(18,17, 0-49)
    4.875041, 4.874127, 4.875218, 4.87795, 4.881939, 4.886819, 4.892274, 
    4.898053, 4.903974, 4.909922, 4.915837, 4.921696, 4.927484, 4.933181, 
    4.938707, 4.951196, 4.952917, 4.958723, 4.965165, 4.971624, 4.977774, 
    4.982686, 4.986784, 4.989913, 4.992849, 4.995311, 4.997171, 4.997947, 
    4.997252, 4.993465, 4.9859, 4.973534, 4.95721, 4.937099, 4.913828, 
    4.888538, 4.862826, 4.838557, 4.817604, 4.801552, 4.791484, 4.787878, 
    4.790633, 4.799174, 4.812584, 4.829738, 4.849395, 4.870271, 4.891096, 
    4.910655,
  // height(18,18, 0-49)
    4.870688, 4.87046, 4.872247, 4.875643, 4.880235, 4.885635, 4.891515, 
    4.897624, 4.90379, 4.909906, 4.91592, 4.921796, 4.927487, 4.932893, 
    4.937829, 4.952391, 4.954152, 4.960028, 4.966936, 4.974069, 4.980973, 
    4.985815, 4.99005, 4.993322, 4.99646, 4.999198, 5.001451, 5.002779, 
    5.002877, 5.000129, 4.994055, 4.982319, 4.966665, 4.947137, 4.924218, 
    4.898921, 4.872756, 4.847573, 4.825289, 4.807601, 4.795727, 4.790283, 
    4.791286, 4.798248, 4.810311, 4.826389, 4.84527, 4.865687, 4.886379, 
    4.906126,
  // height(18,19, 0-49)
    4.86625, 4.86655, 4.868883, 4.872808, 4.877879, 4.883698, 4.889936, 
    4.896357, 4.902807, 4.909202, 4.915492, 4.921624, 4.927492, 4.932897, 
    4.937518, 4.953274, 4.955041, 4.961284, 4.968928, 4.976991, 4.984876, 
    4.989754, 4.994244, 4.997727, 5.001033, 5.003887, 5.006248, 5.007756, 
    5.008227, 5.006122, 5.001248, 4.98988, 4.974717, 4.955695, 4.933158, 
    4.907983, 4.881572, 4.855722, 4.832371, 4.813286, 4.799805, 4.792671, 
    4.792016, 4.797443, 4.808165, 4.823141, 4.841189, 4.861065, 4.881521, 
    4.901341,
  // height(18,20, 0-49)
    4.862615, 4.864183, 4.867981, 4.873559, 4.880429, 4.888097, 4.896105, 
    4.904039, 4.91155, 4.918352, 4.924236, 4.929071, 4.932817, 4.935514, 
    4.937287, 0, 4.967083, 4.970193, 4.974487, 4.979447, 4.9848, 4.986744, 
    4.989418, 4.992031, 4.995424, 4.999174, 5.003032, 5.006403, 5.008925, 
    5.008933, 5.006418, 4.996209, 4.982046, 4.963815, 4.941799, 4.916811, 
    4.8902, 4.86374, 4.83939, 4.818989, 4.803974, 4.79521, 4.792936, 
    4.796848, 4.806228, 4.820079, 4.837255, 4.856534, 4.87668, 4.896485,
  // height(18,21, 0-49)
    4.858526, 4.860593, 4.864909, 4.870983, 4.878288, 4.886311, 4.89458, 
    4.902694, 4.910328, 4.917231, 4.923228, 4.928211, 4.932137, 4.935033, 
    4.936998, 0, 4.96749, 4.971151, 4.976059, 4.981626, 4.987492, 4.988534, 
    4.990527, 4.992525, 4.995533, 4.999171, 5.003212, 5.007048, 5.010316, 
    5.011328, 5.010325, 5.000771, 4.987464, 4.970185, 4.949078, 4.924807, 
    4.898589, 4.872103, 4.847268, 4.82596, 4.809701, 4.799472, 4.795639, 
    4.798006, 4.805933, 4.818489, 4.834568, 4.852976, 4.872499, 4.891943,
  // height(18,22, 0-49)
    4.854605, 4.857058, 4.861805, 4.868328, 4.876069, 4.884493, 4.893115, 
    4.901526, 4.909408, 4.916522, 4.922707, 4.927864, 4.931949, 4.93498, 
    4.937038, 0, 4.968196, 4.972306, 4.977769, 4.98394, 4.990365, 4.990649, 
    4.992125, 4.993677, 4.996429, 5.000011, 5.004191, 5.008338, 5.01208, 
    5.013722, 5.013745, 5.004387, 4.991473, 4.974729, 4.954206, 4.930459, 
    4.904589, 4.878174, 4.853073, 4.831153, 4.813982, 4.802622, 4.797538, 
    4.798625, 4.805327, 4.816769, 4.831888, 4.849522, 4.86848, 4.887581,
  // height(18,23, 0-49)
    4.850917, 4.853661, 4.858761, 4.865675, 4.873829, 4.882668, 4.891686, 
    4.900468, 4.908682, 4.916094, 4.922538, 4.927917, 4.932185, 4.935344, 
    4.93747, 0, 4.969583, 4.973991, 4.979832, 4.98642, 4.993236, 4.992826, 
    4.993824, 4.99496, 4.99745, 5.000928, 5.005152, 5.009469, 5.013495, 
    5.015525, 5.016229, 5.006853, 4.994095, 4.977653, 4.95752, 4.934175, 
    4.908624, 4.882356, 4.857164, 4.834885, 4.817104, 4.804931, 4.798903, 
    4.798989, 4.804698, 4.81521, 4.8295, 4.846437, 4.864852, 4.883585,
  // height(18,24, 0-49)
    4.847519, 4.850479, 4.85586, 4.863112, 4.871647, 4.880895, 4.890332, 
    4.899526, 4.908134, 4.915905, 4.92267, 4.928324, 4.932813, 4.936135, 
    4.938357, 0, 4.971826, 4.976392, 4.982431, 4.989242, 4.996271, 4.995375, 
    4.996037, 4.996878, 4.999168, 5.002536, 5.006739, 5.011106, 5.015255, 
    5.017463, 5.018531, 5.009044, 4.996279, 4.979924, 4.959941, 4.936765, 
    4.911347, 4.885115, 4.859817, 4.837259, 4.819028, 4.806264, 4.799543, 
    4.798884, 4.803843, 4.813639, 4.827281, 4.843661, 4.86163, 4.880041,
  // height(18,25, 0-49)
    4.84447, 4.847589, 4.853196, 4.860741, 4.869628, 4.879272, 4.889136, 
    4.898769, 4.907809, 4.915988, 4.923122, 4.929097, 4.933853, 4.937385, 
    4.939763, 0, 4.974479, 4.979081, 4.985147, 4.991983, 4.999034, 4.997939, 
    4.99846, 4.999179, 5.001375, 5.00467, 5.008821, 5.013151, 5.017279, 
    5.019472, 5.020578, 5.010951, 4.998077, 4.981641, 4.961603, 4.938382, 
    4.91291, 4.88659, 4.861147, 4.838369, 4.819839, 4.806698, 4.799538, 
    4.7984, 4.802862, 4.81217, 4.825348, 4.841312, 4.858924, 4.877048,
  // height(18,26, 0-49)
    4.841846, 4.845082, 4.850876, 4.858679, 4.867893, 4.877924, 4.888223, 
    4.898314, 4.907815, 4.916437, 4.923976, 4.930305, 4.935359, 4.939139, 
    4.941726, 0, 4.977385, 4.981901, 4.98783, 4.994493, 5.001371, 5.000391, 
    5.000994, 5.001788, 5.004019, 5.007303, 5.01139, 5.015614, 5.019589, 
    5.021584, 5.022406, 5.012643, 4.999584, 4.982924, 4.962636, 4.939158, 
    4.913439, 4.886895, 4.861254, 4.838302, 4.819606, 4.806296, 4.798949, 
    4.797599, 4.801824, 4.810872, 4.823782, 4.839473, 4.856821, 4.874699,
  // height(18,27, 0-49)
    4.839744, 4.843068, 4.84902, 4.857059, 4.866587, 4.877005, 4.887747, 
    4.898317, 4.908307, 4.917399, 4.925366, 4.932062, 4.937419, 4.941448, 
    4.944248, 0, 4.980576, 4.984866, 4.990472, 4.996755, 5.003257, 5.002659, 
    5.003529, 5.004568, 5.006943, 5.01026, 5.014267, 5.018305, 5.021995, 
    5.023608, 5.023826, 5.013915, 5.000586, 4.983556, 4.962839, 4.938921, 
    4.912803, 4.885948, 4.860112, 4.837081, 4.818402, 4.805168, 4.797915, 
    4.796639, 4.800896, 4.809918, 4.822744, 4.838297, 4.855458, 4.873108,
  // height(18,28, 0-49)
    4.838279, 4.841671, 4.847761, 4.856022, 4.86586, 4.876674, 4.887884, 
    4.898968, 4.909482, 4.919071, 4.927473, 4.934519, 4.940135, 4.94435, 
    4.94729, 0, 4.984393, 4.988278, 4.993347, 4.999027, 5.004954, 5.004905, 
    5.006158, 5.007552, 5.010141, 5.013506, 5.017393, 5.021155, 5.024417, 
    5.025462, 5.024777, 5.014656, 5.000932, 4.983361, 4.962024, 4.937493, 
    4.910855, 4.883649, 4.857671, 4.834711, 4.816276, 4.803395, 4.796536, 
    4.795633, 4.800196, 4.80943, 4.82236, 4.837905, 4.854949, 4.872379,
  // height(18,29, 0-49)
    4.837578, 4.841016, 4.847223, 4.855696, 4.865859, 4.8771, 4.888828, 
    4.900484, 4.911574, 4.921689, 4.930514, 4.937848, 4.943614, 4.94786, 
    4.950751, 0, 4.988549, 4.991818, 4.996123, 5.000973, 5.006124, 5.006631, 
    5.00827, 5.010037, 5.012847, 5.016247, 5.019962, 5.023355, 5.02604, 
    5.026312, 5.024417, 5.013925, 4.999619, 4.981328, 4.959243, 4.93405, 
    4.906947, 4.879553, 4.853701, 4.831154, 4.813352, 4.801226, 4.795144, 
    4.794957, 4.800112, 4.80978, 4.822963, 4.83858, 4.855508, 4.872646,
  // height(18,30, 0-49)
    4.837201, 4.839952, 4.84534, 4.852841, 4.861905, 4.872, 4.882656, 
    4.893489, 4.904216, 4.914642, 4.924639, 4.934104, 4.942914, 4.950874, 
    4.957664, 4.980512, 4.978384, 4.985451, 4.993881, 5.002621, 5.011064, 
    5.015289, 5.019503, 5.022801, 5.026014, 5.028763, 5.03095, 5.032186, 
    5.032328, 5.02988, 5.02498, 5.012665, 4.996644, 4.97683, 4.95351, 
    4.927465, 4.899968, 4.872666, 4.847361, 4.825732, 4.809091, 4.798231, 
    4.793395, 4.794331, 4.800419, 4.81079, 4.824425, 4.840233, 4.8571, 
    4.873925,
  // height(18,31, 0-49)
    4.838711, 4.841673, 4.847275, 4.855004, 4.864307, 4.874646, 4.885531, 
    4.896559, 4.907419, 4.917896, 4.927857, 4.937228, 4.945951, 4.953948, 
    4.961065, 4.980995, 4.980417, 4.987096, 4.994756, 5.002519, 5.00993, 
    5.014159, 5.018117, 5.021186, 5.024208, 5.026828, 5.028913, 5.029993, 
    5.029801, 5.02675, 5.020671, 5.008065, 4.991631, 4.971384, 4.94774, 
    4.9216, 4.89433, 4.86762, 4.843251, 4.822825, 4.807539, 4.798059, 
    4.794508, 4.796546, 4.803485, 4.814416, 4.828295, 4.844025, 4.860487, 
    4.876597,
  // height(18,32, 0-49)
    4.841342, 4.844412, 4.850084, 4.857855, 4.867183, 4.877531, 4.888418, 
    4.899436, 4.910273, 4.920713, 4.930632, 4.93998, 4.948754, 4.956964, 
    4.964594, 4.980965, 4.981505, 4.988069, 4.995195, 5.002202, 5.00878, 
    5.013144, 5.016983, 5.019907, 5.02272, 5.025066, 5.026776, 5.02734, 
    5.026409, 5.022374, 5.014822, 5.001704, 4.984722, 4.964009, 4.940114, 
    4.914057, 4.88728, 4.861488, 4.838411, 4.819547, 4.80595, 4.798151, 
    4.796151, 4.799515, 4.807491, 4.819123, 4.833344, 4.849035, 4.865076, 
    4.880392,
  // height(18,33, 0-49)
    4.845201, 4.848296, 4.853919, 4.861576, 4.870737, 4.880888, 4.891561, 
    4.902365, 4.912999, 4.923262, 4.933043, 4.942318, 4.951126, 4.959552, 
    4.967697, 4.980441, 4.981912, 4.988523, 4.995258, 5.001646, 5.007523, 
    5.012081, 5.015876, 5.018697, 5.021259, 5.023195, 5.024305, 5.02406, 
    5.022061, 5.016749, 5.007536, 4.993733, 4.976113, 4.954939, 4.930896, 
    4.905118, 4.879101, 4.85454, 4.833084, 4.816096, 4.804484, 4.798627, 
    4.798405, 4.803288, 4.812459, 4.824915, 4.839553, 4.855231, 4.870821, 
    4.885258,
  // height(18,34, 0-49)
    4.850313, 4.853356, 4.858818, 4.866215, 4.875041, 4.884804, 4.895066, 
    4.905462, 4.915716, 4.925641, 4.935148, 4.944232, 4.952967, 4.961494, 
    4.970001, 4.979457, 4.981847, 4.98854, 4.994935, 5.000776, 5.006025, 
    5.010772, 5.014541, 5.01726, 5.019513, 5.020917, 5.02124, 5.019953, 
    5.016633, 5.00984, 4.998881, 4.98429, 4.966008, 4.944437, 4.920403, 
    4.895131, 4.870153, 4.847122, 4.82758, 4.812739, 4.803346, 4.799632, 
    4.801355, 4.8079, 4.818378, 4.831736, 4.846831, 4.862496, 4.877587, 
    4.891049,
  // height(18,35, 0-49)
    4.85662, 4.859527, 4.864711, 4.871711, 4.880044, 4.889249, 4.898926, 
    4.908741, 4.918445, 4.927876, 4.936965, 4.94572, 4.954232, 4.962675, 
    4.971297, 4.978046, 4.981433, 4.988136, 4.99417, 4.999484, 5.004143, 
    5.009024, 5.012743, 5.015333, 5.017207, 5.017971, 5.017355, 5.014852, 
    5.01003, 5.001642, 4.988949, 4.973538, 4.954648, 4.932821, 4.909005, 
    4.884502, 4.860847, 4.839624, 4.822244, 4.809759, 4.80275, 4.801305, 
    4.805072, 4.813345, 4.825176, 4.839457, 4.855005, 4.870616, 4.885136, 
    4.89752,
  // height(18,36, 0-49)
    4.863973, 4.866647, 4.871443, 4.877914, 4.885613, 4.894113, 4.903052, 
    4.912133, 4.921141, 4.929941, 4.938475, 4.946762, 4.954895, 4.963057, 
    4.971507, 4.97621, 4.980695, 4.987263, 4.992869, 4.997642, 5.001723, 
    5.006649, 5.010259, 5.012672, 5.014094, 5.014126, 5.01246, 5.008624, 
    5.0022, 4.992191, 4.977875, 4.961699, 4.942339, 4.920467, 4.897135, 
    4.87369, 4.85164, 4.83247, 4.817447, 4.807454, 4.802914, 4.80378, 
    4.809597, 4.819584, 4.832732, 4.847884, 4.863813, 4.879286, 4.893135, 
    4.904335,
  // height(18,37, 0-49)
    4.872146, 4.874485, 4.878777, 4.884603, 4.891544, 4.899216, 4.907293, 
    4.91552, 4.923715, 4.931767, 4.939631, 4.947328, 4.954942, 4.962633, 
    4.970646, 4.973928, 4.979574, 4.985822, 4.990914, 4.995116, 4.99861, 
    5.003463, 5.006887, 5.00906, 5.009962, 5.009189, 5.006405, 5.001185, 
    4.993144, 4.981586, 4.965855, 4.949062, 4.929453, 4.907815, 4.885276, 
    4.863191, 4.843011, 4.8261, 4.813562, 4.806119, 4.804044, 4.807168, 
    4.814948, 4.826537, 4.840876, 4.856761, 4.872931, 4.888124, 4.901169, 
    4.911073,
  // height(18,38, 0-49)
    4.880842, 4.882741, 4.886423, 4.891498, 4.897586, 4.904336, 4.911465, 
    4.918751, 4.926048, 4.933264, 4.940367, 4.947376, 4.954354, 4.961426, 
    4.968778, 4.971156, 4.977955, 4.983696, 4.988179, 4.991767, 4.994656, 
    4.999306, 5.002451, 5.004314, 5.004631, 5.003013, 4.999096, 4.992517, 
    4.982934, 4.969998, 4.953146, 4.935975, 4.916419, 4.895351, 4.873941, 
    4.853517, 4.83544, 4.820933, 4.810941, 4.806021, 4.806313, 4.811546, 
    4.821102, 4.834083, 4.849388, 4.86578, 4.881971, 4.896688, 4.908768, 
    4.917272,
  // height(18,39, 0-49)
    4.889717, 4.891066, 4.894044, 4.898291, 4.903454, 4.909225, 4.915352, 
    4.921652, 4.927999, 4.934326, 4.940608, 4.946858, 4.953117, 4.959458, 
    4.965996, 4.96784, 4.975702, 4.980766, 4.984552, 4.987484, 4.989732, 
    4.99404, 4.996809, 4.998293, 4.997983, 4.995514, 4.990504, 4.982667, 
    4.971714, 4.957668, 4.940073, 4.922842, 4.903699, 4.883575, 4.863635, 
    4.84515, 4.829363, 4.817347, 4.809879, 4.807374, 4.809848, 4.816947, 
    4.827996, 4.842059, 4.858009, 4.874594, 4.890515, 4.904504, 4.915439, 
    4.922453,
  // height(18,40, 0-49)
    4.8984, 4.899097, 4.90129, 4.904646, 4.908849, 4.913617, 4.91873, 
    4.924032, 4.929419, 4.934838, 4.940274, 4.945725, 4.951211, 4.956755, 
    4.96239, 4.963936, 4.972683, 4.976931, 4.979949, 4.982178, 4.983747, 
    4.987577, 4.989875, 4.990921, 4.989964, 4.98668, 4.98068, 4.971765, 
    4.959704, 4.944898, 4.927004, 4.910091, 4.891764, 4.872965, 4.854824, 
    4.838517, 4.825151, 4.815638, 4.810602, 4.81032, 4.814709, 4.823346, 
    4.835516, 4.850266, 4.866456, 4.882841, 4.898137, 4.911113, 4.920713, 
    4.926178,
  // height(18,41, 0-49)
    4.906529, 4.906476, 4.907814, 4.910242, 4.91347, 4.917244, 4.921369, 
    4.925701, 4.930154, 4.934687, 4.939281, 4.94393, 4.948625, 4.953344, 
    4.958044, 4.959407, 4.968792, 4.97213, 4.974324, 4.975806, 4.976653, 
    4.979882, 4.981626, 4.98219, 4.980597, 4.976579, 4.969752, 4.960011, 
    4.947186, 4.932035, 4.914319, 4.898144, 4.881041, 4.863939, 4.847887, 
    4.833943, 4.823065, 4.816005, 4.813236, 4.814918, 4.820882, 4.830656, 
    4.843504, 4.858468, 4.874428, 4.890163, 4.904439, 4.916101, 4.924196, 
    4.928107,
  // height(18,42, 0-49)
    4.913782, 4.912883, 4.913308, 4.914782, 4.917043, 4.919858, 4.923043, 
    4.926467, 4.93005, 4.933751, 4.937549, 4.941423, 4.945343, 4.949245, 
    4.953024, 4.954234, 4.963964, 4.96634, 4.967675, 4.96837, 4.968452, 
    4.970979, 4.972106, 4.972164, 4.969982, 4.965353, 4.957918, 4.947659, 
    4.934467, 4.919428, 4.902383, 4.887368, 4.871888, 4.856811, 4.843086, 
    4.831631, 4.823244, 4.818518, 4.817794, 4.821123, 4.82827, 4.83873, 
    4.851759, 4.866421, 4.881636, 4.896245, 4.9091, 4.919161, 4.925624, 
    4.928048,
  // height(18,43, 0-49)
    4.919908, 4.918075, 4.917529, 4.918031, 4.919343, 4.921244, 4.923561, 
    4.926164, 4.928969, 4.931925, 4.934999, 4.938159, 4.941349, 4.944471, 
    4.947376, 4.948405, 4.958177, 4.959578, 4.960035, 4.959912, 4.959199, 
    4.960948, 4.961421, 4.960978, 4.958283, 4.953208, 4.945422, 4.934996, 
    4.921866, 4.907401, 4.8915, 4.878047, 4.864542, 4.851766, 4.840542, 
    4.831635, 4.82568, 4.823121, 4.824172, 4.828796, 4.8367, 4.847362, 
    4.860054, 4.873881, 4.887831, 4.900847, 4.911908, 4.920138, 4.924921, 
    4.926015,
  // height(18,44, 0-49)
    4.924776, 4.921913, 4.92034, 4.91985, 4.920226, 4.921264, 4.92279, 
    4.924667, 4.926798, 4.929115, 4.931567, 4.934095, 4.936621, 4.939024, 
    4.941122, 4.941914, 4.951438, 4.951888, 4.951467, 4.95051, 4.94899, 
    4.94992, 4.94973, 4.948813, 4.945714, 4.940386, 4.932531, 4.9223, 
    4.909667, 4.896218, 4.881884, 4.870344, 4.859107, 4.848838, 4.840219, 
    4.833856, 4.830224, 4.829626, 4.832157, 4.837701, 4.845929, 4.856311, 
    4.868156, 4.880635, 4.89284, 4.903851, 4.912822, 4.91908, 4.922236, 
    4.922259,
  // height(18,45, 0-49)
    4.928407, 4.924418, 4.921751, 4.920234, 4.919677, 4.919885, 4.920683, 
    4.921923, 4.923484, 4.925271, 4.927204, 4.929194, 4.931141, 4.932897, 
    4.934264, 4.934757, 4.943786, 4.943328, 4.942047, 4.94026, 4.937941, 
    4.93805, 4.937223, 4.935887, 4.932515, 4.927137, 4.9195, 4.909817, 
    4.898086, 4.886047, 4.873634, 4.864293, 4.855537, 4.847908, 4.841933, 
    4.838057, 4.836599, 4.837729, 4.841436, 4.847537, 4.855672, 4.865327, 
    4.875862, 4.886545, 4.896604, 4.9053, 4.912002, 4.916276, 4.917975, 
    4.917284,
  // height(18,46, 0-49)
    4.931002, 4.925789, 4.921949, 4.919353, 4.917837, 4.917222, 4.917328, 
    4.917989, 4.919061, 4.920411, 4.921917, 4.92346, 4.924904, 4.926087, 
    4.926797, 4.926932, 4.935273, 4.933967, 4.931861, 4.929269, 4.926188, 
    4.925509, 4.924102, 4.922422, 4.918921, 4.9137, 4.906552, 4.897737, 
    4.887263, 4.876956, 4.866735, 4.859797, 4.853657, 4.848723, 4.845367, 
    4.843875, 4.844419, 4.84704, 4.851633, 4.857956, 4.865634, 4.87418, 
    4.883031, 4.891579, 4.899223, 4.905437, 4.90984, 4.912262, 4.912797, 
    4.911825,
  // height(18,47, 0-49)
    4.932955, 4.926421, 4.921322, 4.91757, 4.91504, 4.913567, 4.912973, 
    4.913074, 4.91369, 4.914652, 4.915792, 4.916949, 4.917954, 4.91862, 
    4.918736, 4.91845, 4.925973, 4.923887, 4.921003, 4.917657, 4.913873, 
    4.912481, 4.910572, 4.908642, 4.905159, 4.900286, 4.893863, 4.88618, 
    4.877249, 4.868914, 4.861065, 4.856644, 4.853178, 4.850926, 4.850114, 
    4.850874, 4.853234, 4.85712, 4.862342, 4.86861, 4.875546, 4.88271, 
    4.88963, 4.895852, 4.900975, 4.904717, 4.906961, 4.907805, 4.907571, 
    4.906791,
  // height(18,48, 0-49)
    4.934845, 4.9269, 4.920446, 4.915445, 4.911812, 4.909406, 4.908049, 
    4.907547, 4.907685, 4.908252, 4.909031, 4.909818, 4.910404, 4.910583, 
    4.91014, 4.909373, 4.916004, 4.9132, 4.909599, 4.905562, 4.90116, 
    4.899149, 4.896842, 4.894763, 4.891435, 4.887076, 4.881566, 4.875215, 
    4.868028, 4.861816, 4.856431, 4.854557, 4.85374, 4.854105, 4.855721, 
    4.858578, 4.862577, 4.867533, 4.873183, 4.879201, 4.885219, 4.890858, 
    4.895762, 4.899647, 4.902333, 4.903794, 4.904185, 4.903849, 4.903304, 
    4.90318,
  // height(18,49, 0-49)
    4.943079, 4.933022, 4.92444, 4.917368, 4.911783, 4.907586, 4.904629, 
    4.902708, 4.901586, 4.901, 4.900681, 4.900353, 4.899747, 4.898587, 
    4.896599, 4.894702, 4.907625, 4.902482, 4.896469, 4.890329, 4.884231, 
    4.883526, 4.882961, 4.883486, 4.882074, 4.87913, 4.874318, 4.868094, 
    4.860242, 4.854196, 4.849467, 4.851037, 4.85378, 4.857646, 4.86253, 
    4.868235, 4.874485, 4.880953, 4.887276, 4.893087, 4.898046, 4.901875, 
    4.904406, 4.905601, 4.905601, 4.904716, 4.90344, 4.902396, 4.902278, 
    4.903772,
  // height(19,0, 0-49)
    4.863467, 4.857262, 4.854007, 4.853439, 4.855211, 4.858918, 4.86413, 
    4.870421, 4.877393, 4.884692, 4.892019, 4.899126, 4.905809, 4.911901, 
    4.917256, 4.921696, 4.926414, 4.929109, 4.930936, 4.931877, 4.931879, 
    4.93122, 4.92947, 4.92665, 4.922586, 4.917221, 4.910484, 4.902398, 
    4.893026, 4.882643, 4.871445, 4.860118, 4.848811, 4.838039, 4.828342, 
    4.820229, 4.814119, 4.8103, 4.808887, 4.80981, 4.812818, 4.817494, 
    4.823306, 4.829645, 4.835906, 4.841548, 4.846171, 4.849586, 4.85186, 
    4.853332,
  // height(19,1, 0-49)
    4.865608, 4.859947, 4.857208, 4.857111, 4.8593, 4.863361, 4.868865, 
    4.875392, 4.882556, 4.890017, 4.897492, 4.904748, 4.911586, 4.917842, 
    4.923354, 4.927824, 4.933651, 4.936447, 4.938407, 4.939521, 4.939701, 
    4.939492, 4.938069, 4.935489, 4.931462, 4.925898, 4.918675, 4.909807, 
    4.899339, 4.887649, 4.874897, 4.862156, 4.849326, 4.837008, 4.825834, 
    4.816401, 4.809213, 4.804626, 4.802801, 4.803697, 4.807059, 4.812455, 
    4.8193, 4.826921, 4.834619, 4.841738, 4.847753, 4.85234, 4.855436, 
    4.857277,
  // height(19,2, 0-49)
    4.868079, 4.86294, 4.86067, 4.86098, 4.863502, 4.867823, 4.873523, 
    4.880189, 4.887453, 4.894991, 4.90254, 4.909874, 4.91681, 4.923179, 
    4.928813, 4.933246, 4.940066, 4.942986, 4.945104, 4.946426, 4.946843, 
    4.947165, 4.946175, 4.943969, 4.940157, 4.934615, 4.927167, 4.917808, 
    4.90655, 4.893838, 4.879786, 4.865834, 4.851622, 4.837819, 4.825143, 
    4.814283, 4.805833, 4.800229, 4.7977, 4.798252, 4.801656, 4.807476, 
    4.815114, 4.823852, 4.832918, 4.841565, 4.849153, 4.855217, 4.859553, 
    4.862253,
  // height(19,3, 0-49)
    4.870552, 4.86591, 4.864064, 4.864718, 4.867503, 4.872014, 4.877833, 
    4.884569, 4.891868, 4.899426, 4.906993, 4.914361, 4.921353, 4.927806, 
    4.93355, 4.937875, 4.945512, 4.948591, 4.950888, 4.952444, 4.953139, 
    4.954044, 4.953572, 4.95185, 4.948418, 4.943113, 4.935712, 4.926178, 
    4.914483, 4.901093, 4.886057, 4.871165, 4.855776, 4.840611, 4.826462, 
    4.814105, 4.804229, 4.797366, 4.793829, 4.793693, 4.796775, 4.802673, 
    4.810785, 4.820376, 4.830633, 4.840738, 4.84995, 4.857678, 4.863564, 
    4.867543,
  // height(19,4, 0-49)
    4.872817, 4.868643, 4.867184, 4.868135, 4.871129, 4.875768, 4.881651, 
    4.888405, 4.895691, 4.903227, 4.910775, 4.918141, 4.92516, 4.931677, 
    4.937528, 4.941673, 4.949905, 4.953179, 4.955673, 4.957477, 4.958472, 
    4.959987, 4.960082, 4.958926, 4.956011, 4.951143, 4.944056, 4.934675, 
    4.922916, 4.909231, 4.893579, 4.878071, 4.861773, 4.845433, 4.829899, 
    4.816028, 4.804605, 4.796266, 4.79143, 4.790257, 4.792642, 4.798227, 
    4.806442, 4.816557, 4.827739, 4.839124, 4.849892, 4.859341, 4.866971, 
    4.872547,
  // height(19,5, 0-49)
    4.874774, 4.871048, 4.869942, 4.871148, 4.874307, 4.879029, 4.884934, 
    4.891664, 4.898901, 4.906378, 4.913873, 4.921207, 4.928225, 4.93479, 
    4.940752, 4.944649, 4.953211, 4.956712, 4.959419, 4.961472, 4.962777, 
    4.964893, 4.965576, 4.96503, 4.962738, 4.958478, 4.951951, 4.943034, 
    4.931594, 4.918012, 4.902144, 4.886379, 4.869491, 4.852226, 4.835463, 
    4.820125, 4.807089, 4.797104, 4.790708, 4.788169, 4.789482, 4.79436, 
    4.802285, 4.812552, 4.824332, 4.836738, 4.848891, 4.860003, 4.869445, 
    4.876825,
  // height(19,6, 0-49)
    4.876401, 4.873109, 4.872334, 4.873767, 4.877055, 4.881827, 4.887718, 
    4.894387, 4.901539, 4.90892, 4.916327, 4.923593, 4.930583, 4.937176, 
    4.943255, 4.946844, 4.955447, 4.959205, 4.962132, 4.964428, 4.966038, 
    4.968722, 4.969982, 4.970057, 4.968456, 4.964935, 4.959171, 4.951004, 
    4.94024, 4.92715, 4.911473, 4.895832, 4.878706, 4.860817, 4.843043, 
    4.826352, 4.811706, 4.799966, 4.7918, 4.78761, 4.787505, 4.791297, 
    4.798542, 4.808578, 4.820599, 4.833713, 4.847009, 4.85963, 4.870845, 
    4.880115,
  // height(19,7, 0-49)
    4.877742, 4.87488, 4.87442, 4.876059, 4.879453, 4.884243, 4.890086, 
    4.896661, 4.903688, 4.910936, 4.918213, 4.925372, 4.932297, 4.938896, 
    4.945095, 4.948344, 4.956688, 4.960714, 4.963864, 4.966398, 4.968299, 
    4.971492, 4.973291, 4.973963, 4.973082, 4.970386, 4.965547, 4.958364, 
    4.94859, 4.936349, 4.921254, 4.906102, 4.889108, 4.870925, 4.852411, 
    4.83455, 4.818367, 4.804838, 4.79476, 4.78869, 4.78687, 4.789238, 
    4.795435, 4.80487, 4.816771, 4.830261, 4.844414, 4.858326, 4.871181, 
    4.882321,
  // height(19,8, 0-49)
    4.878867, 4.876438, 4.876289, 4.878121, 4.881602, 4.886387, 4.892151, 
    4.898596, 4.90546, 4.912529, 4.919632, 4.926641, 4.93346, 4.940037, 
    4.946343, 4.94926, 4.957064, 4.961346, 4.964719, 4.967476, 4.969651, 
    4.973279, 4.975556, 4.976775, 4.976603, 4.974774, 4.970967, 4.964946, 
    4.956418, 4.94533, 4.931167, 4.916834, 4.900319, 4.88219, 4.863243, 
    4.844447, 4.826875, 4.811594, 4.799544, 4.791435, 4.787673, 4.788329, 
    4.793161, 4.801657, 4.813101, 4.826638, 4.841345, 4.856289, 4.87059, 
    4.883487,
  // height(19,9, 0-49)
    4.879853, 4.877869, 4.878036, 4.880059, 4.883614, 4.888375, 4.894034, 
    4.900314, 4.906975, 4.913821, 4.920701, 4.927508, 4.934181, 4.940696, 
    4.94708, 4.94973, 4.956745, 4.961252, 4.964836, 4.967809, 4.970237, 
    4.974212, 4.976891, 4.978584, 4.979081, 4.978118, 4.975397, 4.970651, 
    4.963554, 4.953855, 4.940918, 4.927673, 4.911951, 4.894206, 4.875144, 
    4.855691, 4.836935, 4.820017, 4.80601, 4.795788, 4.789926, 4.788655, 
    4.791863, 4.799135, 4.809819, 4.823099, 4.838062, 4.853761, 4.86927, 
    4.883741,
  // height(19,10, 0-49)
    4.880766, 4.879248, 4.879743, 4.881961, 4.885587, 4.890312, 4.895844, 
    4.901929, 4.90835, 4.91493, 4.921543, 4.928103, 4.934577, 4.940979, 
    4.947385, 4.949909, 4.955944, 4.960614, 4.964392, 4.967567, 4.970238, 
    4.974462, 4.977457, 4.979537, 4.980639, 4.980505, 4.978874, 4.975456, 
    4.969903, 4.961752, 4.950266, 4.938305, 4.923625, 4.906556, 4.887687, 
    4.867873, 4.848182, 4.829807, 4.813938, 4.801608, 4.79357, 4.79023, 
    4.79162, 4.797441, 4.807114, 4.819869, 4.834813, 4.850992, 4.867447, 
    4.883266,
  // height(19,11, 0-49)
    4.881644, 4.880621, 4.881466, 4.883892, 4.887596, 4.892278, 4.897672, 
    4.903541, 4.909692, 4.91597, 4.922273, 4.92854, 4.934764, 4.94099, 
    4.94733, 4.949949, 4.954883, 4.959633, 4.963575, 4.966947, 4.969853, 
    4.974226, 4.977445, 4.979825, 4.981448, 4.982079, 4.9815, 4.979406, 
    4.975439, 4.968922, 4.95904, 4.948476, 4.935015, 4.918853, 4.900454, 
    4.880566, 4.860214, 4.840611, 4.823038, 4.80868, 4.798471, 4.792996, 
    4.792449, 4.796651, 4.805115, 4.817122, 4.8318, 4.8482, 4.865337, 4.882246,
  // height(19,12, 0-49)
    4.882496, 4.881999, 4.883224, 4.885882, 4.889676, 4.894325, 4.899577, 
    4.90522, 4.911082, 4.917034, 4.922996, 4.928931, 4.934853, 4.940827, 
    4.946981, 4.949989, 4.95378, 4.958515, 4.962585, 4.966149, 4.969291, 
    4.973717, 4.977075, 4.979658, 4.981715, 4.983027, 4.983429, 4.982606, 
    4.9802, 4.975337, 4.967144, 4.958006, 4.945863, 4.930773, 4.913065, 
    4.893366, 4.872625, 4.852049, 4.832983, 4.816743, 4.804437, 4.796834, 
    4.794295, 4.796777, 4.803885, 4.814964, 4.829169, 4.845552, 4.863111, 
    4.880845,
  // height(19,13, 0-49)
    4.883292, 4.883357, 4.884997, 4.887918, 4.891829, 4.896464, 4.901587, 
    4.907006, 4.912575, 4.918189, 4.923789, 4.929358, 4.934927, 4.940565, 
    4.94639, 4.950139, 4.952823, 4.957446, 4.961614, 4.96537, 4.968758, 
    4.973145, 4.976562, 4.979265, 4.981663, 4.983564, 4.98485, 4.985204, 
    4.984283, 4.981029, 4.974552, 4.966794, 4.955986, 4.942058, 4.9252, 
    4.905908, 4.885034, 4.863748, 4.84343, 4.825501, 4.811233, 4.801569, 
    4.797047, 4.797762, 4.803423, 4.813437, 4.826993, 4.84315, 4.86089, 
    4.879182,
  // height(19,14, 0-49)
    4.883975, 4.884635, 4.886726, 4.889947, 4.894012, 4.898662, 4.903681, 
    4.908897, 4.914186, 4.919464, 4.924696, 4.929881, 4.935049, 4.940267, 
    4.945613, 4.950459, 4.952142, 4.956577, 4.960824, 4.964785, 4.968439, 
    4.972709, 4.976121, 4.978877, 4.981533, 4.983922, 4.985978, 4.987384, 
    4.98782, 4.986081, 4.981294, 4.974806, 4.965281, 4.952532, 4.936615, 
    4.917893, 4.897106, 4.875359, 4.85404, 4.83465, 4.818594, 4.806993, 
    4.800546, 4.799497, 4.803661, 4.812512, 4.825278, 4.841026, 4.858731, 
    4.877334,
  // height(19,15, 0-49)
    4.884464, 4.885746, 4.888322, 4.891884, 4.896142, 4.900849, 4.905801, 
    4.910846, 4.915881, 4.920848, 4.925724, 4.930517, 4.93526, 4.939989, 
    4.94473, 4.95096, 4.951797, 4.956015, 4.960347, 4.964542, 4.968503, 
    4.972597, 4.97596, 4.978716, 4.981555, 4.984333, 4.987031, 4.989339, 
    4.990971, 4.990606, 4.987436, 4.98206, 4.973706, 4.962089, 4.94714, 
    4.929091, 4.908561, 4.886575, 4.864501, 4.843886, 4.82625, 4.812865, 
    4.804594, 4.801823, 4.804478, 4.812106, 4.823973, 4.83916, 4.856639, 
    4.875334,
  // height(19,16, 0-49)
    4.884663, 4.88658, 4.889668, 4.893605, 4.898099, 4.902907, 4.907837, 
    4.912756, 4.917584, 4.922279, 4.926834, 4.931263, 4.935582, 4.939795, 
    4.943863, 4.951606, 4.951766, 4.955799, 4.960267, 4.964756, 4.969089, 
    4.972967, 4.976264, 4.978997, 4.981962, 4.985034, 4.988237, 4.991272, 
    4.993902, 4.994734, 4.993072, 4.988607, 4.981264, 4.970675, 4.956662, 
    4.93933, 4.919178, 4.897139, 4.874533, 4.85293, 4.833932, 4.818943, 
    4.808976, 4.804556, 4.805722, 4.812094, 4.822984, 4.837489, 4.854583, 
    4.873177,
  // height(19,17, 0-49)
    4.884471, 4.887014, 4.890623, 4.894957, 4.899719, 4.904669, 4.909626, 
    4.914478, 4.919161, 4.923654, 4.92796, 4.932091, 4.936043, 4.939777, 
    4.943196, 4.952326, 4.951941, 4.9559, 4.960605, 4.965496, 4.970294, 
    4.973958, 4.977208, 4.979924, 4.982979, 4.986258, 4.989816, 4.993383, 
    4.996779, 4.998592, 4.998283, 4.994504, 4.987976, 4.978271, 4.96511, 
    4.948489, 4.928789, 4.90684, 4.883897, 4.861527, 4.841388, 4.824988, 
    4.813472, 4.8075, 4.807219, 4.81233, 4.822189, 4.835921, 4.852504, 
    4.870842,
  // height(19,18, 0-49)
    4.883793, 4.886919, 4.891025, 4.895751, 4.900793, 4.905913, 4.910947, 
    4.915798, 4.920425, 4.924825, 4.929009, 4.932978, 4.936702, 4.940094, 
    4.94299, 4.953041, 4.952164, 4.956231, 4.961337, 4.966779, 4.972184, 
    4.975669, 4.978938, 4.981686, 4.984823, 4.988232, 4.991991, 4.995869, 
    4.999767, 5.002297, 5.003136, 4.999793, 4.993859, 4.984858, 4.972429, 
    4.956472, 4.937254, 4.915499, 4.892387, 4.869453, 4.848384, 4.830771, 
    4.817868, 4.810457, 4.808792, 4.812659, 4.821465, 4.834362, 4.850341, 
    4.868311,
  // height(19,19, 0-49)
    4.882538, 4.886151, 4.890681, 4.895749, 4.901048, 4.906345, 4.911496, 
    4.916429, 4.921131, 4.92561, 4.929882, 4.933926, 4.937669, 4.94096, 
    4.943571, 4.95371, 4.952253, 4.956655, 4.962374, 4.968572, 4.974777, 
    4.978183, 4.981593, 4.984472, 4.987724, 4.991202, 4.994999, 4.998935, 
    5.003021, 5.00595, 5.007671, 5.004481, 4.998894, 4.990393, 4.978553, 
    4.963183, 4.944447, 4.922963, 4.899824, 4.876513, 4.854719, 4.836087, 
    4.821965, 4.813243, 4.810278, 4.812939, 4.820692, 4.832723, 4.848042, 
    4.865566,
  // height(19,20, 0-49)
    4.881588, 4.886601, 4.892593, 4.899169, 4.905969, 4.912692, 4.919097, 
    4.924998, 4.930258, 4.934787, 4.938541, 4.941516, 4.943758, 4.94535, 
    4.946416, 0, 4.960864, 4.963375, 4.966852, 4.970822, 4.975077, 4.975944, 
    4.977604, 4.979422, 4.982367, 4.986216, 4.99093, 4.996161, 5.00179, 
    5.006393, 5.010077, 5.007852, 5.003162, 4.995485, 4.98438, 4.969624, 
    4.951338, 4.930086, 4.906902, 4.883231, 4.860764, 4.841182, 4.825912, 
    4.815937, 4.811708, 4.813176, 4.819865, 4.831002, 4.845614, 4.862631,
  // height(19,21, 0-49)
    4.87942, 4.884988, 4.891505, 4.898539, 4.905715, 4.912723, 4.919326, 
    4.92536, 4.930717, 4.935334, 4.939191, 4.942301, 4.944708, 4.946493, 
    4.947779, 0, 4.960035, 4.963074, 4.967126, 4.971672, 4.976431, 4.976584, 
    4.977723, 4.979072, 4.98174, 4.985524, 4.990396, 4.995993, 5.002195, 
    5.007564, 5.012428, 5.010612, 5.006535, 4.999634, 4.989399, 4.975526, 
    4.958041, 4.937399, 4.914538, 4.890834, 4.867946, 4.84758, 4.831234, 
    4.819987, 4.814397, 4.814506, 4.819916, 4.829904, 4.843533, 4.859751,
  // height(19,22, 0-49)
    4.876799, 4.882879, 4.889917, 4.897455, 4.905089, 4.912499, 4.919439, 
    4.925747, 4.931327, 4.936132, 4.940154, 4.943415, 4.945968, 4.947898, 
    4.949335, 0, 4.959913, 4.963387, 4.967949, 4.973043, 4.978314, 4.977839, 
    4.978555, 4.979537, 4.982003, 4.985746, 4.990732, 4.996574, 5.003149, 
    5.009007, 5.014683, 5.012933, 5.009101, 5.002608, 4.992905, 4.97964, 
    4.962763, 4.942643, 4.920128, 4.896511, 4.873403, 4.852501, 4.835343, 
    4.823078, 4.816355, 4.815298, 4.819583, 4.828539, 4.841269, 4.856745,
  // height(19,23, 0-49)
    4.873835, 4.880381, 4.887924, 4.895979, 4.904121, 4.912008, 4.91938, 
    4.926068, 4.931972, 4.937049, 4.941298, 4.944747, 4.947457, 4.949518, 
    4.951072, 0, 4.960715, 4.964478, 4.969381, 4.974841, 4.980453, 4.979389, 
    4.979692, 4.980315, 4.982558, 4.986212, 4.991232, 4.997212, 5.004019, 
    5.010185, 5.016409, 5.014583, 5.010819, 5.004539, 4.995176, 4.982343, 
    4.96594, 4.946269, 4.924097, 4.900642, 4.877457, 4.856218, 4.838474, 
    4.825424, 4.817783, 4.815747, 4.819055, 4.827091, 4.838994, 4.853765,
  // height(19,24, 0-49)
    4.870672, 4.877634, 4.885653, 4.894224, 4.902894, 4.911297, 4.91916, 
    4.926295, 4.932595, 4.93801, 4.94254, 4.946218, 4.949106, 4.951304, 
    4.952971, 0, 4.962595, 4.966502, 4.971569, 4.977206, 4.982986, 4.981498, 
    4.981503, 4.981868, 4.98394, 4.987504, 4.992511, 4.998539, 5.005456, 
    5.011777, 5.018311, 5.016373, 5.012581, 5.006359, 4.997128, 4.984486, 
    4.968306, 4.948847, 4.926829, 4.903417, 4.880123, 4.858602, 4.840403, 
    4.826757, 4.818415, 4.815626, 4.818173, 4.82548, 4.836718, 4.850913,
  // height(19,25, 0-49)
    4.867481, 4.874813, 4.883271, 4.892335, 4.901527, 4.91046, 4.918839, 
    4.926459, 4.933195, 4.938988, 4.943835, 4.947769, 4.950856, 4.953206, 
    4.954986, 0, 4.965112, 4.969028, 4.974089, 4.979712, 4.985476, 4.983797, 
    4.983668, 4.983923, 4.985918, 4.989429, 4.994407, 5.000427, 5.007351, 
    5.013689, 5.020282, 5.018254, 5.014394, 5.008122, 4.998861, 4.986204, 
    4.970013, 4.950536, 4.92847, 4.904962, 4.881504, 4.859735, 4.841204, 
    4.827145, 4.818328, 4.815025, 4.817045, 4.823834, 4.834585, 4.848341,
  // height(19,26, 0-49)
    4.864459, 4.87211, 4.880964, 4.890482, 4.900172, 4.909622, 4.918519, 
    4.926631, 4.933817, 4.940006, 4.945184, 4.949382, 4.952669, 4.955164, 
    4.957052, 0, 4.968115, 4.971904, 4.97679, 4.98221, 4.987775, 4.986162, 
    4.986086, 4.986403, 4.988436, 4.991954, 4.996908, 5.002874, 5.009715, 
    5.015938, 5.022344, 5.020271, 5.016323, 5.009913, 5.00047, 4.98759, 
    4.971152, 4.951414, 4.929086, 4.905328, 4.881636, 4.859649, 4.840906, 
    4.826628, 4.817581, 4.814027, 4.815778, 4.822286, 4.832751, 4.846226,
  // height(19,27, 0-49)
    4.861812, 4.869731, 4.878926, 4.888848, 4.898993, 4.908931, 4.918322, 
    4.926916, 4.934547, 4.941125, 4.946622, 4.951062, 4.954522, 4.957128, 
    4.959073, 0, 4.97163, 4.975142, 4.979673, 4.984694, 4.989872, 4.988544, 
    4.988675, 4.989195, 4.991359, 4.994929, 4.999852, 5.005712, 5.012372, 
    5.018343, 5.024315, 5.022226, 5.018149, 5.011499, 5.001717, 4.988418, 
    4.971513, 4.951303, 4.928545, 4.904437, 4.880499, 4.858378, 4.839594, 
    4.825338, 4.816338, 4.812825, 4.814583, 4.821054, 4.831435, 4.844779,
  // height(19,28, 0-49)
    4.859741, 4.867873, 4.877347, 4.887616, 4.898163, 4.908547, 4.918406, 
    4.927459, 4.935514, 4.942453, 4.948228, 4.952856, 4.956412, 4.959038, 
    4.960937, 0, 4.975993, 4.979054, 4.983034, 4.987453, 4.992063, 4.991148, 
    4.991572, 4.99238, 4.994724, 4.998356, 5.003215, 5.008902, 5.015275, 
    5.020853, 5.026161, 5.024028, 5.019733, 5.012695, 5.002378, 4.988438, 
    4.970845, 4.949972, 4.926649, 4.90214, 4.87801, 4.8559, 4.837305, 
    4.823361, 4.814726, 4.811572, 4.813638, 4.820332, 4.830835, 4.844201,
  // height(19,29, 0-49)
    4.858432, 4.866712, 4.876399, 4.88695, 4.897851, 4.908648, 4.918948, 
    4.92844, 4.936892, 4.944144, 4.950123, 4.95483, 4.958349, 4.960835, 
    4.962511, 0, 4.980938, 4.983357, 4.986584, 4.990198, 4.994048, 4.993536, 
    4.994227, 4.995311, 4.997817, 5.001482, 5.006229, 5.011665, 5.017635, 
    5.022667, 5.027061, 5.024763, 5.020088, 5.012481, 5.00145, 4.986721, 
    4.968343, 4.946784, 4.922968, 4.898229, 4.874156, 4.852381, 4.834337, 
    4.821075, 4.813166, 4.810695, 4.81334, 4.820467, 4.831241, 4.8447,
  // height(19,30, 0-49)
    4.857325, 4.864811, 4.87362, 4.883223, 4.89315, 4.903017, 4.912543, 
    4.921545, 4.929926, 4.937651, 4.944711, 4.951098, 4.956753, 4.961548, 
    4.965257, 4.981699, 4.974598, 4.979191, 4.985151, 4.991585, 4.998013, 
    5.000706, 5.003804, 5.006528, 5.009774, 5.013294, 5.017124, 5.021049, 
    5.02509, 5.027961, 5.029866, 5.026049, 5.019855, 5.010766, 4.998342, 
    4.982376, 4.962988, 4.940724, 4.916574, 4.891904, 4.868294, 4.847318, 
    4.830311, 4.818207, 4.811459, 4.810057, 4.813608, 4.821434, 4.832671, 
    4.846352,
  // height(19,31, 0-49)
    4.858174, 4.865802, 4.874738, 4.884463, 4.894507, 4.904485, 4.9141, 
    4.923157, 4.931543, 4.939215, 4.946176, 4.952444, 4.958014, 4.962843, 
    4.966795, 4.981744, 4.976817, 4.98103, 4.986337, 4.99197, 4.997562, 
    5.000377, 5.003357, 5.005968, 5.009114, 5.01259, 5.016417, 5.020319, 
    5.02421, 5.026711, 5.027736, 5.023791, 5.017277, 5.007711, 4.994723, 
    4.978187, 4.958328, 4.935792, 4.911653, 4.88733, 4.8644, 4.844378, 
    4.828509, 4.817608, 4.812016, 4.811631, 4.815988, 4.824363, 4.835867, 
    4.849523,
  // height(19,32, 0-49)
    4.860078, 4.867659, 4.876506, 4.886116, 4.896039, 4.905897, 4.915404, 
    4.924363, 4.932662, 4.940258, 4.947163, 4.953413, 4.959052, 4.964091, 
    4.968487, 4.981169, 4.978074, 4.982155, 4.987026, 4.992065, 4.997014, 
    5.000091, 5.003103, 5.005722, 5.008819, 5.012202, 5.015869, 5.019507, 
    5.02294, 5.024753, 5.024618, 5.020299, 5.013247, 5.003031, 4.989363, 
    4.972216, 4.95193, 4.929254, 4.905345, 4.881649, 4.859718, 4.840992, 
    4.826592, 4.817206, 4.813052, 4.813928, 4.819293, 4.828377, 4.840262, 
    4.853956,
  // height(19,33, 0-49)
    4.863094, 4.870475, 4.879053, 4.888352, 4.897948, 4.907487, 4.916703, 
    4.925407, 4.9335, 4.940943, 4.947758, 4.953999, 4.959738, 4.965044, 
    4.969951, 4.980079, 4.97859, 4.982728, 4.987326, 4.991925, 4.996374, 
    4.999796, 5.002942, 5.005651, 5.008716, 5.011941, 5.015303, 5.018456, 
    5.021159, 5.022017, 5.020511, 5.015593, 5.007808, 4.996795, 4.982359, 
    4.964593, 4.943953, 4.921297, 4.897847, 4.875063, 4.854445, 4.837331, 
    4.824705, 4.817112, 4.814642, 4.816987, 4.823531, 4.833456, 4.845809, 
    4.859584,
  // height(19,34, 0-49)
    4.867206, 4.874252, 4.882409, 4.891233, 4.900333, 4.909385, 4.918148, 
    4.926455, 4.934219, 4.941414, 4.948065, 4.954243, 4.960041, 4.96557, 
    4.970939, 4.978593, 4.978584, 4.98288, 4.987299, 4.991557, 4.995606, 
    4.999401, 5.002732, 5.005574, 5.008594, 5.011591, 5.014505, 5.016977, 
    5.018713, 5.018397, 5.015368, 5.009659, 5.000988, 4.989071, 4.973829, 
    4.955482, 4.934607, 4.912163, 4.889425, 4.867839, 4.848833, 4.833615, 
    4.823024, 4.817452, 4.816856, 4.820828, 4.828676, 4.839528, 4.852401, 
    4.86627,
  // height(19,35, 0-49)
    4.872328, 4.878919, 4.886526, 4.89474, 4.903203, 4.911632, 4.919809, 
    4.927599, 4.934926, 4.941772, 4.948174, 4.954204, 4.959976, 4.965626, 
    4.971318, 4.976828, 4.978239, 4.982703, 4.986978, 4.990948, 4.99466, 
    4.998809, 5.002337, 5.005319, 5.008259, 5.010948, 5.01328, 5.014896, 
    5.015461, 5.013795, 5.009148, 5.002493, 4.992821, 4.979948, 4.963921, 
    4.945088, 4.92415, 4.90215, 4.880391, 4.860284, 4.843158, 4.83008, 
    4.821725, 4.818338, 4.819746, 4.825438, 4.834654, 4.84647, 4.859871, 
    4.873812,
  // height(19,36, 0-49)
    4.878319, 4.884347, 4.891294, 4.898786, 4.906506, 4.914204, 4.921698, 
    4.928871, 4.935667, 4.942079, 4.948146, 4.953941, 4.95958, 4.965217, 
    4.97104, 4.974863, 4.977667, 4.982239, 4.986354, 4.99006, 4.993469, 
    4.997919, 5.001616, 5.004714, 5.007523, 5.009817, 5.011443, 5.012049, 
    5.011275, 5.008129, 5.00182, 4.994109, 4.98338, 4.969563, 4.952835, 
    4.933675, 4.912894, 4.891598, 4.871095, 4.852732, 4.837718, 4.826962, 
    4.820982, 4.819872, 4.823338, 4.830776, 4.841359, 4.854115, 4.868001, 
    4.881951,
  // height(19,37, 0-49)
    4.884991, 4.890361, 4.896557, 4.903244, 4.910141, 4.917033, 4.923767, 
    4.930253, 4.936448, 4.942355, 4.948011, 4.953487, 4.958893, 4.964376, 
    4.97013, 4.972736, 4.976905, 4.981477, 4.985387, 4.988821, 4.991942, 
    4.996607, 5.000417, 5.003583, 5.006192, 5.008002, 5.008813, 5.008285, 
    5.006043, 5.001339, 4.993384, 4.98456, 4.972786, 4.958107, 4.940834, 
    4.921567, 4.901206, 4.880898, 4.861922, 4.845537, 4.832814, 4.824502, 
    4.820959, 4.822139, 4.827637, 4.836768, 4.848647, 4.862257, 4.876529, 
    4.890384,
  // height(19,38, 0-49)
    4.892121, 4.896754, 4.902132, 4.907953, 4.913973, 4.920011, 4.92594, 
    4.931687, 4.937231, 4.942576, 4.947761, 4.952847, 4.957928, 4.963131, 
    4.968633, 4.970451, 4.975925, 4.980362, 4.984005, 4.987148, 4.989974, 
    4.994747, 4.99859, 5.001753, 5.004083, 5.005324, 5.005226, 5.003472, 
    4.999688, 4.993407, 4.983876, 4.973956, 4.96122, 4.945838, 4.928244, 
    4.909145, 4.889503, 4.870472, 4.853275, 4.839058, 4.828744, 4.82292, 
    4.821793, 4.825191, 4.832617, 4.843311, 4.856339, 4.870652, 4.885157, 
    4.898771,
  // height(19,39, 0-49)
    4.899467, 4.903297, 4.907806, 4.912726, 4.917843, 4.923001, 4.928099, 
    4.933086, 4.937946, 4.942693, 4.947358, 4.951997, 4.95668, 4.961504, 
    4.966603, 4.967971, 4.974646, 4.978811, 4.982118, 4.984936, 4.987445, 
    4.992202, 4.995981, 4.999056, 5.00102, 5.001617, 5.000542, 4.997513, 
    4.99217, 4.984358, 4.973391, 4.962465, 4.948932, 4.93308, 4.915452, 
    4.896836, 4.878227, 4.860754, 4.845551, 4.833638, 4.825777, 4.822405, 
    4.823591, 4.829056, 4.838219, 4.850267, 4.864228, 4.879025, 4.893557, 
    4.906746,
  // height(19,40, 0-49)
    4.906766, 4.909746, 4.913357, 4.917359, 4.921566, 4.925843, 4.930111, 
    4.934331, 4.938495, 4.942622, 4.94674, 4.950891, 4.95512, 4.959492, 
    4.964085, 4.965239, 4.97296, 4.976724, 4.979627, 4.98208, 4.984232, 
    4.988842, 4.992447, 4.995337, 4.996855, 4.996744, 4.994654, 4.990354, 
    4.983506, 4.974283, 4.962084, 4.950325, 4.936236, 4.920212, 4.902885, 
    4.885092, 4.867829, 4.852161, 4.839121, 4.829577, 4.824143, 4.823107, 
    4.82642, 4.833713, 4.844347, 4.857467, 4.872072, 4.887079, 4.901387, 
    4.913939,
  // height(19,41, 0-49)
    4.913755, 4.915848, 4.918544, 4.921631, 4.924941, 4.928359, 4.931815, 
    4.935283, 4.938761, 4.942267, 4.945827, 4.949466, 4.953209, 4.957081, 
    4.961106, 4.962186, 4.970744, 4.974006, 4.976444, 4.97848, 4.980226, 
    4.984553, 4.987868, 4.990473, 4.991469, 4.990608, 4.987513, 4.982002, 
    4.973772, 4.963334, 4.950175, 4.93783, 4.923496, 4.90765, 4.890987, 
    4.874359, 4.858728, 4.845076, 4.8343, 4.827125, 4.824011, 4.825119, 
    4.830297, 4.839108, 4.850871, 4.864708, 4.879611, 4.894502, 4.908296, 
    4.919983,
  // height(19,42, 0-49)
    4.92017, 4.921348, 4.923127, 4.925314, 4.927758, 4.930353, 4.933038, 
    4.935792, 4.938614, 4.94152, 4.944527, 4.94765, 4.950894, 4.954247, 
    4.957675, 4.958741, 4.967895, 4.970575, 4.972492, 4.974058, 4.975332, 
    4.979243, 4.982157, 4.984379, 4.984793, 4.983174, 4.979122, 4.97252, 
    4.963109, 4.951718, 4.937935, 4.92532, 4.911098, 4.895811, 4.880182, 
    4.865045, 4.851295, 4.839802, 4.83133, 4.826448, 4.825478, 4.828466, 
    4.835182, 4.845138, 4.857627, 4.871772, 4.886574, 4.900981, 4.913953, 
    4.924549,
  // height(19,43, 0-49)
    4.925763, 4.926003, 4.926868, 4.928182, 4.929801, 4.931626, 4.933599, 
    4.935696, 4.937914, 4.94026, 4.942748, 4.945375, 4.948125, 4.950956, 
    4.953793, 4.954841, 4.96433, 4.966375, 4.967723, 4.968758, 4.969495, 
    4.972867, 4.975272, 4.977025, 4.97682, 4.974465, 4.969556, 4.962043, 
    4.951717, 4.939699, 4.925668, 4.913147, 4.899427, 4.885087, 4.87084, 
    4.857475, 4.845798, 4.836551, 4.830351, 4.827622, 4.828561, 4.833115, 
    4.840987, 4.851663, 4.86443, 4.878427, 4.892694, 4.906231, 4.91807, 
    4.927366,
  // height(19,44, 0-49)
    4.930317, 4.929597, 4.929554, 4.930022, 4.930867, 4.931989, 4.933323, 
    4.934839, 4.936524, 4.938376, 4.940395, 4.942565, 4.944849, 4.94718, 
    4.949445, 4.950438, 4.960001, 4.961379, 4.962115, 4.96256, 4.962694, 
    4.965418, 4.967226, 4.968439, 4.967605, 4.964572, 4.95895, 4.950758, 
    4.93984, 4.927562, 4.913687, 4.901648, 4.888824, 4.875793, 4.863242, 
    4.85188, 4.842403, 4.835417, 4.831395, 4.830625, 4.833188, 4.838951, 
    4.847569, 4.85851, 4.87108, 4.884458, 4.897746, 4.910027, 4.920442, 
    4.928277,
  // height(19,45, 0-49)
    4.933671, 4.931966, 4.931014, 4.930665, 4.930786, 4.931273, 4.932052, 
    4.933077, 4.934319, 4.935762, 4.937385, 4.939156, 4.941019, 4.942884, 
    4.944615, 4.945492, 4.954885, 4.955587, 4.955676, 4.955476, 4.954947, 
    4.956939, 4.958081, 4.958708, 4.957262, 4.953647, 4.947495, 4.938894, 
    4.92774, 4.915594, 4.902283, 4.89111, 4.879552, 4.868159, 4.857555, 
    4.848358, 4.841139, 4.836369, 4.834379, 4.835332, 4.839209, 4.845804, 
    4.854742, 4.86549, 4.877389, 4.889682, 4.901563, 4.912237, 4.920988, 
    4.927265,
  // height(19,46, 0-49)
    4.935753, 4.933025, 4.931156, 4.930007, 4.929449, 4.929368, 4.929675, 
    4.930304, 4.931202, 4.932328, 4.933641, 4.935088, 4.936592, 4.938042, 
    4.939281, 4.939974, 4.948993, 4.949016, 4.948432, 4.947545, 4.946309, 
    4.947513, 4.947949, 4.947968, 4.945961, 4.941886, 4.935413, 4.926697, 
    4.915676, 4.904049, 4.89169, 4.881741, 4.871771, 4.862283, 4.853815, 
    4.846878, 4.841915, 4.83926, 4.839114, 4.841527, 4.846392, 4.853445, 
    4.862292, 4.872415, 4.883203, 4.893989, 4.904093, 4.912873, 4.919795, 
    4.924508,
  // height(19,47, 0-49)
    4.936611, 4.932811, 4.929999, 4.92805, 4.926839, 4.926242, 4.92615, 
    4.92647, 4.927119, 4.928027, 4.929121, 4.930323, 4.931534, 4.932622, 
    4.93342, 4.933862, 4.942347, 4.941703, 4.94043, 4.938825, 4.936858, 
    4.937251, 4.936972, 4.936396, 4.933905, 4.929514, 4.922946, 4.914406, 
    4.903878, 4.893131, 4.882066, 4.873648, 4.86553, 4.858142, 4.851929, 
    4.847281, 4.844512, 4.843832, 4.84532, 4.848924, 4.854459, 4.861622, 
    4.870004, 4.879118, 4.888425, 4.897368, 4.905418, 4.912122, 4.917159, 
    4.920394,
  // height(19,48, 0-49)
    4.936437, 4.931505, 4.927708, 4.924939, 4.923077, 4.921989, 4.921544, 
    4.921619, 4.922096, 4.922868, 4.923826, 4.924857, 4.925838, 4.926618, 
    4.92702, 4.927145, 4.934983, 4.93369, 4.931725, 4.929393, 4.926692, 
    4.926288, 4.925319, 4.924188, 4.921313, 4.916768, 4.910326, 4.90224, 
    4.892526, 4.88297, 4.87348, 4.866836, 4.860761, 4.855598, 4.851686, 
    4.849298, 4.848623, 4.849751, 4.852652, 4.857186, 4.863106, 4.870075, 
    4.877688, 4.885501, 4.89306, 4.89994, 4.905788, 4.910366, 4.913583, 
    4.915535,
  // height(19,49, 0-49)
    4.939479, 4.932686, 4.927199, 4.922946, 4.919828, 4.917706, 4.916431, 
    4.915837, 4.915757, 4.916022, 4.916465, 4.916909, 4.91717, 4.917032, 
    4.916247, 4.915366, 4.929752, 4.926197, 4.921779, 4.917198, 4.912539, 
    4.913105, 4.913378, 4.914213, 4.912521, 4.90855, 4.901885, 4.89297, 
    4.881677, 4.871408, 4.861761, 4.857852, 4.85482, 4.852896, 4.852281, 
    4.853092, 4.855345, 4.858965, 4.86378, 4.869527, 4.875886, 4.882484, 
    4.888945, 4.894903, 4.900057, 4.904189, 4.907223, 4.909227, 4.910436, 
    4.91124,
  // height(20,0, 0-49)
    4.860252, 4.86001, 4.861908, 4.865577, 4.870636, 4.876714, 4.883478, 
    4.890644, 4.897981, 4.905314, 4.912512, 4.919477, 4.926129, 4.932405, 
    4.938227, 4.943402, 4.949084, 4.953224, 4.956752, 4.959602, 4.961658, 
    4.963098, 4.963417, 4.962541, 4.960215, 4.956271, 4.950531, 4.9429, 
    4.933327, 4.921966, 4.908915, 4.894793, 4.879703, 4.864185, 4.848875, 
    4.834458, 4.821619, 4.810974, 4.803027, 4.798102, 4.796328, 4.797613, 
    4.801653, 4.80796, 4.815895, 4.82473, 4.833702, 4.842091, 4.849298, 
    4.854918,
  // height(20,1, 0-49)
    4.862436, 4.862621, 4.86489, 4.86887, 4.874181, 4.880456, 4.887374, 
    4.894657, 4.902087, 4.909499, 4.91677, 4.923805, 4.93053, 4.936876, 
    4.94276, 4.947818, 4.954359, 4.958505, 4.962062, 4.965001, 4.967188, 
    4.969077, 4.969801, 4.969337, 4.967341, 4.963618, 4.957946, 4.950209, 
    4.94033, 4.92852, 4.914805, 4.900119, 4.884272, 4.867824, 4.851451, 
    4.835898, 4.821912, 4.810189, 4.8013, 4.795636, 4.793375, 4.794456, 
    4.798588, 4.805271, 4.813842, 4.823527, 4.833501, 4.842969, 4.851245, 
    4.857827,
  // height(20,2, 0-49)
    4.864428, 4.86499, 4.867573, 4.871808, 4.877315, 4.883739, 4.890766, 
    4.898131, 4.905627, 4.913094, 4.920412, 4.927494, 4.934264, 4.94065, 
    4.946568, 4.951439, 4.958696, 4.962821, 4.966372, 4.969354, 4.971641, 
    4.973957, 4.97509, 4.97507, 4.97349, 4.970134, 4.964743, 4.957186, 
    4.947346, 4.935463, 4.921481, 4.90663, 4.890397, 4.873343, 4.856158, 
    4.839617, 4.824526, 4.811648, 4.801634, 4.794953, 4.791851, 4.792322, 
    4.79611, 4.802735, 4.811536, 4.821715, 4.832422, 4.842813, 4.852137, 
    4.85981,
  // height(20,3, 0-49)
    4.866155, 4.86705, 4.869899, 4.874338, 4.879996, 4.886528, 4.893631, 
    4.90105, 4.908585, 4.916081, 4.923425, 4.930527, 4.937315, 4.943715, 
    4.949641, 4.954255, 4.962042, 4.966132, 4.969641, 4.972626, 4.974976, 
    4.977679, 4.979204, 4.979639, 4.978534, 4.975669, 4.970754, 4.963642, 
    4.954173, 4.94259, 4.928738, 4.914125, 4.897903, 4.880599, 4.862891, 
    4.845562, 4.829454, 4.815392, 4.804106, 4.796156, 4.791875, 4.791333, 
    4.794338, 4.800455, 4.809047, 4.819333, 4.830458, 4.841559, 4.851843, 
    4.860661,
  // height(20,4, 0-49)
    4.867635, 4.868824, 4.871896, 4.876496, 4.882263, 4.888866, 4.896011, 
    4.903454, 4.910999, 4.918499, 4.925837, 4.932927, 4.939702, 4.946087, 
    4.952006, 4.956291, 4.964385, 4.968431, 4.971873, 4.974825, 4.977198, 
    4.980241, 4.982126, 4.982999, 4.982406, 4.980123, 4.975844, 4.969408, 
    4.960617, 4.949678, 4.936331, 4.922343, 4.906526, 4.889344, 4.871434, 
    4.85356, 4.836578, 4.82136, 4.808711, 4.799289, 4.793529, 4.791602, 
    4.793405, 4.798576, 4.80653, 4.816529, 4.827738, 4.8393, 4.850401, 
    4.860345,
  // height(20,5, 0-49)
    4.868941, 4.870391, 4.873652, 4.878376, 4.884216, 4.890854, 4.898007, 
    4.905436, 4.912956, 4.920418, 4.927711, 4.934752, 4.941473, 4.947814, 
    4.953711, 4.957606, 4.965757, 4.969759, 4.973117, 4.976005, 4.978372, 
    4.981693, 4.983891, 4.98517, 4.985097, 4.983453, 4.979932, 4.97436, 
    4.966503, 4.956503, 4.944001, 4.930983, 4.915935, 4.899241, 4.881466, 
    4.863327, 4.845665, 4.82938, 4.815343, 4.80431, 4.796834, 4.793207, 
    4.793438, 4.797264, 4.804183, 4.813521, 4.824488, 4.836249, 4.84799, 
    4.858978,
  // height(20,6, 0-49)
    4.870184, 4.871867, 4.875287, 4.880104, 4.885983, 4.892617, 4.899735, 
    4.907109, 4.914557, 4.921935, 4.929136, 4.936078, 4.942703, 4.948964, 
    4.95482, 4.958287, 4.966236, 4.970192, 4.97346, 4.976264, 4.978598, 
    4.982133, 4.984593, 4.986225, 4.986656, 4.985677, 4.982993, 4.978419, 
    4.971696, 4.962874, 4.95149, 4.939726, 4.925767, 4.9099, 4.892593, 
    4.874488, 4.856383, 4.83918, 4.823804, 4.8111, 4.801749, 4.796178, 
    4.794536, 4.796683, 4.802223, 4.810569, 4.820991, 4.832695, 4.844877, 
    4.856782,
  // height(20,7, 0-49)
    4.871486, 4.873385, 4.876938, 4.881816, 4.887699, 4.894289, 4.901329, 
    4.908598, 4.915922, 4.923161, 4.930209, 4.936997, 4.943477, 4.949618, 
    4.955414, 4.958443, 4.965936, 4.969844, 4.97302, 4.975732, 4.978019, 
    4.981705, 4.984363, 4.986288, 4.987187, 4.986865, 4.985055, 4.981565, 
    4.976113, 4.968638, 4.958585, 4.948279, 4.935663, 4.92091, 4.904378, 
    4.886606, 4.868324, 4.850407, 4.833809, 4.819458, 4.808159, 4.800493, 
    4.796761, 4.796972, 4.800858, 4.807934, 4.81755, 4.828959, 4.841378, 
    4.854039,
  // height(20,8, 0-49)
    4.872965, 4.875064, 4.878729, 4.883643, 4.889493, 4.895999, 4.902913, 
    4.910024, 4.917163, 4.924199, 4.931038, 4.937615, 4.943896, 4.949877, 
    4.955583, 4.958203, 4.965009, 4.968857, 4.971947, 4.974571, 4.976808, 
    4.980578, 4.983373, 4.98552, 4.986834, 4.987137, 4.986202, 4.983829, 
    4.979728, 4.973704, 4.965117, 4.956395, 4.945295, 4.931881, 4.916384, 
    4.899226, 4.88104, 4.862648, 4.845007, 4.829113, 4.815887, 4.806065, 
    4.800118, 4.798223, 4.800258, 4.805854, 4.81445, 4.825356, 4.837813, 
    4.851048,
  // height(20,9, 0-49)
    4.874715, 4.877008, 4.88077, 4.885693, 4.891478, 4.897859, 4.904594, 
    4.911492, 4.918387, 4.925161, 4.931726, 4.938032, 4.944063, 4.949836, 
    4.955409, 4.957707, 4.963628, 4.967393, 4.970406, 4.972955, 4.975152, 
    4.978941, 4.981811, 4.984108, 4.985774, 4.98665, 4.986557, 4.985291, 
    4.982565, 4.978032, 4.970989, 4.96389, 4.954402, 4.942473, 4.928211, 
    4.911908, 4.894079, 4.87547, 4.857014, 4.839749, 4.824699, 4.812755, 
    4.804565, 4.800483, 4.800548, 4.804519, 4.811933, 4.82216, 4.834473, 
    4.848091,
  // height(20,10, 0-49)
    4.876799, 4.879285, 4.883133, 4.888045, 4.893735, 4.899947, 4.906461, 
    4.913087, 4.919682, 4.926131, 4.932365, 4.938345, 4.944074, 4.949587, 
    4.954967, 4.957089, 4.961978, 4.965627, 4.968569, 4.971067, 4.973243, 
    4.97699, 4.979874, 4.98225, 4.984199, 4.985584, 4.986276, 4.986076, 
    4.984701, 4.981645, 4.976162, 4.970654, 4.962789, 4.952418, 4.939521, 
    4.924259, 4.907021, 4.88845, 4.869433, 4.851023, 4.834328, 4.82038, 
    4.810005, 4.803736, 4.801787, 4.804056, 4.810177, 4.819589, 4.831591, 
    4.845403,
  // height(20,11, 0-49)
    4.879239, 4.881923, 4.885851, 4.890735, 4.896304, 4.902315, 4.908561, 
    4.91487, 4.921111, 4.927186, 4.933039, 4.938643, 4.944018, 4.949213, 
    4.954324, 4.956469, 4.960239, 4.963728, 4.966609, 4.969083, 4.971266, 
    4.974913, 4.977757, 4.980145, 4.982306, 4.984129, 4.985535, 4.986328, 
    4.986242, 4.98461, 4.980663, 4.976647, 4.97035, 4.961532, 4.950062, 
    4.935967, 4.919504, 4.901208, 4.881889, 4.862591, 4.844482, 4.828718, 
    4.816289, 4.807916, 4.80398, 4.804524, 4.80929, 4.81778, 4.829328, 
    4.843155,
  // height(20,12, 0-49)
    4.88201, 4.884904, 4.888915, 4.893763, 4.899191, 4.904974, 4.910917, 
    4.916871, 4.922716, 4.928374, 4.933802, 4.938989, 4.943964, 4.948782, 
    4.953533, 4.95595, 4.958569, 4.961857, 4.964685, 4.967168, 4.969397, 
    4.972889, 4.975645, 4.977991, 4.980297, 4.982482, 4.984518, 4.986214, 
    4.987322, 4.987028, 4.984559, 4.981891, 4.977048, 4.969718, 4.959666, 
    4.946801, 4.93125, 4.913426, 4.894051, 4.874133, 4.854875, 4.837531, 
    4.823242, 4.812902, 4.807063, 4.805912, 4.809299, 4.816798, 4.827771, 
    4.841449,
  // height(20,13, 0-49)
    4.885045, 4.888165, 4.892267, 4.897079, 4.902358, 4.907895, 4.913514, 
    4.919086, 4.924509, 4.929721, 4.934696, 4.939434, 4.943967, 4.948348, 
    4.952642, 4.955595, 4.957088, 4.960145, 4.962937, 4.965468, 4.967791, 
    4.971079, 4.973709, 4.975964, 4.978357, 4.980833, 4.98341, 4.985902, 
    4.98809, 4.989025, 4.987952, 4.986454, 4.982911, 4.976952, 4.968254, 
    4.956622, 4.942061, 4.92486, 4.905646, 4.885368, 4.865235, 4.846574, 
    4.830656, 4.818532, 4.810918, 4.808143, 4.810166, 4.816629, 4.826932, 
    4.840311,
  // height(20,14, 0-49)
    4.888229, 4.8916, 4.895807, 4.900593, 4.905726, 4.911015, 4.916304, 
    4.921482, 4.92647, 4.931225, 4.935732, 4.940003, 4.944067, 4.947958, 
    4.951711, 4.955437, 4.955875, 4.958696, 4.961479, 4.964108, 4.966577, 
    4.969624, 4.9721, 4.974234, 4.976667, 4.979364, 4.98239, 4.985562, 
    4.988698, 4.990733, 4.990968, 4.99044, 4.988013, 4.983267, 4.975816, 
    4.965367, 4.951819, 4.935346, 4.916467, 4.896061, 4.875321, 4.855616, 
    4.838318, 4.824619, 4.815388, 4.811089, 4.811786, 4.817195, 4.826753, 
    4.839705,
  // height(20,15, 0-49)
    4.891417, 4.895063, 4.899403, 4.904181, 4.909182, 4.914233, 4.919199, 
    4.923991, 4.928551, 4.932856, 4.936903, 4.940707, 4.944289, 4.947664, 
    4.950818, 4.955467, 4.954948, 4.957564, 4.96039, 4.963179, 4.965862, 
    4.968639, 4.970955, 4.972952, 4.975391, 4.978249, 4.981628, 4.985358, 
    4.989294, 4.99229, 4.993727, 4.993963, 4.99245, 4.988739, 4.982389, 
    4.973036, 4.96048, 4.944787, 4.926372, 4.906035, 4.884928, 4.864438, 
    4.846014, 4.830963, 4.820285, 4.814578, 4.81401, 4.818363, 4.827119, 
    4.839538,
  // height(20,16, 0-49)
    4.894438, 4.898385, 4.902883, 4.90768, 4.912577, 4.917415, 4.922084, 
    4.926518, 4.93068, 4.934565, 4.938181, 4.941544, 4.944665, 4.94753, 
    4.950081, 4.955651, 4.954271, 4.956758, 4.959707, 4.962741, 4.965721, 
    4.968219, 4.970386, 4.972255, 4.974681, 4.977648, 4.981289, 4.985443, 
    4.990022, 4.993821, 4.99635, 4.997137, 4.996331, 4.993463, 4.98805, 
    4.97967, 4.968042, 4.953138, 4.935272, 4.915156, 4.893888, 4.87285, 
    4.853538, 4.837351, 4.825407, 4.818417, 4.816652, 4.819967, 4.827884, 
    4.839682,
  // height(20,17, 0-49)
    4.897111, 4.901378, 4.906057, 4.910903, 4.915725, 4.920388, 4.924805, 
    4.92893, 4.93275, 4.936276, 4.939528, 4.942516, 4.945239, 4.947652, 
    4.949658, 4.955938, 4.95375, 4.956237, 4.959424, 4.962814, 4.966193, 
    4.968428, 4.970485, 4.972262, 4.974679, 4.977714, 4.981524, 4.985966, 
    4.991012, 4.995444, 4.99893, 5.000061, 4.999754, 4.997528, 4.992876, 
    4.985324, 4.974533, 4.960389, 4.943113, 4.92333, 4.90207, 4.880688, 
    4.860705, 4.843585, 4.830546, 4.822402, 4.819518, 4.82182, 4.828876, 
    4.839989,
  // height(20,18, 0-49)
    4.899259, 4.903844, 4.908713, 4.913628, 4.918412, 4.922945, 4.927167, 
    4.931057, 4.934627, 4.9379, 4.940901, 4.943637, 4.946083, 4.948168, 
    4.94976, 4.956294, 4.953275, 4.955921, 4.959491, 4.963376, 4.967283, 
    4.969299, 4.971318, 4.973071, 4.97551, 4.97859, 4.98248, 4.987064, 
    4.992386, 4.997256, 5.001545, 5.002809, 5.002788, 5.001004, 4.996927, 
    4.990052, 4.979986, 4.966546, 4.949867, 4.930487, 4.909364, 4.887812, 
    4.867347, 4.849483, 4.83551, 4.826337, 4.822413, 4.823737, 4.829926, 
    4.840314,
  // height(20,19, 0-49)
    4.900722, 4.905582, 4.910621, 4.915603, 4.920366, 4.924819, 4.928921, 
    4.932685, 4.936142, 4.939328, 4.942264, 4.944942, 4.947306, 4.949254, 
    4.950626, 4.956723, 4.952731, 4.955709, 4.959822, 4.964365, 4.968961, 
    4.970843, 4.972939, 4.974776, 4.977301, 4.980426, 4.984317, 4.988889, 
    4.994273, 4.99935, 5.004237, 5.005415, 5.005468, 5.00392, 5.000231, 
    4.993872, 4.984408, 4.971598, 4.9555, 4.936566, 4.915679, 4.894096, 
    4.873318, 4.854876, 4.840123, 4.83004, 4.825162, 4.825555, 4.830888, 
    4.840529,
  // height(20,20, 0-49)
    4.90239, 4.908547, 4.914843, 4.921025, 4.926898, 4.932327, 4.937214, 
    4.9415, 4.945158, 4.948183, 4.950596, 4.952441, 4.953793, 4.954744, 
    4.955407, 0, 4.958249, 4.960236, 4.962961, 4.965996, 4.969181, 4.968955, 
    4.969491, 4.97025, 4.972277, 4.975456, 4.979868, 4.985317, 4.991841, 
    4.998215, 5.004694, 5.006587, 5.007314, 5.006402, 5.00332, 4.997553, 
    4.988664, 4.976397, 4.960779, 4.942212, 4.921516, 4.899904, 4.878851, 
    4.859899, 4.844436, 4.83351, 4.827723, 4.827208, 4.831687, 4.840559,
  // height(20,21, 0-49)
    4.902546, 4.909152, 4.915813, 4.922264, 4.928308, 4.93382, 4.938725, 
    4.942987, 4.946609, 4.949608, 4.952027, 4.953918, 4.955361, 4.956449, 
    4.957307, 0, 4.95625, 4.958742, 4.96202, 4.965616, 4.96931, 4.968532, 
    4.968688, 4.969118, 4.970976, 4.974154, 4.978734, 4.984498, 4.991485, 
    4.998459, 5.005868, 5.007966, 5.009057, 5.008655, 5.006201, 5.001147, 
    4.99302, 4.981514, 4.966591, 4.948582, 4.928237, 4.906707, 4.885434, 
    4.865964, 4.849724, 4.837832, 4.830966, 4.829334, 4.832719, 4.840568,
  // height(20,22, 0-49)
    4.902033, 4.909122, 4.916215, 4.92303, 4.929366, 4.935092, 4.940144, 
    4.944501, 4.948182, 4.951223, 4.953678, 4.955619, 4.957127, 4.958311, 
    4.959311, 0, 4.955119, 4.958027, 4.96179, 4.965904, 4.970087, 4.968813, 
    4.968649, 4.968804, 4.970531, 4.973706, 4.978404, 4.984384, 4.991682, 
    4.999045, 5.007104, 5.009167, 5.010358, 5.010189, 5.00809, 5.003501, 
    4.995925, 4.985018, 4.970692, 4.953214, 4.933263, 4.911923, 4.89059, 
    4.870792, 4.853981, 4.841319, 4.833551, 4.830953, 4.833365, 4.84028,
  // height(20,23, 0-49)
    4.900946, 4.908532, 4.916096, 4.92334, 4.930048, 4.936085, 4.941385, 
    4.945931, 4.949752, 4.952897, 4.955433, 4.95744, 4.959013, 4.96027, 
    4.961375, 0, 4.954969, 4.958154, 4.962238, 4.966699, 4.971208, 4.969459, 
    4.96897, 4.968847, 4.970413, 4.973536, 4.978281, 4.984387, 4.991886, 
    4.999502, 5.008006, 5.009949, 5.011131, 5.011066, 5.009185, 5.00492, 
    4.99776, 4.987338, 4.973525, 4.956533, 4.936977, 4.915878, 4.894584, 
    4.874597, 4.857371, 4.844103, 4.835588, 4.832156, 4.833704, 4.839765,
  // height(20,24, 0-49)
    4.899428, 4.907504, 4.915555, 4.92326, 4.930388, 4.936795, 4.942407, 
    4.947209, 4.951232, 4.95453, 4.957183, 4.959279, 4.96092, 4.962241, 
    4.963425, 0, 4.95597, 4.959291, 4.963529, 4.968157, 4.972827, 4.970741, 
    4.970021, 4.969701, 4.971145, 4.974215, 4.978966, 4.985128, 4.992729, 
    5.000482, 5.009243, 5.011076, 5.012208, 5.012159, 5.010361, 5.006243, 
    4.999289, 4.98912, 4.975582, 4.958858, 4.939522, 4.918553, 4.897259, 
    4.877122, 4.859592, 4.845881, 4.836812, 4.832757, 4.833642, 4.839036,
  // height(20,25, 0-49)
    4.897653, 4.906196, 4.91472, 4.922887, 4.93045, 4.937253, 4.943209, 
    4.948304, 4.952564, 4.956049, 4.958841, 4.961037, 4.962751, 4.964127, 
    4.965363, 0, 4.957728, 4.961046, 4.96527, 4.969884, 4.974544, 4.972311, 
    4.971497, 4.971106, 4.972506, 4.975554, 4.980302, 4.986476, 4.994102, 
    5.001885, 5.010712, 5.012488, 5.013579, 5.013506, 5.011698, 5.007585, 
    5.000655, 4.990522, 4.977032, 4.960351, 4.941041, 4.920062, 4.898702, 
    4.878432, 4.860693, 4.846697, 4.837277, 4.832819, 4.833266, 4.838201,
  // height(20,26, 0-49)
    4.895818, 4.904783, 4.913742, 4.922344, 4.930325, 4.937515, 4.943821, 
    4.949216, 4.953726, 4.957407, 4.960343, 4.962636, 4.964409, 4.965817, 
    4.967063, 0, 4.960133, 4.963308, 4.967357, 4.971776, 4.976251, 4.974082, 
    4.973327, 4.973009, 4.974462, 4.977538, 4.982289, 4.98844, 4.996022, 
    5.003737, 5.012439, 5.014235, 5.015309, 5.015183, 5.013282, 5.009041, 
    5.001948, 4.99163, 4.97794, 4.961062, 4.941566, 4.920424, 4.898925, 
    4.878536, 4.860688, 4.846581, 4.837034, 4.832421, 4.832682, 4.8374,
  // height(20,27, 0-49)
    4.894114, 4.903435, 4.912771, 4.921757, 4.930116, 4.937665, 4.944301, 
    4.949985, 4.954732, 4.958596, 4.961658, 4.964022, 4.965817, 4.967206, 
    4.968397, 0, 4.96324, 4.966122, 4.969824, 4.973864, 4.97798, 4.976048, 
    4.975473, 4.975338, 4.976915, 4.98005, 4.984796, 4.990885, 4.998345, 
    5.00589, 5.014274, 5.016143, 5.01721, 5.016988, 5.014902, 5.010391, 
    5.002958, 4.992247, 4.978143, 4.960862, 4.941015, 4.919603, 4.897938, 
    4.87749, 4.859674, 4.845661, 4.836235, 4.831735, 4.832074, 4.836821,
  // height(20,28, 0-49)
    4.892716, 4.902316, 4.911954, 4.921258, 4.92994, 4.937809, 4.94474, 
    4.950686, 4.955645, 4.959659, 4.962801, 4.965176, 4.966919, 4.9682, 
    4.969231, 0, 4.967395, 4.969824, 4.972999, 4.976473, 4.980055, 4.978459, 
    4.97812, 4.978223, 4.979947, 4.983134, 4.987837, 4.993802, 5.001053, 
    5.008318, 5.016205, 5.018162, 5.019183, 5.018777, 5.016371, 5.011417, 
    5.00344, 4.992121, 4.977393, 4.95953, 4.939205, 4.917471, 4.895676, 
    4.875288, 4.8577, 4.844033, 4.835011, 4.830916, 4.831614, 4.836638,
  // height(20,29, 0-49)
    4.891768, 4.901561, 4.91142, 4.920973, 4.929929, 4.938075, 4.945275, 
    4.951451, 4.956579, 4.960682, 4.963824, 4.966108, 4.967679, 4.968717, 
    4.969442, 0, 4.972353, 4.974166, 4.976633, 4.979355, 4.982222, 4.980926, 
    4.980772, 4.981068, 4.982892, 4.986081, 4.990681, 4.996451, 5.003397, 
    5.010265, 5.017463, 5.019434, 5.020311, 5.019595, 5.016734, 5.011202, 
    5.002559, 4.990538, 4.975133, 4.956691, 4.935954, 4.914032, 4.892297, 
    4.872213, 4.855128, 4.842093, 4.833755, 4.830319, 4.831594, 4.837072,
  // height(20,30, 0-49)
    4.890552, 4.899473, 4.908428, 4.917069, 4.925149, 4.932522, 4.939125, 
    4.94497, 4.950115, 4.954631, 4.958583, 4.961999, 4.964857, 4.967066, 
    4.968472, 4.979602, 4.96907, 4.971892, 4.976008, 4.980648, 4.98542, 
    4.986781, 4.988743, 4.990612, 4.993301, 4.996634, 5.000715, 5.005429, 
    5.010921, 5.01609, 5.021275, 5.022079, 5.021772, 5.019878, 5.015864, 
    5.009229, 4.99956, 4.986626, 4.970476, 4.951515, 4.930534, 4.90868, 
    4.887331, 4.867914, 4.851709, 4.839678, 4.832371, 4.829907, 4.832027, 
    4.838179,
  // height(20,31, 0-49)
    4.890921, 4.899925, 4.908952, 4.91766, 4.925797, 4.93321, 4.939828, 
    4.945653, 4.950732, 4.95514, 4.958956, 4.962236, 4.965003, 4.967213, 
    4.968752, 4.979363, 4.971177, 4.97361, 4.977141, 4.98109, 4.985148, 
    4.986675, 4.988585, 4.990395, 4.993023, 4.996342, 5.00046, 5.005226, 
    5.010689, 5.015679, 5.020274, 5.021196, 5.02085, 5.01876, 5.014407, 
    5.007318, 4.997122, 4.983652, 4.967027, 4.947731, 4.926632, 4.904924, 
    4.883998, 4.865252, 4.849897, 4.83881, 4.832448, 4.830843, 4.833675, 
    4.840341,
  // height(20,32, 0-49)
    4.891858, 4.900726, 4.909607, 4.918174, 4.926184, 4.933486, 4.940012, 
    4.945757, 4.950766, 4.955113, 4.958885, 4.962158, 4.964985, 4.967364, 
    4.969228, 4.978518, 4.972463, 4.974708, 4.977826, 4.98125, 4.984755, 
    4.986572, 4.988569, 4.990442, 4.993085, 4.996394, 5.000472, 5.005139, 
    5.010365, 5.014951, 5.01875, 5.019603, 5.019039, 5.016583, 5.011744, 
    5.004078, 4.993276, 4.979236, 4.962163, 4.942626, 4.921564, 4.900208, 
    4.879947, 4.86213, 4.847888, 4.837993, 4.832799, 4.832254, 4.835965, 
    4.843286,
  // height(20,33, 0-49)
    4.893402, 4.901961, 4.910522, 4.918782, 4.926514, 4.933579, 4.93991, 
    4.945505, 4.950407, 4.954688, 4.958445, 4.961763, 4.964719, 4.96735, 
    4.96964, 4.977197, 4.973083, 4.975312, 4.978167, 4.981205, 4.984287, 
    4.986477, 4.98866, 4.990693, 4.993394, 4.996678, 5.000629, 5.005051, 
    5.009844, 5.013827, 5.016671, 5.017282, 5.016326, 5.013347, 5.00788, 
    4.999536, 4.988063, 4.973445, 4.955978, 4.936319, 4.915467, 4.894683, 
    4.87533, 4.858694, 4.845803, 4.83732, 4.833489, 4.834168, 4.838899, 
    4.846986,
  // height(20,34, 0-49)
    4.89555, 4.903658, 4.911766, 4.919588, 4.926923, 4.933646, 4.939695, 
    4.945072, 4.949821, 4.954011, 4.957741, 4.961105, 4.964197, 4.967091, 
    4.969819, 4.975549, 4.97322, 4.975553, 4.978248, 4.981001, 4.983756, 
    4.986354, 4.988786, 4.991036, 4.993814, 4.997042, 5.000778, 5.004812, 
    5.008993, 5.012204, 5.01397, 5.014173, 5.01267, 5.009023, 5.002813, 
    4.993709, 4.981535, 4.966369, 4.9486, 4.928967, 4.908524, 4.88854, 
    4.870338, 4.855117, 4.843793, 4.836905, 4.834589, 4.836618, 4.842463, 
    4.851387,
  // height(20,35, 0-49)
    4.898267, 4.905814, 4.913355, 4.920641, 4.92749, 4.933788, 4.939488, 
    4.944591, 4.949139, 4.953203, 4.956876, 4.960257, 4.963455, 4.966567, 
    4.969674, 4.973719, 4.973058, 4.975548, 4.978137, 4.98067, 4.983167, 
    4.986171, 4.988875, 4.991373, 4.994223, 4.997348, 5.000774, 5.004288, 
    5.007689, 5.009979, 5.010575, 5.010211, 5.008013, 5.003575, 4.996533, 
    4.986623, 4.973759, 4.958113, 4.940172, 4.920749, 4.900939, 4.881996, 
    4.865181, 4.851587, 4.842009, 4.83686, 4.836168, 4.83962, 4.846628, 
    4.856417,
  // height(20,36, 0-49)
    4.901495, 4.908389, 4.915284, 4.921958, 4.92825, 4.934066, 4.939364, 
    4.944149, 4.948456, 4.952359, 4.955939, 4.959299, 4.962548, 4.965801, 
    4.969179, 4.971826, 4.972733, 4.975375, 4.977877, 4.980225, 4.982509, 
    4.985884, 4.988856, 4.991599, 4.994495, 4.99746, 5.00048, 5.003342, 
    5.005812, 5.007051, 5.006406, 5.005326, 5.002304, 4.996975, 4.989042, 
    4.97832, 4.964816, 4.948807, 4.930867, 4.911874, 4.892938, 4.87528, 
    4.860076, 4.848299, 4.84061, 4.837299, 4.838289, 4.843188, 4.85136, 
    4.861993,
  // height(20,37, 0-49)
    4.905167, 4.911334, 4.917521, 4.923526, 4.929215, 4.934506, 4.939363, 
    4.943795, 4.947833, 4.95154, 4.954994, 4.958288, 4.961529, 4.964836, 
    4.968349, 4.969948, 4.972336, 4.975077, 4.977478, 4.979656, 4.981754, 
    4.985441, 4.988646, 4.991607, 4.994504, 4.99724, 4.999755, 5.001844, 
    5.003247, 5.003323, 5.001387, 4.999458, 4.995503, 4.989217, 4.980371, 
    4.968874, 4.954834, 4.938624, 4.9209, 4.902584, 4.884777, 4.868644, 
    4.855253, 4.845448, 4.839749, 4.838326, 4.841006, 4.847328, 4.856611, 
    4.868018,
  // height(20,38, 0-49)
    4.909193, 4.914583, 4.920015, 4.925317, 4.930371, 4.935106, 4.939497, 
    4.943548, 4.947289, 4.950776, 4.954073, 4.957259, 4.960435, 4.96371, 
    4.967225, 4.968122, 4.971893, 4.974655, 4.976923, 4.97893, 4.980852, 
    4.984771, 4.988155, 4.991285, 4.994119, 4.996551, 4.998464, 4.999669, 
    4.999884, 4.99871, 4.995449, 4.992558, 4.987595, 4.98032, 4.970589, 
    4.958406, 4.943982, 4.927779, 4.910518, 4.893145, 4.876726, 4.862342, 
    4.85094, 4.84322, 4.839568, 4.840035, 4.844362, 4.852028, 4.862319, 
    4.874377,
  // height(20,39, 0-49)
    4.913477, 4.918053, 4.922704, 4.927279, 4.931678, 4.93584, 4.939745, 
    4.943396, 4.946823, 4.950062, 4.953173, 4.956218, 4.959277, 4.962446, 
    4.965847, 4.966341, 4.971383, 4.974071, 4.976166, 4.977993, 4.979737, 
    4.983795, 4.987283, 4.990516, 4.993211, 4.995252, 4.99647, 4.996691, 
    4.995628, 4.99314, 4.988544, 4.984612, 4.978605, 4.970356, 4.959818, 
    4.94709, 4.932482, 4.916533, 4.900011, 4.883851, 4.869068, 4.856631, 
    4.847351, 4.841784, 4.840184, 4.842492, 4.848373, 4.857256, 4.868401, 
    4.880943,
  // height(20,40, 0-49)
    4.917906, 4.921646, 4.925501, 4.929339, 4.933074, 4.936653, 4.940061, 
    4.9433, 4.946392, 4.949367, 4.952266, 4.955137, 4.958039, 4.961041, 
    4.964238, 4.964564, 4.970736, 4.97326, 4.975143, 4.976772, 4.978323, 
    4.982419, 4.985922, 4.989172, 4.991644, 4.993212, 4.993649, 4.99281, 
    4.990404, 4.98657, 4.980658, 4.975645, 4.968606, 4.959457, 4.948241, 
    4.93516, 4.920611, 4.905192, 4.889691, 4.87501, 4.86208, 4.851747, 
    4.844676, 4.84128, 4.841683, 4.845729, 4.853019, 4.862945, 4.874746, 
    4.887564,
  // height(20,41, 0-49)
    4.922345, 4.925241, 4.928298, 4.9314, 4.934471, 4.937466, 4.940372, 
    4.943191, 4.945935, 4.948627, 4.951293, 4.953965, 4.956676, 4.95947, 
    4.9624, 4.962718, 4.969854, 4.972135, 4.973769, 4.975179, 4.976512, 
    4.980538, 4.983962, 4.987133, 4.989291, 4.9903, 4.98989, 4.987938, 
    4.984165, 4.978992, 4.971818, 4.965739, 4.957735, 4.94781, 4.936104, 
    4.92291, 4.908694, 4.894094, 4.879889, 4.866925, 4.856025, 4.847902, 
    4.84307, 4.841802, 4.844105, 4.849738, 4.858246, 4.868992, 4.881212, 
    4.894058,
  // height(20,42, 0-49)
    4.926642, 4.928699, 4.930964, 4.93334, 4.935758, 4.938178, 4.940584, 
    4.942979, 4.945368, 4.947763, 4.950179, 4.95263, 4.955127, 4.957681, 
    4.960309, 4.96071, 4.96862, 4.970598, 4.971952, 4.973114, 4.974197, 
    4.978046, 4.981288, 4.98428, 4.986035, 4.986415, 4.985108, 4.982025, 
    4.976905, 4.970449, 4.962109, 4.955034, 4.946192, 4.935675, 4.923714, 
    4.910677, 4.897085, 4.88359, 4.870934, 4.859879, 4.851132, 4.845262, 
    4.842635, 4.843394, 4.847439, 4.854456, 4.863945, 4.875252, 4.887619, 
    4.900222,
  // height(20,43, 0-49)
    4.930626, 4.931849, 4.933344, 4.935014, 4.936798, 4.938658, 4.940579, 
    4.942554, 4.944587, 4.94668, 4.948834, 4.951047, 4.953313, 4.955612, 
    4.957922, 4.958442, 4.966921, 4.968552, 4.9696, 4.970482, 4.971275, 
    4.974844, 4.977806, 4.980515, 4.981785, 4.981482, 4.979256, 4.975064, 
    4.968668, 4.961029, 4.951668, 4.943729, 4.934234, 4.923361, 4.911418, 
    4.898832, 4.886153, 4.874021, 4.86312, 4.854114, 4.847578, 4.843935, 
    4.843416, 4.846041, 4.851618, 4.85977, 4.869962, 4.881538, 4.893755, 
    4.905829,
  // height(20,44, 0-49)
    4.93411, 4.934515, 4.935261, 4.936253, 4.937433, 4.938762, 4.940217, 
    4.941791, 4.943477, 4.94527, 4.94716, 4.949131, 4.951157, 4.953195, 
    4.955183, 4.955816, 4.964656, 4.965913, 4.966628, 4.967195, 4.967651, 
    4.970848, 4.973435, 4.975765, 4.976482, 4.975461, 4.972332, 4.967094, 
    4.959548, 4.950883, 4.940692, 4.93208, 4.922171, 4.911213, 4.89958, 
    4.887739, 4.876243, 4.865695, 4.856701, 4.849814, 4.845474, 4.843967, 
    4.845396, 4.84967, 4.856519, 4.865516, 4.876104, 4.887634, 4.899394, 
    4.910653,
  // height(20,45, 0-49)
    4.936903, 4.936502, 4.936521, 4.936871, 4.937485, 4.938321, 4.939349, 
    4.940551, 4.941915, 4.943424, 4.945058, 4.946791, 4.948578, 4.950358, 
    4.952039, 4.952745, 4.961742, 4.962612, 4.962971, 4.963184, 4.963254, 
    4.965993, 4.968124, 4.96999, 4.970107, 4.968362, 4.964381, 4.958209, 
    4.949688, 4.940206, 4.929422, 4.920379, 4.910328, 4.899585, 4.888559, 
    4.877738, 4.867655, 4.858856, 4.851855, 4.847086, 4.844861, 4.845332, 
    4.848487, 4.854145, 4.861969, 4.87149, 4.882148, 4.893308, 4.904304, 
    4.914479,
  // height(20,46, 0-49)
    4.938819, 4.937624, 4.936943, 4.936685, 4.936779, 4.93717, 4.937817, 
    4.938693, 4.939772, 4.94103, 4.942434, 4.943947, 4.945509, 4.947042, 
    4.948433, 4.949158, 4.958127, 4.958603, 4.958583, 4.958401, 4.958039, 
    4.960252, 4.961856, 4.963193, 4.962687, 4.960245, 4.955501, 4.948549, 
    4.939279, 4.929226, 4.918125, 4.908927, 4.899035, 4.888804, 4.878668, 
    4.869109, 4.860616, 4.853668, 4.848677, 4.845958, 4.845698, 4.847935, 
    4.852553, 4.859291, 4.86776, 4.877473, 4.887864, 4.898334, 4.908283, 
    4.91715,
  // height(20,47, 0-49)
    4.93972, 4.937729, 4.936366, 4.935534, 4.935153, 4.935151, 4.935477, 
    4.936083, 4.936932, 4.937986, 4.939202, 4.940526, 4.941891, 4.9432, 
    4.944324, 4.945001, 4.953781, 4.953864, 4.95344, 4.952825, 4.951988, 
    4.953621, 4.954652, 4.955418, 4.954295, 4.951216, 4.945836, 4.938297, 
    4.928536, 4.918194, 4.907071, 4.898016, 4.888585, 4.879151, 4.870152, 
    4.862043, 4.85526, 4.850199, 4.847168, 4.84637, 4.847877, 4.851622, 
    4.857403, 4.864896, 4.873673, 4.883236, 4.893039, 4.902533, 4.911198, 
    4.918588,
  // height(20,48, 0-49)
    4.939519, 4.93672, 4.934682, 4.933303, 4.932487, 4.932148, 4.932213, 
    4.932616, 4.933301, 4.934213, 4.935294, 4.936477, 4.937681, 4.938794, 
    4.939677, 4.940239, 4.948703, 4.94839, 4.94754, 4.946457, 4.945107, 
    4.946132, 4.946567, 4.946746, 4.945043, 4.94142, 4.935561, 4.927656, 
    4.917686, 4.907351, 4.896503, 4.88789, 4.879201, 4.870818, 4.863158, 
    4.856635, 4.85162, 4.848419, 4.847244, 4.848188, 4.851223, 4.856192, 
    4.862821, 4.870739, 4.879495, 4.888591, 4.89752, 4.905799, 4.913006, 
    4.918834,
  // height(20,49, 0-49)
    4.940613, 4.936409, 4.933164, 4.930776, 4.929138, 4.928135, 4.927667, 
    4.927631, 4.927937, 4.928491, 4.9292, 4.92996, 4.930647, 4.931097, 
    4.931102, 4.930818, 4.946164, 4.943949, 4.940964, 4.937904, 4.934816, 
    4.936986, 4.938692, 4.94071, 4.939893, 4.93633, 4.929495, 4.919771, 
    4.907046, 4.894641, 4.882136, 4.8747, 4.867539, 4.861034, 4.855579, 
    4.851521, 4.849131, 4.84859, 4.849968, 4.853214, 4.858169, 4.864559, 
    4.872037, 4.88018, 4.888537, 4.896647, 4.90409, 4.910515, 4.915682, 
    4.919499,
  // height(21,0, 0-49)
    4.867756, 4.87136, 4.876185, 4.881904, 4.888227, 4.894917, 4.901782, 
    4.908686, 4.915534, 4.922264, 4.928842, 4.935246, 4.941461, 4.947464, 
    4.953222, 4.958513, 4.964422, 4.96916, 4.973463, 4.977247, 4.98037, 
    4.982961, 4.984521, 4.984962, 4.984047, 4.981614, 4.977492, 4.971577, 
    4.963781, 4.95417, 4.942726, 4.929893, 4.915575, 4.900093, 4.883879, 
    4.867457, 4.851445, 4.836494, 4.823259, 4.812335, 4.804196, 4.799148, 
    4.797297, 4.798529, 4.802532, 4.808812, 4.816741, 4.82561, 4.834689, 
    4.843285,
  // height(21,1, 0-49)
    4.869227, 4.873135, 4.878213, 4.88414, 4.890633, 4.897455, 4.904428, 
    4.911416, 4.918332, 4.925114, 4.931731, 4.938162, 4.944387, 4.950385, 
    4.956112, 4.961147, 4.967659, 4.972268, 4.976444, 4.980152, 4.983257, 
    4.986171, 4.988067, 4.988924, 4.988447, 4.98646, 4.982759, 4.977232, 
    4.969764, 4.960455, 4.949201, 4.93672, 4.922586, 4.907089, 4.890637, 
    4.87375, 4.857055, 4.841236, 4.827, 4.815002, 4.805791, 4.799745, 
    4.797029, 4.797587, 4.801143, 4.807224, 4.815208, 4.824379, 4.833981, 
    4.843285,
  // height(21,2, 0-49)
    4.87042, 4.874584, 4.879874, 4.885972, 4.892601, 4.899534, 4.906593, 
    4.913648, 4.920613, 4.927431, 4.934066, 4.940497, 4.946706, 4.952666, 
    4.958333, 4.963048, 4.970029, 4.974471, 4.978471, 4.982044, 4.985077, 
    4.988253, 4.990441, 4.991687, 4.991656, 4.99017, 4.987002, 4.982033, 
    4.97512, 4.966384, 4.955632, 4.943846, 4.930265, 4.915128, 4.898799, 
    4.881767, 4.864641, 4.848114, 4.832927, 4.819794, 4.809337, 4.802019, 
    4.798089, 4.79757, 4.800246, 4.805697, 4.813336, 4.822461, 4.832316, 
    4.842153,
  // height(21,3, 0-49)
    4.871417, 4.875794, 4.881257, 4.88749, 4.894225, 4.90124, 4.90836, 
    4.91546, 4.922452, 4.92928, 4.935906, 4.942309, 4.948469, 4.954359, 
    4.959938, 4.964278, 4.971559, 4.975809, 4.979591, 4.982981, 4.985889, 
    4.989264, 4.991691, 4.993279, 4.993685, 4.992729, 4.990175, 4.985899, 
    4.979735, 4.971802, 4.96182, 4.951028, 4.938334, 4.923909, 4.908056, 
    4.891205, 4.873922, 4.856891, 4.840857, 4.826586, 4.81477, 4.805964, 
    4.800524, 4.798568, 4.799973, 4.804396, 4.811304, 4.820037, 4.829866, 
    4.840038,
  // height(21,4, 0-49)
    4.872332, 4.876885, 4.882481, 4.888814, 4.895623, 4.902688, 4.909839, 
    4.916954, 4.923941, 4.930746, 4.937329, 4.943668, 4.949744, 4.955535, 
    4.961005, 4.964917, 4.972301, 4.976346, 4.979885, 4.983051, 4.985792, 
    4.989301, 4.991906, 4.993781, 4.994592, 4.994171, 4.992283, 4.9888, 
    4.983535, 4.976586, 4.967588, 4.958031, 4.946498, 4.933095, 4.91804, 
    4.90169, 4.884544, 4.867239, 4.850518, 4.835167, 4.821952, 4.811521, 
    4.804342, 4.800659, 4.800459, 4.8035, 4.809333, 4.817359, 4.826887, 
    4.837183,
  // height(21,5, 0-49)
    4.873298, 4.87799, 4.883683, 4.890078, 4.896924, 4.904002, 4.91115, 
    4.91824, 4.925184, 4.931925, 4.938425, 4.94466, 4.950615, 4.956275, 
    4.961616, 4.965065, 4.972339, 4.976171, 4.979454, 4.982371, 4.984913, 
    4.988491, 4.99121, 4.993308, 4.994482, 4.994578, 4.993377, 4.990749, 
    4.986489, 4.980652, 4.972798, 4.964639, 4.954481, 4.942347, 4.928371, 
    4.912815, 4.896089, 4.878769, 4.861557, 4.845256, 4.830675, 4.818562, 
    4.809506, 4.803884, 4.801821, 4.803196, 4.807662, 4.8147, 4.823673, 
    4.833878,
  // height(21,6, 0-49)
    4.874443, 4.879241, 4.884993, 4.891414, 4.898254, 4.905306, 4.912405, 
    4.919427, 4.926284, 4.932917, 4.939289, 4.945377, 4.951174, 4.956671, 
    4.961865, 4.964837, 4.971784, 4.975398, 4.97842, 4.981078, 4.983403, 
    4.986985, 4.989758, 4.992006, 4.993488, 4.994068, 4.99355, 4.991801, 
    4.988611, 4.983963, 4.977353, 4.970687, 4.962039, 4.951355, 4.938675, 
    4.924161, 4.908125, 4.891047, 4.87358, 4.856506, 4.840674, 4.826908, 
    4.815924, 4.808243, 4.804142, 4.803638, 4.806506, 4.812325, 4.820523, 
    4.830435,
  // height(21,7, 0-49)
    4.87588, 4.880752, 4.88653, 4.892937, 4.899731, 4.90671, 4.913714, 
    4.920619, 4.927339, 4.933815, 4.940012, 4.945911, 4.951509, 4.956812, 
    4.961838, 4.964347, 4.970757, 4.97415, 4.976916, 4.979318, 4.981421, 
    4.98495, 4.987716, 4.990044, 4.991772, 4.992788, 4.992926, 4.992055, 
    4.989957, 4.986527, 4.981206, 4.976059, 4.968983, 4.959855, 4.948626, 
    4.93535, 4.92023, 4.903647, 4.886172, 4.868548, 4.851635, 4.836328, 
    4.823456, 4.813686, 4.807459, 4.804945, 4.806056, 4.810474, 4.81771, 
    4.82715,
  // height(21,8, 0-49)
    4.8777, 4.882618, 4.888388, 4.894741, 4.901444, 4.908303, 4.915162, 
    4.9219, 4.928433, 4.934703, 4.940678, 4.946343, 4.951704, 4.95678, 
    4.961609, 4.963711, 4.969393, 4.972557, 4.975082, 4.977241, 4.979133, 
    4.982553, 4.985257, 4.987593, 4.989506, 4.990901, 4.99165, 4.991627, 
    4.990613, 4.988391, 4.984363, 4.980696, 4.975188, 4.967651, 4.957954, 
    4.946052, 4.932031, 4.916164, 4.898924, 4.880996, 4.863228, 4.846558, 
    4.831919, 4.82012, 4.811763, 4.807185, 4.806442, 4.80934, 4.81547, 
    4.824277,
  // height(21,9, 0-49)
    4.879959, 4.884899, 4.890628, 4.89689, 4.903462, 4.910154, 4.916817, 
    4.923337, 4.929632, 4.935648, 4.941355, 4.946746, 4.951833, 4.956645, 
    4.961241, 4.963027, 4.967825, 4.970748, 4.97305, 4.974993, 4.976692, 
    4.979956, 4.982547, 4.98483, 4.986863, 4.988575, 4.989882, 4.990657, 
    4.99069, 4.989635, 4.986869, 4.984592, 4.98059, 4.974617, 4.966471, 
    4.956012, 4.943221, 4.928251, 4.911475, 4.893493, 4.87512, 4.857318, 
    4.8411, 4.827405, 4.816993, 4.810369, 4.807745, 4.80905, 4.813972, 
    4.822018,
  // height(21,10, 0-49)
    4.882683, 4.887622, 4.893283, 4.899419, 4.905817, 4.912298, 4.918719, 
    4.924973, 4.930984, 4.936702, 4.942099, 4.947176, 4.951952, 4.956465, 
    4.960778, 4.962388, 4.966177, 4.968843, 4.970945, 4.972705, 4.974249, 
    4.977313, 4.979748, 4.98192, 4.984013, 4.985978, 4.98778, 4.989291, 
    4.99031, 4.990362, 4.988803, 4.987789, 4.985182, 4.980694, 4.97406, 
    4.965057, 4.953567, 4.939633, 4.923513, 4.905717, 4.887003, 4.868331, 
    4.85077, 4.835371, 4.823044, 4.814457, 4.809978, 4.809673, 4.813326, 
    4.820508,
  // height(21,11, 0-49)
    4.885859, 4.890782, 4.896351, 4.902331, 4.90852, 4.914749, 4.920887, 
    4.926834, 4.932517, 4.937896, 4.942946, 4.947676, 4.952104, 4.956275, 
    4.960248, 4.961854, 4.964558, 4.966954, 4.968882, 4.970501, 4.971934, 
    4.974759, 4.977002, 4.979015, 4.981116, 4.983275, 4.985504, 4.987677, 
    4.989609, 4.990688, 4.990268, 4.990361, 4.989007, 4.985883, 4.980674, 
    4.973091, 4.962924, 4.950112, 4.934801, 4.917403, 4.898602, 4.879333, 
    4.860695, 4.843828, 4.829777, 4.819361, 4.813109, 4.811215, 4.813574, 
    4.819819,
  // height(21,12, 0-49)
    4.88944, 4.894337, 4.899799, 4.905598, 4.911548, 4.917494, 4.923313, 
    4.928915, 4.934238, 4.939242, 4.943916, 4.948267, 4.952316, 4.956103, 
    4.959673, 4.961469, 4.963051, 4.965169, 4.966954, 4.968485, 4.96986, 
    4.972414, 4.974438, 4.976257, 4.978319, 4.980617, 4.983204, 4.985958, 
    4.988717, 4.990734, 4.99138, 4.99241, 4.992143, 4.990234, 4.986331, 
    4.980086, 4.971216, 4.959564, 4.945173, 4.928348, 4.909691, 4.890091, 
    4.870652, 4.852578, 4.837027, 4.824958, 4.81705, 4.813632, 4.814701, 
    4.819964,
  // height(21,13, 0-49)
    4.893345, 4.898217, 4.90356, 4.909164, 4.914856, 4.920492, 4.925966, 
    4.931196, 4.936131, 4.94074, 4.945012, 4.948959, 4.952602, 4.955966, 
    4.959073, 4.961245, 4.961709, 4.963559, 4.96524, 4.96674, 4.96812, 
    4.970376, 4.972166, 4.973768, 4.975757, 4.978142, 4.981021, 4.984272, 
    4.987758, 4.990619, 4.99226, 4.994047, 4.99469, 4.993832, 4.991089, 
    4.98607, 4.978432, 4.967936, 4.954527, 4.93841, 4.920095, 4.900408, 
    4.880437, 4.861424, 4.844614, 4.831095, 4.821679, 4.816827, 4.816639, 
    4.820898,
  // height(21,14, 0-49)
    4.897468, 4.902321, 4.907547, 4.912951, 4.918373, 4.923688, 4.928799, 
    4.93364, 4.93817, 4.942365, 4.946223, 4.949754, 4.95297, 4.95588, 
    4.958479, 4.961169, 4.960548, 4.962161, 4.963795, 4.965333, 4.966787, 
    4.968728, 4.97028, 4.971656, 4.973548, 4.975982, 4.979085, 4.982744, 
    4.986854, 4.990458, 4.993018, 4.995389, 4.996763, 4.99678, 4.995036, 
    4.991111, 4.98461, 4.975227, 4.962822, 4.947505, 4.929689, 4.910128, 
    4.889874, 4.870183, 4.852361, 4.837605, 4.826849, 4.820671, 4.819281, 
    4.822535,
  // height(21,15, 0-49)
    4.901683, 4.906533, 4.911652, 4.916859, 4.922011, 4.927, 4.931743, 
    4.936191, 4.94031, 4.944088, 4.94753, 4.950641, 4.953424, 4.955871, 
    4.957943, 4.96121, 4.959546, 4.960984, 4.962644, 4.9643, 4.965909, 
    4.967529, 4.968853, 4.970014, 4.971802, 4.974249, 4.977513, 4.981489, 
    4.986113, 4.990354, 4.993762, 4.996544, 4.998473, 4.999189, 4.998278, 
    4.995298, 4.989818, 4.981478, 4.970063, 4.955593, 4.938392, 4.919131, 
    4.898813, 4.878683, 4.860091, 4.844313, 4.832389, 4.825014, 4.822492, 
    4.824755,
  // height(21,16, 0-49)
    4.905852, 4.910719, 4.915746, 4.92077, 4.925663, 4.930331, 4.934713, 
    4.938773, 4.942492, 4.945868, 4.948905, 4.951612, 4.953979, 4.955981, 
    4.95755, 4.961321, 4.958642, 4.960001, 4.961782, 4.963653, 4.965511, 
    4.966817, 4.967943, 4.968918, 4.970611, 4.973051, 4.976418, 4.980618, 
    4.985636, 4.9904, 4.994579, 4.99761, 4.999923, 5.001165, 5.00092, 
    4.99873, 4.994142, 4.986749, 4.976277, 4.962667, 4.946156, 4.927331, 
    4.907132, 4.886779, 4.86764, 4.851046, 4.838132, 4.82969, 4.826118, 
    4.82742,
  // height(21,17, 0-49)
    4.909837, 4.914738, 4.919692, 4.924548, 4.929195, 4.93356, 4.9376, 
    4.941293, 4.944641, 4.947648, 4.950324, 4.95267, 4.954671, 4.956281, 
    4.957415, 4.961463, 4.957752, 4.959157, 4.961174, 4.963372, 4.965584, 
    4.966605, 4.967587, 4.968428, 4.970053, 4.97248, 4.975895, 4.980227, 
    4.985517, 4.99068, 4.995541, 4.998661, 5.001194, 5.002797, 5.003052, 
    5.001498, 4.997662, 4.991107, 4.98151, 4.968741, 4.95296, 4.934667, 
    4.914736, 4.894343, 4.874856, 4.857644, 4.843911, 4.834536, 4.83, 4.830382,
  // height(21,18, 0-49)
    4.913497, 4.918441, 4.923331, 4.928032, 4.932451, 4.936535, 4.940263, 
    4.943635, 4.946665, 4.949371, 4.951762, 4.953833, 4.955557, 4.956873, 
    4.957686, 4.961622, 4.956789, 4.958377, 4.96076, 4.963412, 4.9661, 
    4.966885, 4.967799, 4.968584, 4.970194, 4.972615, 4.97604, 4.980412, 
    4.985839, 4.991264, 4.996696, 4.999753, 5.002348, 5.004149, 5.004743, 
    5.003669, 5.000443, 4.994608, 4.985798, 4.973829, 4.958785, 4.94109, 
    4.921543, 4.901266, 4.881607, 4.863956, 4.849568, 4.839391, 4.833985, 
    4.833497,
  // height(21,19, 0-49)
    4.9167, 4.921665, 4.926477, 4.931019, 4.93522, 4.939054, 4.942522, 
    4.945646, 4.948455, 4.950972, 4.953205, 4.955136, 4.956722, 4.957885, 
    4.958528, 4.961836, 4.95568, 4.957586, 4.960464, 4.963702, 4.967002, 
    4.967633, 4.968585, 4.96942, 4.971097, 4.973547, 4.976954, 4.981276, 
    4.986701, 4.992226, 4.998084, 5.00092, 5.003414, 5.00525, 5.006023, 
    5.005275, 5.00252, 4.997281, 4.989166, 4.977938, 4.963619, 4.94656, 
    4.927482, 4.90745, 4.887774, 4.869849, 4.854956, 4.84411, 4.837931, 
    4.836633,
  // height(21,20, 0-49)
    4.920373, 4.926408, 4.932198, 4.937615, 4.942574, 4.947017, 4.95092, 
    4.954266, 4.957061, 4.959322, 4.961086, 4.962402, 4.963344, 4.963996, 
    4.96446, 0, 4.958336, 4.959911, 4.962055, 4.964373, 4.966731, 4.965669, 
    4.965298, 4.965133, 4.966242, 4.968559, 4.972223, 4.977122, 4.983384, 
    4.989923, 4.997092, 5.000469, 5.003476, 5.005798, 5.007044, 5.006776, 
    5.004527, 4.999839, 4.992319, 4.981717, 4.96802, 4.951524, 4.932887, 
    4.913119, 4.893489, 4.875374, 4.860076, 4.848648, 4.841766, 4.839701,
  // height(21,21, 0-49)
    4.922716, 4.928973, 4.934875, 4.9403, 4.945176, 4.949471, 4.95318, 
    4.956317, 4.958914, 4.96101, 4.962654, 4.963908, 4.964848, 4.965567, 
    4.966182, 0, 4.955145, 4.957202, 4.959885, 4.962759, 4.965636, 4.964164, 
    4.963536, 4.963161, 4.964198, 4.966575, 4.970424, 4.975614, 4.982278, 
    4.989311, 4.997245, 5.000715, 5.003937, 5.006592, 5.008276, 5.008539, 
    5.006902, 5.002893, 4.996096, 4.986228, 4.97323, 4.957343, 4.939162, 
    4.919639, 4.900001, 4.881614, 4.865797, 4.85364, 4.845881, 4.842846,
  // height(21,22, 0-49)
    4.924577, 4.931123, 4.937216, 4.942735, 4.947618, 4.951845, 4.955435, 
    4.958422, 4.960857, 4.962803, 4.964324, 4.965492, 4.966395, 4.967139, 
    4.967857, 0, 4.952854, 4.955309, 4.958461, 4.96184, 4.965202, 4.963355, 
    4.962503, 4.961944, 4.962914, 4.96533, 4.96931, 4.974701, 4.981636, 
    4.988995, 4.997468, 5.000855, 5.004099, 5.006884, 5.008801, 5.009401, 
    5.008202, 5.004722, 4.998529, 4.989316, 4.976982, 4.961714, 4.944051, 
    4.92488, 4.905382, 4.886895, 4.870741, 4.858034, 4.849556, 4.845685,
  // height(21,23, 0-49)
    4.925975, 4.932854, 4.939191, 4.944864, 4.949818, 4.954044, 4.957575, 
    4.960462, 4.962778, 4.964598, 4.966004, 4.967083, 4.967932, 4.968668, 
    4.969452, 0, 4.951511, 4.954235, 4.957705, 4.961428, 4.965119, 4.962908, 
    4.961822, 4.961064, 4.961936, 4.964339, 4.968385, 4.973899, 4.98101, 
    4.988581, 4.997424, 5.000678, 5.003872, 5.006702, 5.008762, 5.009603, 
    5.008744, 5.0057, 5.000029, 4.9914, 4.97968, 4.96501, 4.947873, 4.929098, 
    4.909818, 4.891339, 4.874972, 4.861847, 4.852779, 4.848183,
  // height(21,24, 0-49)
    4.926955, 4.934186, 4.940796, 4.946662, 4.951729, 4.956, 4.959518, 
    4.962349, 4.964579, 4.966302, 4.96761, 4.968601, 4.969385, 4.970094, 
    4.970906, 0, 4.951337, 4.954191, 4.957818, 4.961719, 4.965586, 4.963124, 
    4.961879, 4.96099, 4.961792, 4.964177, 4.968248, 4.973822, 4.981027, 
    4.988714, 4.997774, 5.000921, 5.004061, 5.006891, 5.009009, 5.009973, 
    5.009304, 5.006517, 5.001168, 4.992916, 4.981607, 4.967354, 4.950599, 
    4.932136, 4.913054, 4.894632, 4.878164, 4.864782, 4.855316, 4.850201,
  // height(21,25, 0-49)
    4.927581, 4.93516, 4.94205, 4.948121, 4.953326, 4.957671, 4.961206, 
    4.964014, 4.96619, 4.967835, 4.969058, 4.969966, 4.970678, 4.971337, 
    4.972132, 0, 4.951993, 4.954841, 4.958466, 4.962369, 4.966248, 4.963695, 
    4.962402, 4.961487, 4.962284, 4.964675, 4.968763, 4.974359, 4.981592, 
    4.989312, 4.998431, 5.001542, 5.004662, 5.007491, 5.009628, 5.010636, 
    5.010038, 5.007354, 5.002141, 4.994059, 4.982945, 4.968903, 4.952358, 
    4.934081, 4.915137, 4.896785, 4.880301, 4.866809, 4.857136, 4.851721,
  // height(21,26, 0-49)
    4.927925, 4.935825, 4.942978, 4.949254, 4.954605, 4.959037, 4.962613, 
    4.965418, 4.967557, 4.969142, 4.970285, 4.971105, 4.971728, 4.972306, 
    4.973034, 0, 4.953425, 4.95613, 4.959591, 4.963326, 4.96705, 4.964577, 
    4.963362, 4.962536, 4.963402, 4.965837, 4.969944, 4.975535, 4.982742, 
    4.990416, 4.999442, 5.002605, 5.005761, 5.008602, 5.010732, 5.011711, 
    5.011069, 5.008329, 5.003057, 4.994917, 4.983764, 4.969701, 4.953165, 
    4.934923, 4.91604, 4.89776, 4.881342, 4.867894, 4.858222, 4.852753,
  // height(21,27, 0-49)
    4.92806, 4.936237, 4.943624, 4.950087, 4.955577, 4.960105, 4.963733, 
    4.96655, 4.968665, 4.970191, 4.971249, 4.971961, 4.972464, 4.972912, 
    4.973501, 0, 4.955719, 4.958138, 4.961273, 4.964661, 4.968061, 4.965804, 
    4.964757, 4.964105, 4.965088, 4.967585, 4.971696, 4.977244, 4.98436, 
    4.99191, 5.000689, 5.003982, 5.007212, 5.01007, 5.012156, 5.013031, 
    5.01223, 5.009284, 5.00377, 4.995371, 4.983961, 4.969677, 4.952976, 
    4.93465, 4.915774, 4.897588, 4.881337, 4.868097, 4.85864, 4.853362,
  // height(21,28, 0-49)
    4.928054, 4.936454, 4.944035, 4.950661, 4.956285, 4.960913, 4.964603, 
    4.967442, 4.969531, 4.970989, 4.971935, 4.972499, 4.972823, 4.973068, 
    4.973427, 0, 4.959241, 4.961226, 4.963868, 4.966732, 4.969642, 4.967668, 
    4.96682, 4.966366, 4.967466, 4.969997, 4.974066, 4.979512, 4.986459, 
    4.993795, 5.002191, 5.005653, 5.008963, 5.011804, 5.013775, 5.014439, 
    5.013337, 5.010012, 5.004061, 4.995199, 4.983335, 4.968651, 4.951647, 
    4.933157, 4.914279, 4.896254, 4.880302, 4.867464, 4.858457, 4.853627,
  // height(21,29, 0-49)
    4.92797, 4.936532, 4.944271, 4.951048, 4.956806, 4.961545, 4.965309, 
    4.968172, 4.970227, 4.971584, 4.972364, 4.972703, 4.972755, 4.972694, 
    4.972711, 0, 4.963769, 4.965175, 4.967158, 4.969325, 4.971568, 4.96982, 
    4.969094, 4.968768, 4.969911, 4.972406, 4.976363, 4.981632, 4.988328, 
    4.995357, 5.003223, 5.006826, 5.010169, 5.01293, 5.014711, 5.015079, 
    5.013591, 5.0098, 5.003335, 4.99394, 4.981572, 4.966462, 4.949168, 
    4.930563, 4.911772, 4.894035, 4.878546, 4.866288, 4.85792, 4.853728,
  // height(21,30, 0-49)
    4.926956, 4.934618, 4.941468, 4.947391, 4.952364, 4.956439, 4.959708, 
    4.962296, 4.964333, 4.965935, 4.967184, 4.968123, 4.968738, 4.968968, 
    4.968709, 4.975595, 4.962874, 4.964472, 4.967275, 4.970613, 4.974156, 
    4.97453, 4.975579, 4.976661, 4.978667, 4.98145, 4.985137, 4.989669, 
    4.995262, 5.000958, 5.007199, 5.009936, 5.012409, 5.014312, 5.015257, 
    5.014821, 5.012557, 5.008026, 5.000863, 4.990838, 4.977942, 4.962452, 
    4.944969, 4.926406, 4.9079, 4.890683, 4.875904, 4.864484, 4.857009, 
    4.853695,
  // height(21,31, 0-49)
    4.926929, 4.934672, 4.941601, 4.947601, 4.95264, 4.956754, 4.960025, 
    4.962573, 4.964523, 4.965997, 4.967094, 4.96788, 4.968374, 4.968542, 
    4.968293, 4.975252, 4.964764, 4.96593, 4.968161, 4.970851, 4.97374, 
    4.974269, 4.975286, 4.976324, 4.978278, 4.981052, 4.98479, 4.98941, 
    4.995051, 5.0007, 5.006574, 5.009628, 5.012319, 5.014328, 5.015259, 
    5.014685, 5.012158, 5.007254, 4.999632, 4.989102, 4.975713, 4.959807, 
    4.942053, 4.923415, 4.905064, 4.888221, 4.874006, 4.863276, 4.856546, 
    4.853962,
  // height(21,32, 0-49)
    4.926838, 4.934477, 4.941327, 4.947276, 4.952287, 4.956389, 4.959658, 
    4.962198, 4.964133, 4.965584, 4.966657, 4.967435, 4.967957, 4.968214, 
    4.968139, 4.974419, 4.966065, 4.966943, 4.968725, 4.970888, 4.973237, 
    4.974019, 4.975111, 4.976216, 4.978195, 4.980991, 4.984751, 4.989377, 
    4.994931, 5.000389, 5.005764, 5.009021, 5.011818, 5.013818, 5.014621, 
    5.013795, 5.0109, 5.005525, 4.997361, 4.986272, 4.972367, 4.956063, 
    4.938097, 4.919488, 4.901426, 4.885119, 4.871639, 4.861775, 4.855964, 
    4.854273,
  // height(21,33, 0-49)
    4.926754, 4.934147, 4.940796, 4.946594, 4.951506, 4.955551, 4.958797, 
    4.961343, 4.963299, 4.964785, 4.96591, 4.966764, 4.967407, 4.967854, 
    4.968068, 4.973201, 4.966861, 4.967598, 4.969047, 4.970792, 4.972705, 
    4.973806, 4.97506, 4.976316, 4.978374, 4.981203, 4.984944, 4.989483, 
    4.994825, 4.999962, 5.004738, 5.008092, 5.010881, 5.012757, 5.013318, 
    5.012129, 5.00876, 5.002823, 4.994051, 4.982362, 4.967942, 4.951282, 
    4.93319, 4.914731, 4.897108, 4.881502, 4.868926, 4.86009, 4.855348, 
    4.854691,
  // height(21,34, 0-49)
    4.926736, 4.933774, 4.940129, 4.945702, 4.950455, 4.954404, 4.95761, 
    4.960158, 4.962151, 4.9637, 4.964916, 4.96589, 4.966699, 4.967385, 
    4.967942, 4.971733, 4.967276, 4.967985, 4.969195, 4.970612, 4.972173, 
    4.973621, 4.975093, 4.976563, 4.978733, 4.98159, 4.98526, 4.989622, 
    4.994627, 4.999331, 5.003438, 5.006778, 5.009446, 5.011085, 5.011292, 
    5.009635, 5.005699, 4.999127, 4.989699, 4.977401, 4.962496, 4.945557, 
    4.927455, 4.909292, 4.892269, 4.877531, 4.866017, 4.858353, 4.854806, 
    4.855289,
  // height(21,35, 0-49)
    4.926836, 4.933433, 4.939422, 4.944709, 4.949258, 4.953081, 4.956228, 
    4.95877, 4.960804, 4.96243, 4.96375, 4.964861, 4.965849, 4.966776, 
    4.967676, 4.970145, 4.967444, 4.968202, 4.969242, 4.970393, 4.971665, 
    4.973465, 4.975183, 4.976903, 4.979197, 4.982062, 4.985603, 4.989695, 
    4.994246, 4.998414, 5.001794, 5.005006, 5.007436, 5.008721, 5.008463, 
    5.00624, 5.001657, 4.994396, 4.984295, 4.971416, 4.9561, 4.938995, 
    4.921033, 4.903339, 4.887095, 4.873391, 4.863085, 4.856715, 4.854457, 
    4.856152,
  // height(21,36, 0-49)
    4.927101, 4.933189, 4.938755, 4.943709, 4.948019, 4.951687, 4.954755, 
    4.957284, 4.959356, 4.961058, 4.962487, 4.963735, 4.964891, 4.966037, 
    4.967238, 4.96855, 4.967488, 4.968328, 4.969235, 4.970166, 4.9712, 
    4.973329, 4.975299, 4.977283, 4.979695, 4.982537, 4.985882, 4.989611, 
    4.993591, 4.997127, 4.999732, 5.00269, 5.004757, 5.005571, 5.00474, 
    5.00186, 4.996566, 4.988592, 4.977838, 4.964443, 4.948833, 4.931724, 
    4.91409, 4.897061, 4.881786, 4.869282, 4.860319, 4.855337, 4.85443, 
    4.857368,
  // height(21,37, 0-49)
    4.927572, 4.933101, 4.938197, 4.942782, 4.946818, 4.950309, 4.95328, 
    4.955783, 4.957885, 4.959661, 4.961193, 4.962566, 4.963869, 4.965193, 
    4.966624, 4.967034, 4.967501, 4.96842, 4.969209, 4.969953, 4.970782, 
    4.9732, 4.975408, 4.97765, 4.980156, 4.982931, 4.986008, 4.989279, 
    4.992575, 4.995385, 4.997163, 4.999734, 5.00131, 5.001532, 5.000024, 
    4.996412, 4.990367, 4.981685, 4.970336, 4.956542, 4.940803, 4.923894, 
    4.906811, 4.890669, 4.876559, 4.865418, 4.857912, 4.854388, 4.854856, 
    4.859026,
  // height(21,38, 0-49)
    4.928286, 4.933214, 4.937806, 4.941989, 4.945725, 4.949013, 4.951869, 
    4.954332, 4.956453, 4.95829, 4.959915, 4.9614, 4.962823, 4.964279, 
    4.965862, 4.965644, 4.967535, 4.968503, 4.969175, 4.969752, 4.970407, 
    4.97306, 4.975472, 4.977946, 4.980508, 4.983161, 4.985892, 4.988606, 
    4.991111, 4.993099, 4.993998, 4.996039, 4.99699, 4.996502, 4.994226, 
    4.989821, 4.983016, 4.97367, 4.961834, 4.947803, 4.932146, 4.915679, 
    4.899399, 4.884381, 4.87164, 4.86201, 4.856055, 4.854027, 4.85586, 
    4.861211,
  // height(21,39, 0-49)
    4.929265, 4.933565, 4.937625, 4.941379, 4.944791, 4.947852, 4.950571, 
    4.952974, 4.955095, 4.95698, 4.958681, 4.960257, 4.961775, 4.963317, 
    4.964976, 4.964395, 4.967595, 4.96857, 4.969121, 4.969549, 4.97005, 
    4.972878, 4.975447, 4.978108, 4.980676, 4.983141, 4.985444, 4.987503, 
    4.989108, 4.990186, 4.990143, 4.991511, 4.991702, 4.990395, 4.987274, 
    4.982047, 4.974504, 4.964581, 4.952405, 4.938348, 4.923028, 4.907279, 
    4.892075, 4.878423, 4.867244, 4.859259, 4.854925, 4.8544, 4.857553, 
    4.863996,
  // height(21,40, 0-49)
    4.930509, 4.934163, 4.937672, 4.940976, 4.944041, 4.946851, 4.949409, 
    4.951728, 4.953829, 4.95574, 4.957498, 4.959143, 4.96073, 4.962318, 
    4.963991, 4.96327, 4.967656, 4.968591, 4.969017, 4.969309, 4.969671, 
    4.972606, 4.975278, 4.97807, 4.980577, 4.982781, 4.984569, 4.985875, 
    4.986485, 4.986562, 4.985514, 4.986065, 4.985376, 4.983157, 4.979137, 
    4.973087, 4.964869, 4.954496, 4.942178, 4.928343, 4.913644, 4.898909, 
    4.885057, 4.873009, 4.86357, 4.857339, 4.854666, 4.855622, 4.860014, 
    4.867422,
  // height(21,41, 0-49)
    4.931998, 4.934996, 4.937942, 4.94078, 4.943478, 4.946014, 4.948385, 
    4.950592, 4.952645, 4.954556, 4.956345, 4.958038, 4.959667, 4.961271, 
    4.962908, 4.962221, 4.967657, 4.968509, 4.968806, 4.968975, 4.969211, 
    4.972187, 4.974899, 4.977754, 4.980126, 4.981987, 4.983173, 4.983639, 
    4.983162, 4.982157, 4.980039, 4.979643, 4.977969, 4.974769, 4.969831, 
    4.962996, 4.954207, 4.943558, 4.931327, 4.917993, 4.904217, 4.890792, 
    4.878562, 4.868335, 4.860787, 4.856392, 4.855388, 4.857768, 4.863286, 
    4.8715,
  // height(21,42, 0-49)
    4.933681, 4.93602, 4.938399, 4.940762, 4.943074, 4.945315, 4.947473, 
    4.949539, 4.951512, 4.953393, 4.955186, 4.9569, 4.958545, 4.960138, 
    4.961708, 4.961169, 4.967508, 4.968248, 4.968419, 4.968473, 4.968589, 
    4.971543, 4.97423, 4.977072, 4.979232, 4.980669, 4.981169, 4.980713, 
    4.979079, 4.976922, 4.973677, 4.972228, 4.969491, 4.965276, 4.95944, 
    4.951901, 4.942686, 4.931967, 4.920083, 4.907539, 4.894986, 4.883152, 
    4.872786, 4.864562, 4.859018, 4.856503, 4.857143, 4.860859, 4.867363, 
    4.876194,
  // height(21,43, 0-49)
    4.935478, 4.937166, 4.938977, 4.940857, 4.942774, 4.9447, 4.946618, 
    4.948514, 4.950376, 4.952195, 4.953959, 4.955664, 4.957301, 4.958864, 
    4.960346, 4.960024, 4.967107, 4.967718, 4.967767, 4.967717, 4.967713, 
    4.970584, 4.973182, 4.975931, 4.977798, 4.978734, 4.978477, 4.977031, 
    4.974191, 4.970835, 4.966425, 4.963848, 4.960012, 4.95479, 4.948117, 
    4.939998, 4.930539, 4.919984, 4.908716, 4.897247, 4.886191, 4.876195, 
    4.867887, 4.861801, 4.858331, 4.857696, 4.859924, 4.86486, 4.87218, 
    4.88142,
  // height(21,44, 0-49)
    4.937275, 4.938323, 4.939574, 4.940974, 4.942487, 4.944084, 4.945742, 
    4.947441, 4.949162, 4.950884, 4.95259, 4.954257, 4.955863, 4.957377, 
    4.958764, 4.958681, 4.966344, 4.966816, 4.966756, 4.966607, 4.966479, 
    4.969213, 4.971659, 4.974236, 4.975735, 4.976098, 4.975027, 4.972552, 
    4.968484, 4.96391, 4.958328, 4.954591, 4.949665, 4.943493, 4.936093, 
    4.927554, 4.91806, 4.907915, 4.897525, 4.887393, 4.878069, 4.8701, 
    4.863985, 4.860114, 4.858732, 4.859934, 4.863651, 4.869663, 4.877614, 
    4.887039,
  // height(21,45, 0-49)
    4.938926, 4.939353, 4.940056, 4.940982, 4.942094, 4.943354, 4.944736, 
    4.946219, 4.947771, 4.949369, 4.950988, 4.952592, 4.954145, 4.955598, 
    4.956888, 4.957033, 4.965114, 4.965453, 4.965286, 4.965036, 4.964778, 
    4.967328, 4.969562, 4.97189, 4.972956, 4.972693, 4.970773, 4.967258, 
    4.961981, 4.956205, 4.949481, 4.944608, 4.938652, 4.931637, 4.923662, 
    4.914896, 4.905593, 4.896097, 4.886826, 4.878241, 4.870824, 4.865007, 
    4.861149, 4.859497, 4.860159, 4.863107, 4.868181, 4.875099, 4.883481, 
    4.892863,
  // height(21,46, 0-49)
    4.940262, 4.940084, 4.940259, 4.940728, 4.941444, 4.942371, 4.943476, 
    4.944729, 4.946098, 4.947554, 4.949063, 4.950583, 4.952066, 4.953447, 
    4.954642, 4.95498, 4.963323, 4.963535, 4.963268, 4.96291, 4.962506, 
    4.964828, 4.9668, 4.968812, 4.969393, 4.968471, 4.965699, 4.961167, 
    4.954741, 4.947829, 4.940039, 4.934107, 4.927235, 4.919528, 4.911165, 
    4.902386, 4.893498, 4.884871, 4.876911, 4.870032, 4.864622, 4.861, 
    4.859388, 4.859892, 4.862491, 4.867044, 4.873307, 4.880941, 4.889546, 
    4.898666,
  // height(21,47, 0-49)
    4.941096, 4.940332, 4.939998, 4.940029, 4.940372, 4.940979, 4.941815, 
    4.942842, 4.944026, 4.945332, 4.94672, 4.948144, 4.949549, 4.950854, 
    4.951961, 4.952435, 4.960899, 4.960996, 4.960621, 4.960141, 4.959572, 
    4.961631, 4.963296, 4.964937, 4.965001, 4.963412, 4.959817, 4.954334, 
    4.946867, 4.938931, 4.930195, 4.923338, 4.915718, 4.907512, 4.898972, 
    4.890397, 4.882132, 4.874554, 4.868045, 4.862955, 4.859578, 4.858113, 
    4.858655, 4.861183, 4.865554, 4.871528, 4.878778, 4.886925, 4.895541, 
    4.904192,
  // height(21,48, 0-49)
    4.941243, 4.939906, 4.939085, 4.938703, 4.938699, 4.939013, 4.939602, 
    4.940422, 4.941435, 4.942599, 4.943874, 4.945204, 4.946529, 4.947761, 
    4.948786, 4.949333, 4.957789, 4.957774, 4.957283, 4.956659, 4.955901, 
    4.95767, 4.958993, 4.960226, 4.959764, 4.95753, 4.953178, 4.946849, 
    4.938492, 4.929691, 4.920184, 4.91259, 4.904428, 4.895942, 4.887444, 
    4.879278, 4.871814, 4.865419, 4.860435, 4.857142, 4.855741, 4.856319, 
    4.858856, 4.863209, 4.869135, 4.876301, 4.884318, 4.892757, 4.901187, 
    4.909195,
  // height(21,49, 0-49)
    4.941844, 4.93949, 4.937799, 4.936679, 4.936049, 4.935833, 4.935967, 
    4.936391, 4.937048, 4.937884, 4.938838, 4.939832, 4.94078, 4.941552, 
    4.941981, 4.941836, 4.957452, 4.955976, 4.953788, 4.951624, 4.94955, 
    4.952877, 4.955788, 4.959049, 4.959525, 4.957204, 4.951482, 4.942688, 
    4.930685, 4.918662, 4.906098, 4.898111, 4.889776, 4.881432, 4.873471, 
    4.866293, 4.860284, 4.855782, 4.853061, 4.852297, 4.853556, 4.856781, 
    4.861804, 4.868344, 4.876037, 4.88445, 4.893135, 4.901632, 4.909525, 
    4.916467,
  // height(22,0, 0-49)
    4.880537, 4.886049, 4.892055, 4.89834, 4.90474, 4.911143, 4.917471, 
    4.923685, 4.92976, 4.935697, 4.941501, 4.947173, 4.952713, 4.958113, 
    4.963342, 4.968148, 4.973527, 4.977929, 4.981947, 4.985516, 4.988526, 
    4.991129, 4.992905, 4.993828, 4.99375, 4.992583, 4.990228, 4.986621, 
    4.981689, 4.975449, 4.967793, 4.959002, 4.948776, 4.937156, 4.924249, 
    4.910238, 4.895406, 4.880136, 4.864914, 4.850298, 4.836879, 4.825234, 
    4.815861, 4.809134, 4.805259, 4.804258, 4.805966, 4.810053, 4.816054, 
    4.823408,
  // height(22,1, 0-49)
    4.881404, 4.887128, 4.893311, 4.899741, 4.906262, 4.912758, 4.919157, 
    4.925417, 4.93152, 4.937462, 4.943248, 4.948881, 4.954358, 4.959669, 
    4.964782, 4.969224, 4.975, 4.979175, 4.982958, 4.986339, 4.989226, 
    4.992044, 4.994077, 4.995368, 4.995728, 4.995061, 4.993247, 4.99022, 
    4.985889, 4.980306, 4.973286, 4.96537, 4.95594, 4.94499, 4.932577, 
    4.918843, 4.904028, 4.888497, 4.872729, 4.857299, 4.842846, 4.830007, 
    4.819363, 4.81137, 4.806323, 4.804312, 4.805237, 4.808805, 4.814574, 
    4.821985,
  // height(22,2, 0-49)
    4.882138, 4.888039, 4.894367, 4.900916, 4.907531, 4.914097, 4.920544, 
    4.926829, 4.932936, 4.938857, 4.944596, 4.950159, 4.955542, 4.960733, 
    4.965704, 4.969741, 4.975807, 4.979735, 4.983255, 4.986413, 4.989146, 
    4.992136, 4.994386, 4.996001, 4.99677, 4.996595, 4.995338, 4.992937, 
    4.989284, 4.984453, 4.978187, 4.971295, 4.962846, 4.952787, 4.941124, 
    4.927945, 4.913436, 4.897918, 4.881842, 4.865784, 4.850403, 4.836392, 
    4.824409, 4.815003, 4.808563, 4.805276, 4.805117, 4.807853, 4.813084, 
    4.820271,
  // height(22,3, 0-49)
    4.88286, 4.888899, 4.895341, 4.901977, 4.908658, 4.915267, 4.921736, 
    4.92802, 4.9341, 4.93997, 4.945633, 4.951095, 4.956351, 4.961398, 
    4.966206, 4.969803, 4.976026, 4.979697, 4.982938, 4.98585, 4.988398, 
    4.991513, 4.99393, 4.995817, 4.996953, 4.997241, 4.996539, 4.994784, 
    4.991858, 4.987838, 4.982406, 4.976634, 4.969298, 4.960302, 4.949604, 
    4.937222, 4.923286, 4.908053, 4.891929, 4.875461, 4.859316, 4.844221, 
    4.830904, 4.820007, 4.812023, 4.807248, 4.80575, 4.807377, 4.811787, 
    4.818478,
  // height(22,4, 0-49)
    4.883684, 4.889828, 4.896346, 4.903038, 4.90975, 4.916372, 4.922831, 
    4.929082, 4.935105, 4.940893, 4.946448, 4.951777, 4.956883, 4.96176, 
    4.966392, 4.969527, 4.975749, 4.97916, 4.982116, 4.984766, 4.987107, 
    4.990293, 4.992825, 4.99492, 4.996367, 4.997078, 4.996912, 4.995807, 
    4.993631, 4.990452, 4.985897, 4.981287, 4.975144, 4.96733, 4.957751, 
    4.94637, 4.93324, 4.918549, 4.902637, 4.886006, 4.869302, 4.853272, 
    4.838696, 4.826305, 4.8167, 4.810288, 4.807254, 4.807538, 4.810874, 
    4.816814,
  // height(22,5, 0-49)
    4.884719, 4.890928, 4.897486, 4.904196, 4.910906, 4.917505, 4.92392, 
    4.930103, 4.936036, 4.941709, 4.947129, 4.952298, 4.957226, 4.961914, 
    4.96636, 4.969028, 4.97508, 4.978233, 4.980904, 4.983284, 4.985404, 
    4.98861, 4.991196, 4.993429, 4.995127, 4.99621, 4.996547, 4.996074, 
    4.994657, 4.992321, 4.988653, 4.985206, 4.980282, 4.973714, 4.96536, 
    4.955123, 4.942988, 4.929064, 4.913613, 4.897071, 4.880046, 4.86328, 
    4.847586, 4.833769, 4.822536, 4.814412, 4.809701, 4.80846, 4.81051, 
    4.815478,
  // height(22,6, 0-49)
    4.886049, 4.892287, 4.898846, 4.905535, 4.912204, 4.918742, 4.925076, 
    4.931158, 4.936968, 4.942498, 4.947752, 4.952737, 4.957466, 4.961949, 
    4.9662, 4.968412, 4.974121, 4.97702, 4.979414, 4.981527, 4.983417, 
    4.986587, 4.98917, 4.991468, 4.99335, 4.994747, 4.995544, 4.99568, 
    4.995009, 4.993502, 4.990707, 4.988382, 4.984662, 4.979352, 4.972273, 
    4.963274, 4.952274, 4.9393, 4.924531, 4.908326, 4.89123, 4.873957, 
    4.857336, 4.842224, 4.829421, 4.819574, 4.813116, 4.810222, 4.810823, 
    4.814631,
  // height(22,7, 0-49)
    4.887733, 4.893962, 4.900485, 4.907114, 4.913703, 4.920143, 4.92636, 
    4.932308, 4.937963, 4.94332, 4.948382, 4.953161, 4.957674, 4.961939, 
    4.965983, 4.967781, 4.972977, 4.975623, 4.977752, 4.979605, 4.981266, 
    4.984348, 4.986871, 4.989161, 4.991158, 4.992808, 4.994019, 4.994727, 
    4.994781, 4.994075, 4.992127, 4.990852, 4.98828, 4.984199, 4.978396, 
    4.970678, 4.960901, 4.949014, 4.935112, 4.919465, 4.902544, 4.885012, 
    4.867685, 4.851458, 4.837206, 4.825689, 4.817468, 4.812854, 4.811893, 
    4.814398,
  // height(22,8, 0-49)
    4.88981, 4.895993, 4.902441, 4.908971, 4.915441, 4.921747, 4.927812, 
    4.933593, 4.939067, 4.944226, 4.949075, 4.953628, 4.957908, 4.96194, 
    4.965762, 4.967212, 4.971738, 4.974128, 4.976008, 4.977619, 4.979063, 
    4.982004, 4.98441, 4.986624, 4.988671, 4.990512, 4.992086, 4.993325, 
    4.994076, 4.994135, 4.992996, 4.992678, 4.991173, 4.988257, 4.983695, 
    4.977253, 4.968738, 4.958027, 4.945134, 4.930234, 4.913712, 4.896164, 
    4.878372, 4.86124, 4.845705, 4.832624, 4.822687, 4.816338, 4.813755, 
    4.814858,
  // height(22,9, 0-49)
    4.892284, 4.898389, 4.904727, 4.911123, 4.917439, 4.923574, 4.929457, 
    4.935043, 4.94031, 4.945249, 4.949864, 4.954177, 4.958208, 4.96199, 
    4.965567, 4.966765, 4.970487, 4.972616, 4.974267, 4.975658, 4.976905, 
    4.979655, 4.981893, 4.983966, 4.986002, 4.987977, 4.989863, 4.991588, 
    4.993001, 4.993782, 4.993412, 4.993945, 4.993408, 4.991569, 4.988178, 
    4.982973, 4.975715, 4.966225, 4.954433, 4.940427, 4.924498, 4.90716, 
    4.889142, 4.871335, 4.854712, 4.84022, 4.828661, 4.820616, 4.8164, 
    4.816047,
  // height(22,10, 0-49)
    4.895145, 4.901142, 4.907338, 4.913567, 4.919698, 4.925632, 4.931304, 
    4.93667, 4.941706, 4.946405, 4.950773, 4.95483, 4.958596, 4.96211, 
    4.965409, 4.96648, 4.969285, 4.971148, 4.972591, 4.973794, 4.974871, 
    4.977384, 4.979412, 4.981291, 4.983261, 4.985313, 4.987463, 4.989625, 
    4.991659, 4.993119, 4.993484, 4.99475, 4.995069, 4.994203, 4.991892, 
    4.987855, 4.981818, 4.973549, 4.96291, 4.949902, 4.93472, 4.917789, 
    4.899768, 4.881516, 4.864025, 4.8483, 4.835255, 4.825601, 4.819786, 
    4.817967,
  // height(22,11, 0-49)
    4.898359, 4.904222, 4.910252, 4.916286, 4.922204, 4.927913, 4.93335, 
    4.938472, 4.943258, 4.947702, 4.951809, 4.955594, 4.959082, 4.962301, 
    4.965283, 4.966367, 4.968176, 4.969769, 4.971031, 4.972083, 4.973031, 
    4.975266, 4.977045, 4.978685, 4.980544, 4.98263, 4.984991, 4.987542, 
    4.990149, 4.992247, 4.993314, 4.995196, 4.996253, 4.996246, 4.994911, 
    4.991952, 4.987071, 4.979993, 4.970516, 4.958566, 4.944244, 4.927882, 
    4.910058, 4.891582, 4.873441, 4.856687, 4.842321, 4.831179, 4.823837, 
    4.82058,
  // height(22,12, 0-49)
    4.901878, 4.907592, 4.913434, 4.919252, 4.924936, 4.930398, 4.935579, 
    4.940441, 4.944962, 4.949134, 4.952963, 4.956466, 4.959656, 4.962557, 
    4.965181, 4.966418, 4.967177, 4.968506, 4.96962, 4.970567, 4.97143, 
    4.973352, 4.974858, 4.976231, 4.977943, 4.980022, 4.98255, 4.985436, 
    4.988568, 4.991255, 4.992997, 4.995377, 4.997054, 4.99779, 4.997318, 
    4.995336, 4.991525, 4.98558, 4.977245, 4.966374, 4.952986, 4.937315, 
    4.919857, 4.901359, 4.882782, 4.865209, 4.849709, 4.837227, 4.828466, 
    4.823829,
  // height(22,13, 0-49)
    4.90565, 4.911202, 4.916841, 4.922431, 4.927863, 4.933063, 4.937972, 
    4.942556, 4.946795, 4.950685, 4.954226, 4.957429, 4.960305, 4.962861, 
    4.96509, 4.966601, 4.96628, 4.967366, 4.968375, 4.969272, 4.970106, 
    4.971691, 4.97291, 4.973999, 4.975545, 4.977583, 4.980232, 4.9834, 
    4.986999, 4.990225, 4.992621, 4.995386, 4.997564, 4.998925, 4.999202, 
    4.998087, 4.99525, 4.990359, 4.983118, 4.973319, 4.960899, 4.946009, 
    4.92905, 4.910706, 4.891897, 4.873711, 4.857275, 4.843622, 4.83357, 
    4.827637,
  // height(22,14, 0-49)
    4.909611, 4.915001, 4.920432, 4.925782, 4.930954, 4.935875, 4.940499, 
    4.944792, 4.948737, 4.952328, 4.955569, 4.958461, 4.961009, 4.963201, 
    4.965012, 4.966866, 4.965448, 4.966335, 4.967295, 4.968207, 4.969079, 
    4.970313, 4.971245, 4.97205, 4.973421, 4.975398, 4.978127, 4.981521, 
    4.985519, 4.989235, 4.992261, 4.995299, 4.997867, 4.999737, 5.000646, 
    5.000288, 4.998318, 4.994392, 4.988178, 4.979414, 4.96797, 4.953912, 
    4.937561, 4.919518, 4.900659, 4.882061, 4.864886, 4.850241, 4.839045, 
    4.831921,
  // height(22,15, 0-49)
    4.913706, 4.918937, 4.924161, 4.929266, 4.934164, 4.938797, 4.943122, 
    4.947111, 4.950749, 4.954034, 4.956963, 4.959537, 4.961747, 4.96357, 
    4.964959, 4.967154, 4.964622, 4.965373, 4.966358, 4.967362, 4.968349, 
    4.96923, 4.969894, 4.970437, 4.971638, 4.973541, 4.976313, 4.979875, 
    4.984203, 4.988347, 4.99198, 4.995186, 4.998031, 5.000298, 5.001725, 
    5.002008, 5.000802, 4.997742, 4.992472, 4.984691, 4.974206, 4.96101, 
    4.945339, 4.927721, 4.908974, 4.89015, 4.87243, 4.856977, 4.844789, 
    4.836594,
  // height(22,16, 0-49)
    4.917878, 4.922956, 4.927972, 4.932827, 4.937447, 4.94178, 4.945793, 
    4.949466, 4.952789, 4.95576, 4.958376, 4.960632, 4.962512, 4.963979, 
    4.964971, 4.967404, 4.963717, 4.964427, 4.965526, 4.966713, 4.967906, 
    4.968447, 4.96888, 4.969199, 4.970256, 4.972084, 4.974867, 4.978536, 
    4.983116, 4.987617, 4.991826, 4.995096, 4.998113, 5.000667, 5.002501, 
    5.003314, 5.00276, 5.000465, 4.996054, 4.989187, 4.979626, 4.967295, 
    4.952357, 4.935261, 4.916767, 4.897888, 4.879806, 4.863722, 4.850706, 
    4.841565,
  // height(22,17, 0-49)
    4.92207, 4.926999, 4.931807, 4.936404, 4.940733, 4.944755, 4.948444, 
    4.951794, 4.9548, 4.957461, 4.959776, 4.961733, 4.963308, 4.964456, 
    4.965109, 4.967572, 4.962652, 4.963425, 4.964743, 4.966219, 4.967717, 
    4.967952, 4.96821, 4.968366, 4.96932, 4.971087, 4.973859, 4.977577, 
    4.982324, 4.9871, 4.991838, 4.99507, 4.998154, 5.000888, 5.00302, 
    5.004251, 5.00424, 5.002608, 4.998962, 4.992938, 4.984252, 4.972774, 
    4.9586, 4.942105, 4.923982, 4.905201, 4.886931, 4.870391, 4.856705, 
    4.846749,
  // height(22,18, 0-49)
    4.926219, 4.930993, 4.935577, 4.939902, 4.943923, 4.94762, 4.950982, 
    4.954012, 4.956714, 4.95909, 4.961139, 4.96284, 4.964164, 4.96506, 
    4.965462, 4.967654, 4.961352, 4.962304, 4.963949, 4.965824, 4.967738, 
    4.967719, 4.967881, 4.967954, 4.96887, 4.970606, 4.973351, 4.977064, 
    4.981887, 4.986845, 4.99204, 4.995138, 4.998181, 5.000986, 5.003305, 
    5.004848, 5.005273, 5.004199, 5.001225, 4.995965, 4.988102, 4.977455, 
    4.964059, 4.948224, 4.930574, 4.912029, 4.893728, 4.876899, 4.862697, 
    4.852058,
  // height(22,19, 0-49)
    4.930254, 4.934838, 4.939164, 4.943184, 4.946876, 4.950236, 4.953277, 
    4.95601, 4.958449, 4.960598, 4.962448, 4.963972, 4.965132, 4.96587, 
    4.966131, 4.967701, 4.959782, 4.961017, 4.963089, 4.965472, 4.967917, 
    4.967721, 4.967884, 4.967977, 4.968936, 4.970692, 4.973415, 4.977076, 
    4.981885, 4.986914, 4.992465, 4.995318, 4.998209, 5.000971, 5.003365, 
    5.005108, 5.005862, 5.005246, 5.002851, 4.998276, 4.991178, 4.981333, 
    4.968722, 4.953592, 4.936501, 4.918311, 4.900126, 4.883163, 4.868595, 
    4.857404,
  // height(22,20, 0-49)
    4.935121, 4.940522, 4.945562, 4.95019, 4.954374, 4.958099, 4.961357, 
    4.964148, 4.966482, 4.968373, 4.969851, 4.970959, 4.971753, 4.972302, 
    4.972693, 0, 4.959976, 4.961293, 4.963098, 4.965001, 4.966878, 4.965349, 
    4.964415, 4.963618, 4.964009, 4.965533, 4.968349, 4.972388, 4.97783, 
    4.983681, 4.990357, 4.993667, 4.997002, 5.000195, 5.003012, 5.00518, 
    5.006382, 5.006256, 5.004407, 5.000442, 4.994011, 4.984875, 4.972975, 
    4.958509, 4.941978, 4.924188, 4.906198, 4.8892, 4.874375, 4.862727,
  // height(22,21, 0-49)
    4.939007, 4.944368, 4.949268, 4.953667, 4.957558, 4.960947, 4.963851, 
    4.966298, 4.968316, 4.969938, 4.971203, 4.972163, 4.972878, 4.973427, 
    4.973916, 0, 4.955731, 4.957488, 4.959795, 4.962227, 4.964609, 4.962763, 
    4.96166, 4.960739, 4.961128, 4.962759, 4.965786, 4.970114, 4.975934, 
    4.982237, 4.989596, 4.992975, 4.996485, 4.999949, 5.003128, 5.00574, 
    5.007459, 5.007914, 5.006705, 5.003426, 4.997713, 4.989299, 4.978093, 
    4.964244, 4.948203, 4.930723, 4.912822, 4.895671, 4.880454, 4.868197,
  // height(22,22, 0-49)
    4.942727, 4.948107, 4.952914, 4.957129, 4.960762, 4.96384, 4.966405, 
    4.968505, 4.970191, 4.971513, 4.972527, 4.973292, 4.973882, 4.974389, 
    4.974936, 0, 4.952352, 4.954473, 4.957218, 4.960129, 4.962974, 4.960836, 
    4.959574, 4.958531, 4.958904, 4.960607, 4.963778, 4.968307, 4.974384, 
    4.980988, 4.988835, 4.992147, 4.995678, 4.999262, 5.002652, 5.005566, 
    5.007674, 5.008605, 5.007951, 5.005296, 5.000262, 4.99256, 4.982064, 
    4.968881, 4.953407, 4.936348, 4.918674, 4.901524, 4.886073, 4.873363,
  // height(22,23, 0-49)
    4.946211, 4.951646, 4.956401, 4.960465, 4.963868, 4.966659, 4.968901, 
    4.970664, 4.972017, 4.973031, 4.973774, 4.974321, 4.974754, 4.975182, 
    4.975747, 0, 4.949856, 4.952229, 4.955276, 4.958517, 4.961682, 4.959258, 
    4.957822, 4.956636, 4.956953, 4.958671, 4.961921, 4.966574, 4.97282, 
    4.979625, 4.98781, 4.991016, 4.994521, 4.998165, 5.001703, 5.004858, 
    5.007296, 5.008648, 5.0085, 5.006428, 5.002038, 4.995022, 4.98522, 
    4.972703, 4.957818, 4.94122, 4.923836, 4.906774, 4.891189, 4.878129,
  // height(22,24, 0-49)
    4.949394, 4.954908, 4.959633, 4.963575, 4.966775, 4.969305, 4.971246, 
    4.972689, 4.973722, 4.97443, 4.9749, 4.975216, 4.975473, 4.975791, 
    4.976331, 0, 4.948518, 4.951012, 4.954212, 4.957628, 4.960968, 4.958356, 
    4.95681, 4.955535, 4.955814, 4.957535, 4.960822, 4.965538, 4.971878, 
    4.978793, 4.987182, 4.990316, 4.993803, 4.997482, 5.001118, 5.004433, 
    5.007102, 5.008749, 5.008963, 5.007317, 5.003409, 4.996915, 4.987658, 
    4.975676, 4.961286, 4.945103, 4.928017, 4.911108, 4.895511, 4.882263,
  // height(22,25, 0-49)
    4.952204, 4.957809, 4.962523, 4.966364, 4.969392, 4.971691, 4.973362, 
    4.97451, 4.975244, 4.975662, 4.975863, 4.975944, 4.97601, 4.976191, 
    4.976657, 0, 4.948055, 4.950538, 4.953739, 4.957167, 4.960527, 4.957858, 
    4.956294, 4.955017, 4.955307, 4.957049, 4.960361, 4.965107, 4.971481, 
    4.978438, 4.986895, 4.990032, 4.993546, 4.99728, 5.001002, 5.004436, 
    5.00726, 5.0091, 5.009548, 5.008173, 5.004572, 4.998418, 4.989519, 
    4.977905, 4.96387, 4.948008, 4.931185, 4.914455, 4.898934, 4.885649,
  // height(22,26, 0-49)
    4.95458, 4.960278, 4.964995, 4.96876, 4.971643, 4.973747, 4.975185, 
    4.976077, 4.97654, 4.97669, 4.976631, 4.976472, 4.976333, 4.976344, 
    4.976682, 0, 4.948453, 4.950796, 4.953845, 4.957116, 4.960338, 4.957754, 
    4.956271, 4.955087, 4.95545, 4.95724, 4.960577, 4.965328, 4.97169, 
    4.978623, 4.98702, 4.990255, 4.993862, 4.997688, 5.001496, 5.005016, 
    5.007926, 5.009855, 5.010394, 5.00912, 5.00563, 4.999599, 4.990843, 
    4.979391, 4.965537, 4.949868, 4.933245, 4.916705, 4.901348, 4.888179,
  // height(22,27, 0-49)
    4.95647, 4.962255, 4.966988, 4.970704, 4.973483, 4.975435, 4.976684, 
    4.977357, 4.977584, 4.977483, 4.977173, 4.976769, 4.976398, 4.976196, 
    4.976342, 0, 4.94983, 4.951895, 4.954633, 4.957582, 4.960505, 4.958111, 
    4.956778, 4.955749, 4.956214, 4.95806, 4.961405, 4.966125, 4.972418, 
    4.979264, 4.98748, 4.990894, 4.994651, 4.998594, 5.002487, 5.006057, 
    5.008984, 5.010896, 5.011392, 5.010053, 5.006485, 5.000376, 4.991556, 
    4.98007, 4.96623, 4.950636, 4.934154, 4.917815, 4.902705, 4.889807,
  // height(22,28, 0-49)
    4.957836, 4.963705, 4.968472, 4.972172, 4.974893, 4.976745, 4.977857, 
    4.978356, 4.978376, 4.978041, 4.977476, 4.976804, 4.976159, 4.975689, 
    4.975567, 0, 4.952566, 4.954219, 4.956491, 4.958948, 4.961411, 4.95925, 
    4.958077, 4.957208, 4.95776, 4.959622, 4.962923, 4.967553, 4.973707, 
    4.980392, 4.988312, 4.991958, 4.995893, 4.999952, 5.003895, 5.00745, 
    5.010296, 5.012068, 5.012367, 5.010787, 5.006949, 5.000559, 4.991478, 
    4.979781, 4.965812, 4.950198, 4.933821, 4.917719, 4.90296, 4.890495,
  // height(22,29, 0-49)
    4.95867, 4.964626, 4.969453, 4.973186, 4.975905, 4.977718, 4.978745, 
    4.979113, 4.978947, 4.978374, 4.97753, 4.976545, 4.975567, 4.974751, 
    4.974271, 0, 4.95646, 4.95757, 4.959221, 4.961021, 4.962852, 4.960859, 
    4.959756, 4.958962, 4.95951, 4.961305, 4.96448, 4.968947, 4.974889, 
    4.981332, 4.988841, 4.992712, 4.996807, 5.000953, 5.004909, 5.008403, 
    5.011117, 5.012687, 5.012722, 5.010827, 5.006638, 4.999887, 4.990465, 
    4.978487, 4.964337, 4.94868, 4.932421, 4.916602, 4.902275, 4.890357,
  // height(22,30, 0-49)
    4.958047, 4.963116, 4.967086, 4.970015, 4.972012, 4.973216, 4.973781, 
    4.973852, 4.973566, 4.973029, 4.972315, 4.97146, 4.970461, 4.969284, 
    4.96787, 4.971422, 4.957416, 4.958146, 4.959991, 4.962359, 4.964968, 
    4.964603, 4.964927, 4.965328, 4.966667, 4.968801, 4.971864, 4.975824, 
    4.980929, 4.98633, 4.992523, 4.995769, 4.999239, 5.002778, 5.006158, 
    5.009108, 5.011305, 5.01238, 5.011932, 5.009561, 5.00491, 4.997726, 
    4.987928, 4.975666, 4.961368, 4.945735, 4.929695, 4.914293, 4.900559, 
    4.889373,
  // height(22,31, 0-49)
    4.95789, 4.963067, 4.967144, 4.970172, 4.972244, 4.973488, 4.974046, 
    4.974065, 4.973676, 4.972998, 4.972118, 4.97109, 4.969933, 4.968622, 
    4.967101, 4.971066, 4.959039, 4.959276, 4.960526, 4.96225, 4.964221, 
    4.963971, 4.964255, 4.964615, 4.965906, 4.968037, 4.971161, 4.975234, 
    4.980437, 4.98588, 4.991862, 4.995546, 4.999402, 5.003253, 5.00686, 
    5.009934, 5.012142, 5.013105, 5.012422, 5.009698, 5.004597, 4.9969, 
    4.986571, 4.973823, 4.959142, 4.94329, 4.927226, 4.912013, 4.898664, 
    4.888015,
  // height(22,32, 0-49)
    4.957166, 4.962335, 4.966437, 4.969514, 4.971652, 4.972965, 4.973582, 
    4.97364, 4.973271, 4.972588, 4.971687, 4.970632, 4.969455, 4.968151, 
    4.96666, 4.970359, 4.96031, 4.960156, 4.960892, 4.962051, 4.963462, 
    4.963401, 4.963728, 4.964138, 4.96545, 4.967617, 4.970803, 4.974948, 
    4.980169, 4.985564, 4.991252, 4.995315, 4.999488, 5.003579, 5.007331, 
    5.010444, 5.012566, 5.013313, 5.012284, 5.009094, 5.003433, 4.995127, 
    4.984194, 4.970913, 4.955841, 4.939794, 4.923772, 4.908843, 4.895998, 
    4.886026,
  // height(22,33, 0-49)
    4.955983, 4.961055, 4.965122, 4.968218, 4.970413, 4.971811, 4.972531, 
    4.972694, 4.972424, 4.971832, 4.971011, 4.970033, 4.968942, 4.967745, 
    4.966402, 4.969375, 4.961257, 4.960827, 4.96114, 4.961818, 4.962752, 
    4.962927, 4.963367, 4.963902, 4.965289, 4.967519, 4.970751, 4.974916, 
    4.980073, 4.985337, 4.990673, 4.995048, 4.999469, 5.003721, 5.007534, 
    5.010592, 5.01253, 5.012957, 5.011473, 5.007711, 5.001394, 4.992397, 
    4.980807, 4.966975, 4.951529, 4.935343, 4.919448, 4.904913, 4.892695, 
    4.883534,
  // height(22,34, 0-49)
    4.954448, 4.95936, 4.963346, 4.966434, 4.968682, 4.970178, 4.971027, 
    4.971339, 4.971222, 4.970782, 4.970108, 4.969277, 4.968343, 4.967324, 
    4.966204, 4.968204, 4.961935, 4.961338, 4.961315, 4.96159, 4.962114, 
    4.962554, 4.963157, 4.963874, 4.965377, 4.967681, 4.970933, 4.975061, 
    4.980067, 4.985126, 4.99007, 4.994689, 4.999281, 5.003613, 5.007399, 
    5.010306, 5.01196, 5.011963, 5.009924, 5.005498, 4.998452, 4.988713, 
    4.976445, 4.962076, 4.946308, 4.930067, 4.914408, 4.900389, 4.888928, 
    4.880701,
  // height(22,35, 0-49)
    4.952672, 4.957375, 4.961246, 4.964301, 4.966592, 4.968191, 4.969186, 
    4.969673, 4.969746, 4.969497, 4.969015, 4.968374, 4.967635, 4.966836, 
    4.965979, 4.966949, 4.962429, 4.961751, 4.961463, 4.961401, 4.961579, 
    4.962293, 4.96309, 4.964033, 4.965674, 4.968048, 4.971286, 4.975313, 
    4.980082, 4.984866, 4.989388, 4.994173, 4.99885, 5.00317, 5.006832, 
    5.00949, 5.010759, 5.010242, 5.00756, 5.002398, 4.994569, 4.984073, 
    4.971148, 4.9563, 4.940302, 4.924123, 4.908833, 4.895466, 4.88489, 
    4.877709,
  // height(22,36, 0-49)
    4.950771, 4.955221, 4.958945, 4.961947, 4.96427, 4.965969, 4.967115, 
    4.96779, 4.968071, 4.968041, 4.967778, 4.967352, 4.96683, 4.966259, 
    4.965673, 4.965696, 4.962821, 4.962123, 4.961627, 4.961285, 4.961173, 
    4.96215, 4.963158, 4.96435, 4.96614, 4.968571, 4.97175, 4.975606, 
    4.980051, 4.984489, 4.988561, 4.993416, 4.99808, 5.002285, 5.005719, 
    5.008024, 5.008811, 5.007683, 5.004285, 4.998341, 4.98972, 4.978488, 
    4.96497, 4.949749, 4.933655, 4.917694, 4.902929, 4.890361, 4.880794, 
    4.874759,
  // height(22,37, 0-49)
    4.948856, 4.953017, 4.956562, 4.959488, 4.961827, 4.963615, 4.964911, 
    4.965777, 4.966276, 4.966475, 4.966443, 4.966245, 4.965945, 4.9656, 
    4.965266, 4.964514, 4.963181, 4.962499, 4.961835, 4.961262, 4.960908, 
    4.962128, 4.963348, 4.964801, 4.966734, 4.969196, 4.972267, 4.975879, 
    4.979912, 4.983932, 4.987516, 4.992332, 4.996866, 5.000842, 5.003934, 
    5.005777, 5.005983, 5.004169, 5.000006, 4.993264, 4.983874, 4.971982, 
    4.957987, 4.942545, 4.926535, 4.910977, 4.896918, 4.885301, 4.876864, 
    4.872054,
  // height(22,38, 0-49)
    4.947029, 4.95087, 4.954208, 4.957035, 4.959365, 4.961228, 4.962661, 
    4.96371, 4.964424, 4.964855, 4.965057, 4.965089, 4.965008, 4.964876, 
    4.964758, 4.963451, 4.963553, 4.962902, 4.962105, 4.961343, 4.960793, 
    4.962229, 4.963652, 4.965358, 4.967416, 4.969876, 4.972776, 4.976065, 
    4.979594, 4.983118, 4.98617, 4.990817, 4.995093, 4.99871, 5.00134, 
    5.002613, 5.00215, 4.999588, 4.994634, 4.987115, 4.977029, 4.964597, 
    4.950294, 4.934833, 4.919126, 4.904189, 4.891028, 4.880522, 4.873323, 
    4.869796,
  // height(22,39, 0-49)
    4.945388, 4.948878, 4.95198, 4.954679, 4.956977, 4.958889, 4.960439, 
    4.961655, 4.962572, 4.963227, 4.96366, 4.963917, 4.964046, 4.964107, 
    4.964168, 4.96253, 4.963966, 4.963343, 4.962438, 4.96153, 4.960828, 
    4.962446, 4.964049, 4.965991, 4.968144, 4.970555, 4.973221, 4.976102, 
    4.979031, 4.981975, 4.984433, 4.988768, 4.992643, 4.995764, 4.997804, 
    4.9984, 4.997189, 4.993839, 4.988104, 4.979869, 4.969203, 4.956405, 
    4.94201, 4.926777, 4.911627, 4.89755, 4.885493, 4.876248, 4.870383, 
    4.868177,
  // height(22,40, 0-49)
    4.944005, 4.947119, 4.949958, 4.952499, 4.954735, 4.956668, 4.958309, 
    4.959668, 4.960769, 4.96163, 4.962281, 4.962752, 4.96308, 4.963314, 
    4.963518, 4.961757, 4.964414, 4.963816, 4.962826, 4.961812, 4.960998, 
    4.962762, 4.964519, 4.966666, 4.968871, 4.971179, 4.973535, 4.975921, 
    4.978155, 4.980425, 4.982213, 4.986079, 4.989399, 4.99188, 4.993204, 
    4.993023, 4.991001, 4.986851, 4.980374, 4.971526, 4.960449, 4.947505, 
    4.933281, 4.918559, 4.904246, 4.891278, 4.880527, 4.87269, 4.868237, 
    4.867364,
  // height(22,41, 0-49)
    4.942934, 4.945651, 4.948199, 4.950552, 4.952695, 4.954617, 4.956311, 
    4.957786, 4.959041, 4.960086, 4.960935, 4.961604, 4.962116, 4.962505, 
    4.962822, 4.961109, 4.964873, 4.964289, 4.963243, 4.96216, 4.961271, 
    4.963148, 4.965024, 4.967335, 4.969543, 4.971682, 4.973652, 4.975451, 
    4.976894, 4.978395, 4.979421, 4.98265, 4.985257, 4.986954, 4.987439, 
    4.986394, 4.983522, 4.978585, 4.971448, 4.962138, 4.950858, 4.938031, 
    4.924275, 4.910371, 4.897185, 4.885581, 4.876331, 4.870027, 4.86704, 
    4.867486,
  // height(22,42, 0-49)
    4.942198, 4.944501, 4.946737, 4.948874, 4.950887, 4.952759, 4.954475, 
    4.956024, 4.957401, 4.9586, 4.959621, 4.960468, 4.961146, 4.961676, 
    4.962083, 4.960546, 4.965296, 4.964724, 4.963648, 4.962533, 4.961604, 
    4.963559, 4.96552, 4.967943, 4.970094, 4.971998, 4.973501, 4.974625, 
    4.975183, 4.975811, 4.975973, 4.978401, 4.980134, 4.980906, 4.980445, 
    4.978471, 4.974735, 4.969062, 4.961384, 4.951796, 4.940564, 4.928149, 
    4.91518, 4.90241, 4.890639, 4.880638, 4.873065, 4.868399, 4.866908, 
    4.868633,
  // height(22,43, 0-49)
    4.941798, 4.943673, 4.945574, 4.947466, 4.949317, 4.951102, 4.952796, 
    4.954382, 4.95584, 4.957156, 4.958319, 4.959318, 4.960145, 4.9608, 
    4.961287, 4.960012, 4.965619, 4.965061, 4.963984, 4.962872, 4.961929, 
    4.963934, 4.965942, 4.968421, 4.970454, 4.972047, 4.973005, 4.973367, 
    4.972955, 4.97261, 4.971803, 4.973268, 4.973981, 4.973707, 4.972209, 
    4.969264, 4.964683, 4.958358, 4.950296, 4.940651, 4.929743, 4.918052, 
    4.906193, 4.894865, 4.884781, 4.876598, 4.870849, 4.867894, 4.867904, 
    4.870842,
  // height(22,44, 0-49)
    4.941687, 4.943127, 4.944678, 4.9463, 4.947957, 4.949617, 4.95125, 
    4.952827, 4.954327, 4.955722, 4.956991, 4.958113, 4.959068, 4.959835, 
    4.960393, 4.959428, 4.965758, 4.965227, 4.96418, 4.963101, 4.962169, 
    4.964197, 4.966213, 4.968689, 4.970536, 4.971749, 4.972087, 4.97161, 
    4.970154, 4.968743, 4.966866, 4.967227, 4.966793, 4.965372, 4.962781, 
    4.958857, 4.953483, 4.946626, 4.938364, 4.928908, 4.918612, 4.907955, 
    4.897513, 4.88791, 4.87975, 4.87356, 4.869744, 4.868541, 4.870022, 
    4.874084,
  // height(22,45, 0-49)
    4.941793, 4.942795, 4.943985, 4.945317, 4.946753, 4.948253, 4.949785, 
    4.951314, 4.952811, 4.954244, 4.955584, 4.9568, 4.957859, 4.958724, 
    4.959352, 4.958708, 4.965632, 4.96514, 4.964149, 4.963128, 4.962224, 
    4.964252, 4.966239, 4.96865, 4.97025, 4.971015, 4.97067, 4.969294, 
    4.966736, 4.964185, 4.961152, 4.960292, 4.958618, 4.955986, 4.952279, 
    4.947404, 4.941326, 4.934086, 4.92583, 4.916817, 4.907412, 4.898078, 
    4.889328, 4.881688, 4.875639, 4.87157, 4.869749, 4.870298, 4.873192, 
    4.878266,
  // height(22,46, 0-49)
    4.942007, 4.942574, 4.943394, 4.944422, 4.945613, 4.946927, 4.948323, 
    4.949766, 4.951222, 4.952654, 4.954029, 4.955307, 4.956448, 4.957397, 
    4.958094, 4.957758, 4.965144, 4.964711, 4.963798, 4.962851, 4.961987, 
    4.963995, 4.965917, 4.968205, 4.969499, 4.96976, 4.968681, 4.966363, 
    4.962676, 4.958935, 4.954689, 4.952533, 4.949564, 4.9457, 4.940897, 
    4.935141, 4.928477, 4.921025, 4.91299, 4.904661, 4.896404, 4.888639, 
    4.881803, 4.876304, 4.87249, 4.870608, 4.870795, 4.873055, 4.877275, 
    4.88323,
  // height(22,47, 0-49)
    4.942184, 4.942324, 4.942777, 4.943493, 4.944427, 4.94553, 4.946764, 
    4.948091, 4.949472, 4.950871, 4.952249, 4.95356, 4.954759, 4.955781, 
    4.956546, 4.956481, 4.964205, 4.963849, 4.963029, 4.962167, 4.961345, 
    4.963313, 4.965137, 4.967248, 4.968189, 4.967905, 4.966066, 4.96279, 
    4.957972, 4.953028, 4.947546, 4.944068, 4.939801, 4.934735, 4.928899, 
    4.922368, 4.915265, 4.907782, 4.900171, 4.892743, 4.885846, 4.879838, 
    4.875064, 4.87181, 4.870286, 4.870596, 4.872749, 4.876638, 4.882066, 
    4.888757,
  // height(22,48, 0-49)
    4.942157, 4.941879, 4.941971, 4.942379, 4.943048, 4.943933, 4.94499, 
    4.94618, 4.947465, 4.948805, 4.95016, 4.951481, 4.952719, 4.953801, 
    4.954633, 4.95479, 4.962732, 4.962471, 4.961751, 4.960971, 4.960187, 
    4.962099, 4.963796, 4.965682, 4.966233, 4.965381, 4.962782, 4.958564, 
    4.952653, 4.946531, 4.939835, 4.935065, 4.929556, 4.923367, 4.916611, 
    4.909441, 4.902061, 4.894722, 4.887719, 4.881363, 4.875974, 4.871838, 
    4.869196, 4.86821, 4.868954, 4.871396, 4.875418, 4.880815, 4.887309, 
    4.894578,
  // height(22,49, 0-49)
    4.942302, 4.941273, 4.940712, 4.94055, 4.940726, 4.94118, 4.941866, 
    4.942734, 4.943739, 4.944835, 4.945973, 4.947086, 4.948108, 4.94893, 
    4.949424, 4.949001, 4.964243, 4.962885, 4.960816, 4.958843, 4.957083, 
    4.960893, 4.964464, 4.968607, 4.970275, 4.969415, 4.9654, 4.958524, 
    4.948629, 4.938767, 4.928291, 4.922237, 4.915466, 4.908151, 4.900531, 
    4.892879, 4.885505, 4.878732, 4.872895, 4.868293, 4.865188, 4.863756, 
    4.864096, 4.866197, 4.869948, 4.875145, 4.881518, 4.888731, 4.896425, 
    4.904231,
  // height(23,0, 0-49)
    4.895426, 4.901486, 4.90759, 4.913628, 4.919533, 4.92527, 4.930825, 
    4.936199, 4.941404, 4.946454, 4.951359, 4.956124, 4.960742, 4.965197, 
    4.969453, 4.973246, 4.977482, 4.980842, 4.983828, 4.986425, 4.988595, 
    4.990544, 4.991959, 4.992893, 4.993297, 4.993151, 4.992422, 4.991085, 
    4.989092, 4.986431, 4.982956, 4.978846, 4.973688, 4.967337, 4.959653, 
    4.950525, 4.939891, 4.927777, 4.914315, 4.899775, 4.884562, 4.869212, 
    4.85435, 4.840641, 4.828725, 4.819151, 4.812321, 4.808452, 4.807563, 
    4.809484,
  // height(23,1, 0-49)
    4.896116, 4.90232, 4.908538, 4.914664, 4.920634, 4.92641, 4.931978, 
    4.937342, 4.942514, 4.947505, 4.952327, 4.956984, 4.961471, 4.965774, 
    4.969862, 4.97324, 4.977746, 4.980855, 4.983581, 4.985966, 4.987989, 
    4.990112, 4.991745, 4.993001, 4.993792, 4.994096, 4.993859, 4.993059, 
    4.991638, 4.989619, 4.986797, 4.983615, 4.979371, 4.973888, 4.966999, 
    4.958545, 4.948429, 4.936629, 4.923249, 4.908527, 4.892865, 4.876808, 
    4.861016, 4.846209, 4.8331, 4.822316, 4.814339, 4.809461, 4.807758, 
    4.809104,
  // height(23,2, 0-49)
    4.896848, 4.903163, 4.909467, 4.915654, 4.921661, 4.927448, 4.933006, 
    4.938334, 4.943444, 4.948349, 4.953061, 4.957585, 4.961919, 4.966052, 
    4.96996, 4.972911, 4.977615, 4.980476, 4.982946, 4.985118, 4.986993, 
    4.989272, 4.991097, 4.992633, 4.993772, 4.994483, 4.9947, 4.994403, 
    4.993524, 4.99211, 4.989905, 4.987619, 4.98428, 4.979692, 4.973659, 
    4.965992, 4.956553, 4.945277, 4.932223, 4.917595, 4.901763, 4.885261, 
    4.868759, 4.853016, 4.838797, 4.826807, 4.81761, 4.81158, 4.808866, 
    4.809398,
  // height(23,3, 0-49)
    4.897707, 4.904102, 4.910461, 4.91668, 4.922695, 4.928468, 4.933987, 
    4.939251, 4.944274, 4.949068, 4.953646, 4.958017, 4.962181, 4.966132, 
    4.969855, 4.972373, 4.977182, 4.979805, 4.98203, 4.983992, 4.985715, 
    4.988125, 4.990106, 4.991872, 4.993307, 4.994374, 4.994997, 4.99516, 
    4.994784, 4.993926, 4.992285, 4.990835, 4.988363, 4.984661, 4.979513, 
    4.972706, 4.964067, 4.953493, 4.940991, 4.926718, 4.910996, 4.894328, 
    4.877372, 4.860893, 4.845701, 4.832562, 4.822122, 4.814842, 4.810956, 
    4.810467,
  // height(23,4, 0-49)
    4.898767, 4.905207, 4.911588, 4.917809, 4.923801, 4.929531, 4.934984, 
    4.940162, 4.945074, 4.949735, 4.954161, 4.958361, 4.962342, 4.966105, 
    4.969644, 4.971735, 4.976532, 4.978934, 4.980926, 4.982686, 4.984258, 
    4.986763, 4.988861, 4.990802, 4.992469, 4.993831, 4.994809, 4.995383, 
    4.99547, 4.995112, 4.993973, 4.993282, 4.991616, 4.988761, 4.984494, 
    4.978585, 4.970834, 4.9611, 4.949344, 4.935659, 4.920317, 4.903763, 
    4.886617, 4.869635, 4.853644, 4.839461, 4.827805, 4.819223, 4.814049, 
    4.812364,
  // height(23,5, 0-49)
    4.900073, 4.906525, 4.912896, 4.919085, 4.925028, 4.930689, 4.93605, 
    4.941118, 4.945899, 4.950413, 4.95467, 4.958691, 4.962481, 4.966052, 
    4.969409, 4.971094, 4.975749, 4.977942, 4.979719, 4.981287, 4.982709, 
    4.985273, 4.987438, 4.989486, 4.991323, 4.992917, 4.994195, 4.995135, 
    4.995642, 4.995732, 4.995035, 4.995014, 4.994076, 4.992012, 4.988597, 
    4.983593, 4.976781, 4.967987, 4.957124, 4.94423, 4.929503, 4.913324, 
    4.896254, 4.879013, 4.862425, 4.847337, 4.834532, 4.824646, 4.818106, 
    4.815096,
  // height(23,6, 0-49)
    4.901654, 4.908082, 4.914409, 4.920537, 4.926403, 4.931969, 4.937221, 
    4.94216, 4.946796, 4.951147, 4.95523, 4.959061, 4.962658, 4.966038, 
    4.969217, 4.970532, 4.974907, 4.976904, 4.978485, 4.979873, 4.981148, 
    4.983724, 4.985905, 4.987993, 4.989932, 4.991693, 4.993219, 4.994479, 
    4.995372, 4.995861, 4.995553, 4.996108, 4.995815, 4.994474, 4.991864, 
    4.987747, 4.98189, 4.974093, 4.964232, 4.952282, 4.938368, 4.922791, 
    4.906042, 4.888782, 4.87181, 4.855984, 4.842136, 4.830983, 4.823049, 
    4.818624,
  // height(23,7, 0-49)
    4.903516, 4.909886, 4.916139, 4.922179, 4.927942, 4.933392, 4.938515, 
    4.943311, 4.947791, 4.951973, 4.955874, 4.959517, 4.96292, 4.966109, 
    4.96911, 4.97011, 4.974067, 4.975875, 4.977278, 4.9785, 4.979634, 
    4.982173, 4.984315, 4.986372, 4.988348, 4.990219, 4.991941, 4.99348, 
    4.994731, 4.995581, 4.995622, 4.996662, 4.996929, 4.996234, 4.994371, 
    4.991102, 4.986189, 4.979417, 4.970619, 4.959719, 4.946767, 4.931982, 
    4.915766, 4.898709, 4.881564, 4.86518, 4.85042, 4.838073, 4.82876, 4.82288,
  // height(23,8, 0-49)
    4.905653, 4.911932, 4.918082, 4.924006, 4.929646, 4.934963, 4.939943, 
    4.944586, 4.948904, 4.952912, 4.956631, 4.960085, 4.963297, 4.966295, 
    4.969112, 4.969871, 4.973276, 4.974898, 4.97614, 4.977212, 4.978214, 
    4.980665, 4.982713, 4.984673, 4.986623, 4.988544, 4.990419, 4.992204, 
    4.99379, 4.994974, 4.995334, 4.996774, 4.997522, 4.997402, 4.996218, 
    4.993746, 4.989747, 4.98399, 4.976279, 4.966488, 4.954601, 4.940746, 
    4.925236, 4.908576, 4.891455, 4.874695, 4.859173, 4.845736, 4.835096, 
    4.827761,
  // height(23,9, 0-49)
    4.908045, 4.914205, 4.920225, 4.926012, 4.931508, 4.936678, 4.941504, 
    4.945988, 4.95014, 4.953975, 4.957514, 4.960781, 4.963801, 4.966605, 
    4.969224, 4.969835, 4.972563, 4.973999, 4.975098, 4.976038, 4.976922, 
    4.979229, 4.981129, 4.982932, 4.984797, 4.986721, 4.988709, 4.99071, 
    4.992615, 4.994116, 4.994787, 4.996551, 4.997704, 4.998085, 4.997517, 
    4.995781, 4.992645, 4.987872, 4.981241, 4.972581, 4.961812, 4.948979, 
    4.934303, 4.918199, 4.901276, 4.884313, 4.868188, 4.853786, 4.841904, 
    4.833155,
  // height(23,10, 0-49)
    4.910669, 4.916684, 4.922551, 4.928182, 4.93352, 4.938529, 4.943195, 
    4.947515, 4.951498, 4.955161, 4.958521, 4.961602, 4.96443, 4.967033, 
    4.969435, 4.969999, 4.971944, 4.973189, 4.97416, 4.974993, 4.975775, 
    4.977887, 4.979592, 4.981181, 4.982915, 4.984797, 4.986864, 4.989058, 
    4.991269, 4.993081, 4.994066, 4.996086, 4.997576, 4.998394, 4.998374, 
    4.997312, 4.994981, 4.991141, 4.985553, 4.978009, 4.968371, 4.956611, 
    4.942855, 4.927424, 4.910847, 4.893844, 4.877275, 4.862051, 4.849038, 
    4.838949,
  // height(23,11, 0-49)
    4.9135, 4.919349, 4.925044, 4.930502, 4.935669, 4.94051, 4.945008, 
    4.94916, 4.952974, 4.956462, 4.959645, 4.96254, 4.965172, 4.967559, 
    4.969719, 4.970341, 4.971409, 4.972464, 4.973328, 4.974075, 4.974782, 
    4.976649, 4.978117, 4.979452, 4.981015, 4.982821, 4.984939, 4.9873, 
    4.989808, 4.991928, 4.993247, 4.995461, 4.997231, 4.998425, 4.998889, 
    4.998437, 4.996847, 4.993878, 4.989277, 4.98281, 4.974285, 4.963607, 
    4.950817, 4.936144, 4.92003, 4.903127, 4.886267, 4.870369, 4.856357, 
    4.845033,
  // height(23,12, 0-49)
    4.916521, 4.922186, 4.927694, 4.932967, 4.937951, 4.942612, 4.946934, 
    4.950913, 4.954554, 4.957866, 4.960867, 4.963572, 4.965996, 4.968154, 
    4.970044, 4.970819, 4.970935, 4.971805, 4.972583, 4.973278, 4.97394, 
    4.975521, 4.976722, 4.97777, 4.979136, 4.98084, 4.982984, 4.985491, 
    4.988282, 4.990713, 4.99239, 4.994746, 4.996741, 4.998255, 4.999147, 
    4.999241, 4.998323, 4.996156, 4.992476, 4.987025, 4.97957, 4.969954, 
    4.958146, 4.944283, 4.928721, 4.912042, 4.895033, 4.878615, 4.863748, 
    4.851315,
  // height(23,13, 0-49)
    4.919718, 4.925189, 4.930497, 4.935571, 4.940359, 4.944829, 4.948966, 
    4.952762, 4.956221, 4.95935, 4.962162, 4.964666, 4.966873, 4.968783, 
    4.970378, 4.971375, 4.97047, 4.971176, 4.971901, 4.972583, 4.97324, 
    4.9745, 4.975414, 4.976161, 4.977314, 4.978903, 4.981051, 4.983681, 
    4.98674, 4.989478, 4.991546, 4.993996, 4.996167, 4.997951, 4.999214, 
    4.999793, 4.999481, 4.998042, 4.995209, 4.990702, 4.984257, 4.975666, 
    4.964827, 4.951798, 4.936854, 4.920501, 4.903476, 4.886686, 4.871117, 
    4.857717,
  // height(23,14, 0-49)
    4.92309, 4.928356, 4.933453, 4.938313, 4.942891, 4.947155, 4.95109, 
    4.954689, 4.957953, 4.960886, 4.963496, 4.96579, 4.967766, 4.969412, 
    4.970696, 4.97194, 4.96995, 4.970529, 4.971247, 4.971963, 4.972665, 
    4.973577, 4.974202, 4.97465, 4.975592, 4.977057, 4.979191, 4.981923, 
    4.985222, 4.988264, 4.990751, 4.99325, 4.995551, 4.997555, 4.999138, 
    5.000143, 5.000372, 4.999589, 4.997525, 4.993887, 4.988383, 4.980763, 
    4.970865, 4.958676, 4.944394, 4.928452, 4.91153, 4.894514, 4.878398, 
    4.864184,
  // height(23,15, 0-49)
    4.926639, 4.931692, 4.936564, 4.941194, 4.945542, 4.949579, 4.95329, 
    4.956672, 4.959722, 4.962442, 4.964838, 4.966904, 4.968638, 4.970015, 
    4.970989, 4.972441, 4.969296, 4.969801, 4.970569, 4.97138, 4.972188, 
    4.972746, 4.973093, 4.973263, 4.974007, 4.975351, 4.977458, 4.980263, 
    4.983772, 4.9871, 4.99003, 4.992534, 4.99492, 4.997099, 4.99895, 
    5.000324, 5.001028, 5.000831, 4.999461, 4.996616, 4.99198, 4.985271, 
    4.976275, 4.96492, 4.95133, 4.93587, 4.919161, 4.902054, 4.885547, 
    4.870674,
  // height(23,16, 0-49)
    4.93037, 4.935199, 4.939828, 4.944206, 4.948298, 4.952079, 4.95554, 
    4.958678, 4.961491, 4.96398, 4.966144, 4.967977, 4.969463, 4.970573, 
    4.971258, 4.972813, 4.968417, 4.968924, 4.969812, 4.970793, 4.971777, 
    4.971989, 4.972089, 4.97202, 4.972597, 4.973833, 4.975907, 4.978754, 
    4.982432, 4.986019, 4.989403, 4.991866, 4.994292, 4.996596, 4.998665, 
    5.000351, 5.00147, 5.001792, 5.001044, 4.998916, 4.995078, 4.989218, 
    4.981081, 4.970545, 4.957668, 4.942747, 4.926349, 4.909281, 4.892532, 
    4.877156,
  // height(23,17, 0-49)
    4.934283, 4.938868, 4.943231, 4.947325, 4.951125, 4.954617, 4.957797, 
    4.960662, 4.963215, 4.965456, 4.967381, 4.968978, 4.970225, 4.971089, 
    4.971526, 4.973015, 4.967241, 4.967832, 4.968923, 4.970154, 4.971397, 
    4.971285, 4.971189, 4.970938, 4.971395, 4.972552, 4.974586, 4.97745, 
    4.981249, 4.985054, 4.988883, 4.991256, 4.99367, 4.99605, 4.998283, 
    5.000228, 5.001703, 5.002481, 5.002286, 5.000806, 4.997698, 4.992626, 
    4.985308, 4.975571, 4.96342, 4.94909, 4.933088, 4.91618, 4.89933, 4.883603,
  // height(23,18, 0-49)
    4.938361, 4.942673, 4.946726, 4.950492, 4.953959, 4.957124, 4.95999, 
    4.962561, 4.964844, 4.966834, 4.968524, 4.969899, 4.970932, 4.971589, 
    4.971833, 4.973045, 4.96572, 4.966478, 4.967849, 4.969416, 4.971005, 
    4.970614, 4.970387, 4.970029, 4.97043, 4.971549, 4.973553, 4.976407, 
    4.980273, 4.98424, 4.988482, 4.990712, 4.993061, 4.995459, 4.9978, 
    4.999946, 5.001716, 5.002888, 5.003185, 5.00229, 4.99985, 4.995514, 
    4.988973, 4.980016, 4.968597, 4.9549, 4.939373, 4.922735, 4.905919, 
    4.889985,
  // height(23,19, 0-49)
    4.942561, 4.94654, 4.950226, 4.953609, 4.956694, 4.959494, 4.962023, 
    4.964293, 4.96631, 4.96807, 4.969558, 4.970748, 4.971611, 4.972114, 
    4.972234, 4.972956, 4.963853, 4.964847, 4.966568, 4.968548, 4.970571, 
    4.969965, 4.969689, 4.969313, 4.969736, 4.970868, 4.972862, 4.97569, 
    4.979569, 4.98363, 4.988221, 4.990247, 4.992464, 4.994816, 4.9972, 
    4.999482, 5.001488, 5.002994, 5.003723, 5.003355, 5.001528, 4.99788, 
    4.992079, 4.983882, 4.973204, 4.960176, 4.945191, 4.928922, 4.912266, 
    4.896266,
  // height(23,20, 0-49)
    4.947812, 4.952392, 4.956592, 4.960402, 4.963821, 4.966853, 4.969504, 
    4.971782, 4.973697, 4.975266, 4.976511, 4.977463, 4.978164, 4.978666, 
    4.97904, 0, 4.962282, 4.963513, 4.965213, 4.966989, 4.9687, 4.967034, 
    4.965853, 4.964697, 4.964581, 4.965442, 4.967443, 4.970533, 4.974926, 
    4.979701, 4.98531, 4.987769, 4.990425, 4.993213, 4.996024, 4.998729, 
    5.001162, 5.003111, 5.004313, 5.004456, 5.003191, 5.000156, 4.995014, 
    4.987504, 4.977509, 4.965121, 4.950686, 4.934827, 4.918398, 4.902422,
  // height(23,21, 0-49)
    4.952321, 4.956649, 4.960524, 4.963956, 4.966967, 4.969578, 4.971817, 
    4.973706, 4.975272, 4.97654, 4.977539, 4.978305, 4.978885, 4.979341, 
    4.979759, 0, 4.957336, 4.958926, 4.96105, 4.963284, 4.965437, 4.96349, 
    4.962173, 4.960936, 4.960859, 4.961868, 4.964108, 4.967514, 4.972302, 
    4.977538, 4.983817, 4.986392, 4.989252, 4.992331, 4.995506, 4.998638, 
    5.001549, 5.004018, 5.005775, 5.006501, 5.005841, 5.003427, 4.99891, 
    4.992016, 4.982603, 4.970729, 4.956704, 4.941106, 4.924758, 4.90866,
  // height(23,22, 0-49)
    4.956862, 4.960968, 4.964542, 4.967612, 4.970216, 4.972399, 4.974205, 
    4.975675, 4.97685, 4.977767, 4.978467, 4.978996, 4.979407, 4.979776, 
    4.98021, 0, 4.953183, 4.955079, 4.957577, 4.960221, 4.962775, 4.960561, 
    4.959106, 4.957771, 4.957701, 4.958802, 4.961205, 4.96483, 4.969896, 
    4.975457, 4.982234, 4.984813, 4.987763, 4.991016, 4.994449, 4.997913, 
    5.001224, 5.004153, 5.00642, 5.0077, 5.007632, 5.005837, 5.001956, 
    4.995699, 4.986902, 4.975594, 4.962046, 4.946799, 4.930641, 4.914544,
  // height(23,23, 0-49)
    4.961319, 4.96523, 4.968522, 4.971242, 4.973449, 4.975204, 4.976571, 
    4.977608, 4.978371, 4.97891, 4.979281, 4.979536, 4.979744, 4.979992, 
    4.980406, 0, 4.949828, 4.951932, 4.954688, 4.957613, 4.960438, 4.957965, 
    4.956351, 4.954892, 4.954782, 4.955913, 4.958411, 4.962177, 4.967437, 
    4.973226, 4.980362, 4.982919, 4.985924, 4.989314, 4.992963, 4.996723, 
    5.000404, 5.00377, 5.006535, 5.008361, 5.008878, 5.007699, 5.004451, 
    4.998827, 4.990645, 4.979904, 4.966846, 4.951975, 4.936047, 4.920007,
  // height(23,24, 0-49)
    4.965569, 4.969304, 4.972334, 4.974724, 4.976551, 4.977893, 4.978831, 
    4.979438, 4.979786, 4.97994, 4.979965, 4.979927, 4.979905, 4.98, 4.98035, 
    0, 4.947584, 4.949786, 4.952665, 4.955732, 4.958699, 4.956051, 4.954333, 
    4.952793, 4.952653, 4.953795, 4.956342, 4.960189, 4.965566, 4.971498, 
    4.97887, 4.981437, 4.984508, 4.988023, 4.991858, 4.995862, 4.999844, 
    5.003561, 5.006723, 5.008988, 5.009978, 5.009296, 5.006564, 5.001464, 
    4.993795, 4.983542, 4.970922, 4.956411, 4.940742, 4.924834,
  // height(23,25, 0-49)
    4.969476, 4.973059, 4.975853, 4.977944, 4.97942, 4.980377, 4.980908, 
    4.981107, 4.981056, 4.98083, 4.980508, 4.980166, 4.979897, 4.979808, 
    4.980052, 0, 4.946215, 4.948393, 4.951257, 4.954316, 4.95728, 4.954575, 
    4.95283, 4.951283, 4.951154, 4.952318, 4.9549, 4.958794, 4.96423, 
    4.970243, 4.97773, 4.980377, 4.983562, 4.987227, 4.991247, 4.995472, 
    4.999707, 5.003707, 5.007178, 5.009773, 5.011113, 5.010795, 5.008437, 
    5.003716, 4.996426, 4.986541, 4.974265, 4.960062, 4.944643, 4.928911,
  // height(23,26, 0-49)
    4.972922, 4.976376, 4.97897, 4.980797, 4.981965, 4.982578, 4.982746, 
    4.982569, 4.982144, 4.981558, 4.980897, 4.980248, 4.979712, 4.979408, 
    4.979493, 0, 4.945743, 4.947777, 4.950482, 4.953379, 4.956195, 4.95355, 
    4.951866, 4.950394, 4.950324, 4.951531, 4.954144, 4.95806, 4.963513, 
    4.969546, 4.977036, 4.979848, 4.983212, 4.987065, 4.991282, 4.995709, 
    5.000151, 5.00436, 5.008039, 5.010841, 5.012385, 5.012269, 5.010112, 
    5.005596, 4.998515, 4.988846, 4.976793, 4.962817, 4.947624, 4.932106,
  // height(23,27, 0-49)
    4.975794, 4.979151, 4.981586, 4.983203, 4.984118, 4.984444, 4.9843, 
    4.983793, 4.983029, 4.982104, 4.981112, 4.980152, 4.979331, 4.978775, 
    4.978641, 0, 4.946302, 4.948066, 4.950467, 4.953045, 4.955564, 4.953069, 
    4.9515, 4.950153, 4.950165, 4.951417, 4.954041, 4.957945, 4.963362, 
    4.969354, 4.976735, 4.979789, 4.983385, 4.987454, 4.991872, 4.996479, 
    5.001076, 5.005418, 5.009205, 5.012092, 5.013698, 5.013628, 5.011506, 
    5.007021, 4.999983, 4.990378, 4.978427, 4.964598, 4.9496, 4.934321,
  // height(23,28, 0-49)
    4.978009, 4.981311, 4.983644, 4.985114, 4.985842, 4.985948, 4.985551, 
    4.984766, 4.983699, 4.982455, 4.981137, 4.979851, 4.978716, 4.977863, 
    4.977447, 0, 4.948286, 4.949656, 4.951609, 4.953715, 4.955791, 4.953478, 
    4.952028, 4.950802, 4.950869, 4.952122, 4.9547, 4.958529, 4.963839, 
    4.969721, 4.97689, 4.98023, 4.984081, 4.988367, 4.992958, 4.997692, 
    5.002371, 5.006748, 5.010526, 5.01336, 5.014878, 5.014691, 5.012437, 
    5.007819, 5.000664, 4.990985, 4.979025, 4.965273, 4.950454, 4.935455,
  // height(23,29, 0-49)
    4.979519, 4.98282, 4.985117, 4.98652, 4.987142, 4.987102, 4.986516, 
    4.985497, 4.984156, 4.982601, 4.980945, 4.979306, 4.977814, 4.976609, 
    4.975844, 0, 4.951502, 4.952365, 4.95373, 4.955213, 4.956685, 4.954491, 
    4.953069, 4.951875, 4.951902, 4.953065, 4.955513, 4.959191, 4.964319, 
    4.970014, 4.976858, 4.980478, 4.984567, 4.989044, 4.993778, 4.998605, 
    5.003326, 5.007692, 5.011411, 5.01414, 5.015511, 5.015141, 5.012679, 
    5.007847, 5.000496, 4.990666, 4.978632, 4.964911, 4.95025, 4.93554,
  // height(23,30, 0-49)
    4.979384, 4.981814, 4.983278, 4.983901, 4.98382, 4.983175, 4.9821, 
    4.980711, 4.979107, 4.977366, 4.975537, 4.973642, 4.971686, 4.969653, 
    4.967526, 4.968501, 4.95388, 4.953983, 4.955086, 4.956669, 4.958492, 
    4.957497, 4.95718, 4.956963, 4.957675, 4.959179, 4.961603, 4.964932, 
    4.969421, 4.974288, 4.980054, 4.983217, 4.986848, 4.990884, 4.995209, 
    4.999662, 5.004045, 5.008105, 5.011535, 5.013987, 5.015082, 5.014435, 
    5.011695, 5.006598, 4.999016, 4.98902, 4.976917, 4.96326, 4.948817, 
    4.934488,
  // height(23,31, 0-49)
    4.979453, 4.981999, 4.983564, 4.984265, 4.984229, 4.983586, 4.982464, 
    4.980983, 4.979244, 4.977332, 4.97531, 4.973215, 4.971061, 4.968839, 
    4.966521, 4.968116, 4.955175, 4.954739, 4.955228, 4.956167, 4.957366, 
    4.956451, 4.956088, 4.955835, 4.956506, 4.958014, 4.960509, 4.963962, 
    4.96857, 4.97352, 4.979156, 4.9828, 4.986884, 4.991324, 4.995992, 
    5.000715, 5.005282, 5.009428, 5.012842, 5.01517, 5.016033, 5.015054, 
    5.011901, 5.006335, 4.99827, 4.987822, 4.975352, 4.961461, 4.94695, 
    4.932743,
  // height(23,32, 0-49)
    4.978727, 4.981336, 4.98298, 4.983766, 4.983811, 4.983236, 4.982162, 
    4.980702, 4.978957, 4.977013, 4.974936, 4.972773, 4.970546, 4.968249, 
    4.965855, 4.967472, 4.956299, 4.9554, 4.955333, 4.955686, 4.956318, 
    4.955542, 4.955204, 4.95499, 4.955684, 4.95724, 4.959817, 4.963375, 
    4.968049, 4.97302, 4.978463, 4.982544, 4.987028, 4.991814, 4.996756, 
    5.001674, 5.006341, 5.010485, 5.013781, 5.015877, 5.016394, 5.014968, 
    5.011288, 5.00515, 4.996514, 4.985552, 4.97268, 4.958555, 4.944016, 
    4.929998,
  // height(23,33, 0-49)
    4.977302, 4.979942, 4.981656, 4.982538, 4.982697, 4.982244, 4.981289, 
    4.979935, 4.97828, 4.976404, 4.974379, 4.972252, 4.970052, 4.967782, 
    4.965415, 4.966619, 4.957237, 4.955972, 4.955427, 4.955264, 4.955398, 
    4.954807, 4.954551, 4.954451, 4.955221, 4.956857, 4.959517, 4.963147, 
    4.967824, 4.972751, 4.977959, 4.982429, 4.987256, 4.992321, 4.997468, 
    5.002501, 5.007183, 5.011227, 5.014306, 5.01606, 5.016119, 5.014136, 
    5.009826, 5.003026, 4.99375, 4.982231, 4.968952, 4.954619, 4.940107, 
    4.926363,
  // height(23,34, 0-49)
    4.975289, 4.977936, 4.979716, 4.98071, 4.981011, 4.98072, 4.979937, 
    4.978752, 4.977258, 4.975528, 4.97363, 4.971616, 4.969521, 4.967354, 
    4.965097, 4.965625, 4.958004, 4.956473, 4.955529, 4.954925, 4.954628, 
    4.954253, 4.954134, 4.954203, 4.955094, 4.956829, 4.959558, 4.963218, 
    4.967833, 4.972657, 4.977599, 4.982405, 4.987512, 4.992789, 4.998067, 
    5.003136, 5.007743, 5.011593, 5.01435, 5.015658, 5.015156, 5.012516, 
    5.007489, 4.99996, 4.990002, 4.977917, 4.964249, 4.94976, 4.935356, 
    4.921988,
  // height(23,35, 0-49)
    4.972805, 4.975446, 4.977287, 4.978399, 4.978864, 4.978765, 4.978192, 
    4.977223, 4.97594, 4.97441, 4.972696, 4.970852, 4.968914, 4.966905, 
    4.964818, 4.964561, 4.958642, 4.956938, 4.955672, 4.954696, 4.954036, 
    4.953892, 4.953948, 4.954236, 4.955279, 4.957119, 4.959894, 4.963537, 
    4.96802, 4.972685, 4.977338, 4.982416, 4.987737, 4.993151, 4.998478, 
    5.003494, 5.007935, 5.011493, 5.013832, 5.014596, 5.013438, 5.010059, 
    5.004251, 4.995952, 4.985302, 4.972674, 4.958676, 4.944117, 4.929926, 
    4.917049,
  // height(23,36, 0-49)
    4.969972, 4.972589, 4.974487, 4.975722, 4.97636, 4.976475, 4.976136, 
    4.975414, 4.974378, 4.973086, 4.971597, 4.969959, 4.968216, 4.966397, 
    4.964516, 4.963494, 4.959198, 4.957397, 4.955878, 4.954597, 4.953636, 
    4.953732, 4.95399, 4.954529, 4.955745, 4.957692, 4.960482, 4.964052, 
    4.968329, 4.972781, 4.977126, 4.9824, 4.987854, 4.993322, 4.99861, 
    5.00348, 5.007657, 5.010827, 5.01265, 5.01278, 5.01089, 5.006711, 
    5.000083, 4.991011, 4.979698, 4.966591, 4.952356, 4.937846, 4.924, 
    4.911744,
  // height(23,37, 0-49)
    4.966919, 4.969494, 4.971436, 4.972788, 4.973604, 4.973938, 4.973849, 
    4.973393, 4.972626, 4.971597, 4.970358, 4.968953, 4.967428, 4.965818, 
    4.964155, 4.96248, 4.959714, 4.957877, 4.956165, 4.954644, 4.953441, 
    4.953775, 4.954249, 4.955064, 4.95646, 4.9585, 4.961268, 4.964707, 
    4.968708, 4.972888, 4.976903, 4.982288, 4.987783, 4.99321, 4.998359, 
    5.002985, 5.006799, 5.009483, 5.010701, 5.010118, 5.007432, 5.002418, 
    4.994967, 4.985151, 4.973249, 4.959768, 4.945435, 4.931123, 4.917774, 
    4.906282,
  // height(23,38, 0-49)
    4.963768, 4.966279, 4.968248, 4.969707, 4.970693, 4.971244, 4.971407, 
    4.971223, 4.970736, 4.969985, 4.969013, 4.967857, 4.966562, 4.96517, 
    4.963725, 4.96156, 4.96023, 4.958398, 4.956545, 4.954842, 4.953458, 
    4.95402, 4.954714, 4.955815, 4.95739, 4.959505, 4.962207, 4.965453, 
    4.969102, 4.972951, 4.976608, 4.982003, 4.987434, 4.992712, 4.997617, 
    5.001892, 5.005239, 5.007343, 5.007872, 5.006511, 5.002993, 4.997136, 
    4.988894, 4.978408, 4.96603, 4.952328, 4.938067, 4.924137, 4.911459, 
    4.90088,
  // height(23,39, 0-49)
    4.960637, 4.963058, 4.965035, 4.96658, 4.967719, 4.968476, 4.968884, 
    4.968968, 4.968763, 4.968296, 4.967598, 4.966702, 4.965645, 4.964471, 
    4.963233, 4.960762, 4.96077, 4.958971, 4.957023, 4.955193, 4.953681, 
    4.954453, 4.955369, 4.956755, 4.958495, 4.960657, 4.963246, 4.966229, 
    4.969455, 4.972909, 4.976169, 4.981458, 4.986709, 4.99172, 4.996265, 
    5.000077, 5.002857, 5.00429, 5.004058, 5.001873, 4.997508, 4.990834, 
    4.981874, 4.970839, 4.958142, 4.944409, 4.930429, 4.917086, 4.905265, 
    4.895751,
  // height(23,40, 0-49)
    4.95763, 4.959937, 4.961891, 4.963499, 4.964767, 4.965711, 4.966346, 
    4.966689, 4.966758, 4.96657, 4.966147, 4.965512, 4.964697, 4.963742, 
    4.962697, 4.960098, 4.961344, 4.959596, 4.957597, 4.95569, 4.954103, 
    4.95507, 4.956193, 4.957851, 4.959733, 4.961905, 4.964325, 4.966981, 
    4.969707, 4.972701, 4.975508, 4.980567, 4.98551, 4.990129, 4.99419, 
    4.997423, 4.999531, 5.000209, 4.99916, 4.996129, 4.990932, 4.983507, 
    4.973942, 4.962516, 4.949704, 4.936168, 4.922704, 4.910172, 4.8994, 
    4.891098,
  // height(23,41, 0-49)
    4.95484, 4.957002, 4.958905, 4.960543, 4.961915, 4.963018, 4.963856, 
    4.964436, 4.964763, 4.964844, 4.96469, 4.964315, 4.963742, 4.963002, 
    4.962139, 4.959574, 4.961953, 4.96027, 4.958256, 4.956322, 4.954705, 
    4.955848, 4.957162, 4.959065, 4.961057, 4.963192, 4.965388, 4.967646, 
    4.9698, 4.972257, 4.974547, 4.979238, 4.983736, 4.987826, 4.991275, 
    4.993814, 4.995153, 4.995003, 4.993098, 4.989223, 4.983247, 4.975173, 
    4.965159, 4.953546, 4.940858, 4.927775, 4.915082, 4.903592, 4.89406, 
    4.887104,
  // height(23,42, 0-49)
    4.952335, 4.954322, 4.956143, 4.957779, 4.959219, 4.960448, 4.961461, 
    4.962251, 4.962814, 4.963148, 4.963252, 4.963131, 4.962798, 4.962269, 
    4.961581, 4.959179, 4.962581, 4.960975, 4.958985, 4.95707, 4.955463, 
    4.956761, 4.958241, 4.960354, 4.962413, 4.964461, 4.966369, 4.96816, 
    4.96967, 4.971512, 4.973205, 4.977383, 4.981291, 4.984713, 4.987421, 
    4.989151, 4.989631, 4.988597, 4.985819, 4.981133, 4.974466, 4.965889, 
    4.955624, 4.944065, 4.931768, 4.919414, 4.907753, 4.897533, 4.889417, 
    4.883925,
  // height(23,43, 0-49)
    4.950162, 4.951948, 4.953654, 4.955253, 4.956722, 4.958042, 4.959195, 
    4.960165, 4.960937, 4.9615, 4.961845, 4.961969, 4.961868, 4.961549, 
    4.961031, 4.958889, 4.963201, 4.961686, 4.959754, 4.957897, 4.956337, 
    4.957767, 4.959386, 4.961664, 4.963741, 4.965644, 4.967198, 4.968454, 
    4.96925, 4.970394, 4.971401, 4.97492, 4.97809, 4.980704, 4.982542, 
    4.983356, 4.982902, 4.980946, 4.977309, 4.971876, 4.964646, 4.955748, 
    4.945463, 4.934228, 4.922611, 4.91127, 4.900899, 4.892162, 4.885618, 
    4.881681,
  // height(23,44, 0-49)
    4.948341, 4.9499, 4.951458, 4.952984, 4.954449, 4.955821, 4.957075, 
    4.958187, 4.959137, 4.959904, 4.96047, 4.960821, 4.960945, 4.960835, 
    4.960487, 4.958665, 4.963771, 4.962362, 4.960526, 4.958759, 4.957273, 
    4.958815, 4.960539, 4.962932, 4.96497, 4.966668, 4.967808, 4.968459, 
    4.968475, 4.968838, 4.96906, 4.971774, 4.974064, 4.975734, 4.976582, 
    4.976389, 4.974941, 4.972054, 4.967598, 4.961523, 4.953889, 4.944887, 
    4.934844, 4.92422, 4.913573, 4.903521, 4.894681, 4.887616, 4.882772, 
    4.88045,
  // height(23,45, 0-49)
    4.946861, 4.948171, 4.949554, 4.950976, 4.952395, 4.95378, 4.955097, 
    4.956316, 4.957407, 4.958346, 4.959108, 4.95967, 4.960007, 4.960099, 
    4.959925, 4.958453, 4.964239, 4.962955, 4.961242, 4.959595, 4.958201, 
    4.959833, 4.961634, 4.964084, 4.966026, 4.967455, 4.968119, 4.968105, 
    4.967281, 4.966781, 4.966122, 4.967893, 4.969166, 4.96977, 4.969526, 
    4.968252, 4.96578, 4.961977, 4.956776, 4.950191, 4.942346, 4.933481, 
    4.923957, 4.914234, 4.904842, 4.896333, 4.889235, 4.883993, 4.880938, 
    4.880261,
  // height(23,46, 0-49)
    4.945683, 4.946728, 4.947913, 4.949197, 4.950539, 4.951898, 4.953238, 
    4.954524, 4.955721, 4.9568, 4.957727, 4.958476, 4.959012, 4.959301, 
    4.959304, 4.958188, 4.964537, 4.963399, 4.961836, 4.96033, 4.959041, 
    4.960747, 4.962584, 4.965035, 4.966822, 4.967922, 4.968055, 4.967322, 
    4.965609, 4.964171, 4.962538, 4.963241, 4.963384, 4.962819, 4.961406, 
    4.959006, 4.955505, 4.950835, 4.944994, 4.938061, 4.930218, 4.921744, 
    4.913013, 4.904469, 4.896591, 4.889844, 4.884655, 4.881347, 4.88013, 
    4.881088,
  // height(23,47, 0-49)
    4.944736, 4.945503, 4.946472, 4.947594, 4.948827, 4.950127, 4.951453, 
    4.952766, 4.954033, 4.955215, 4.956281, 4.957191, 4.957909, 4.958385, 
    4.958569, 4.957788, 4.964588, 4.96362, 4.962227, 4.960876, 4.959701, 
    4.961462, 4.963302, 4.965695, 4.96727, 4.967989, 4.967543, 4.96605, 
    4.96341, 4.960971, 4.958283, 4.957822, 4.956746, 4.954939, 4.952308, 
    4.948769, 4.944271, 4.938815, 4.932464, 4.925364, 4.917743, 4.909908, 
    4.902228, 4.895111, 4.888963, 4.884154, 4.880991, 4.879674, 4.8803, 
    4.882845,
  // height(23,48, 0-49)
    4.943918, 4.9444, 4.945139, 4.946082, 4.947184, 4.948393, 4.949674, 
    4.950984, 4.952284, 4.953536, 4.954707, 4.955752, 4.956629, 4.957283, 
    4.957647, 4.957171, 4.964309, 4.96353, 4.962326, 4.961139, 4.960081, 
    4.961879, 4.963689, 4.965969, 4.967283, 4.967573, 4.966515, 4.964235, 
    4.960649, 4.957168, 4.953364, 4.951672, 4.949322, 4.946239, 4.942382, 
    4.93773, 4.932302, 4.926166, 4.919459, 4.91238, 4.905197, 4.898226, 
    4.891818, 4.886326, 4.882068, 4.87931, 4.878233, 4.878918, 4.881347, 
    4.885399,
  // height(23,49, 0-49)
    4.943139, 4.943075, 4.943346, 4.94389, 4.944658, 4.945593, 4.946653, 
    4.94779, 4.948959, 4.950121, 4.951228, 4.952226, 4.953055, 4.953636, 
    4.953867, 4.95286, 4.96727, 4.965607, 4.963223, 4.960995, 4.959105, 
    4.962934, 4.966742, 4.971398, 4.97398, 4.974425, 4.972114, 4.967323, 
    4.959898, 4.952757, 4.94517, 4.942115, 4.938286, 4.93369, 4.928385, 
    4.922455, 4.916029, 4.909282, 4.902445, 4.895787, 4.889615, 4.884236, 
    4.879951, 4.877014, 4.875607, 4.87583, 4.877696, 4.881118, 4.885932, 
    4.8919,
  // height(24,0, 0-49)
    4.910848, 4.916671, 4.922301, 4.927701, 4.932858, 4.937772, 4.942453, 
    4.946915, 4.951171, 4.955228, 4.959091, 4.962752, 4.9662, 4.969418, 
    4.972382, 4.974842, 4.97764, 4.97967, 4.981387, 4.98284, 4.984052, 
    4.985279, 4.986291, 4.987188, 4.987974, 4.988667, 4.989259, 4.989744, 
    4.990077, 4.99023, 4.990046, 4.989658, 4.988633, 4.986763, 4.983824, 
    4.979576, 4.973786, 4.966261, 4.95687, 4.945582, 4.932493, 4.917852, 
    4.902067, 4.8857, 4.869432, 4.854009, 4.840175, 4.8286, 4.81981, 4.81415,
  // height(24,1, 0-49)
    4.911695, 4.917596, 4.923278, 4.928706, 4.933865, 4.938758, 4.943394, 
    4.94779, 4.951956, 4.955903, 4.959635, 4.963151, 4.96644, 4.969491, 
    4.972285, 4.974345, 4.977362, 4.979176, 4.980673, 4.981947, 4.983039, 
    4.984436, 4.985643, 4.986808, 4.987906, 4.988943, 4.989892, 4.990752, 
    4.991471, 4.992055, 4.9923, 4.992604, 4.992283, 4.991125, 4.988891, 
    4.985327, 4.980186, 4.973246, 4.964348, 4.95343, 4.940554, 4.92594, 
    4.909973, 4.89321, 4.876342, 4.860144, 4.845407, 4.832861, 4.823102, 
    4.816533,
  // height(24,2, 0-49)
    4.912669, 4.91862, 4.924327, 4.929756, 4.934893, 4.93974, 4.944309, 
    4.948617, 4.952674, 4.956494, 4.960084, 4.963445, 4.966572, 4.969456, 
    4.972089, 4.973764, 4.97696, 4.978581, 4.979879, 4.980993, 4.981977, 
    4.983537, 4.984918, 4.986313, 4.987674, 4.988997, 4.990244, 4.99141, 
    4.992443, 4.993364, 4.993931, 4.994814, 4.995092, 4.994552, 4.992957, 
    4.990049, 4.985571, 4.979286, 4.97101, 4.96065, 4.948229, 4.933926, 
    4.918087, 4.901238, 4.884052, 4.867312, 4.851837, 4.8384, 4.827665, 
    4.820106,
  // height(24,3, 0-49)
    4.91381, 4.919782, 4.925487, 4.93089, 4.935981, 4.940762, 4.945244, 
    4.949446, 4.953381, 4.957063, 4.960503, 4.963704, 4.966669, 4.969393, 
    4.971877, 4.973185, 4.976495, 4.977949, 4.979077, 4.98005, 4.980939, 
    4.982646, 4.984173, 4.98575, 4.987319, 4.988866, 4.990348, 4.991757, 
    4.993032, 4.994204, 4.994997, 4.996337, 4.997099, 4.997078, 4.996046, 
    4.993749, 4.98993, 4.984341, 4.976785, 4.967137, 4.955381, 4.941644, 
    4.92622, 4.909581, 4.892362, 4.875326, 4.859296, 4.845084, 4.833405, 
    4.824807,
  // height(24,4, 0-49)
    4.915136, 4.921102, 4.926778, 4.932133, 4.937155, 4.941853, 4.946233, 
    4.950315, 4.954117, 4.957655, 4.960942, 4.963984, 4.966791, 4.969364, 
    4.971712, 4.972683, 4.976027, 4.977337, 4.978322, 4.979175, 4.979979, 
    4.981809, 4.983449, 4.985155, 4.986871, 4.988581, 4.990238, 4.991829, 
    4.993289, 4.994633, 4.995562, 4.997245, 4.998381, 4.99878, 4.998229, 
    4.996487, 4.993301, 4.988431, 4.98166, 4.972841, 4.961918, 4.948961, 
    4.934201, 4.918041, 4.901056, 4.883966, 4.867583, 4.852731, 4.840173, 
    4.830526,
  // height(24,5, 0-49)
    4.916652, 4.922581, 4.928205, 4.933492, 4.938432, 4.943027, 4.947294, 
    4.951252, 4.954916, 4.958307, 4.961441, 4.964331, 4.966985, 4.969419, 
    4.971646, 4.972317, 4.975591, 4.976784, 4.977652, 4.978406, 4.979137, 
    4.981061, 4.982773, 4.984549, 4.986351, 4.988163, 4.989937, 4.99166, 
    4.993255, 4.994709, 4.995702, 4.997621, 4.999029, 4.999756, 4.999607, 
    4.99836, 4.995777, 4.99162, 4.985671, 4.977759, 4.967791, 4.95578, 
    4.941885, 4.926431, 4.909919, 4.893005, 4.876468, 4.861129, 4.847784, 
    4.837109,
  // height(24,6, 0-49)
    4.918346, 4.924214, 4.929765, 4.934965, 4.939806, 4.944293, 4.948441, 
    4.952268, 4.955794, 4.959041, 4.962029, 4.96477, 4.967284, 4.969589, 
    4.971706, 4.972129, 4.975222, 4.976313, 4.97709, 4.977765, 4.978433, 
    4.980412, 4.982152, 4.983939, 4.985767, 4.98762, 4.989464, 4.991274, 
    4.992972, 4.994491, 4.995498, 4.997561, 4.999152, 5.000124, 5.000306, 
    4.999494, 4.997471, 4.994012, 4.988893, 4.98193, 4.972991, 4.96204, 
    4.949162, 4.934595, 4.918754, 4.902222, 4.885718, 4.870051, 4.856028, 
    4.844377,
  // height(24,7, 0-49)
    4.920202, 4.925986, 4.931444, 4.936544, 4.941278, 4.945648, 4.949674, 
    4.953372, 4.956764, 4.959872, 4.962719, 4.965323, 4.967707, 4.969892, 
    4.971903, 4.972137, 4.97493, 4.975934, 4.976643, 4.977257, 4.977875, 
    4.979867, 4.981587, 4.983323, 4.985119, 4.986961, 4.988832, 4.990698, 
    4.992476, 4.994034, 4.995025, 4.997155, 4.998858, 5.000006, 5.000455, 
    5.000026, 4.99852, 4.995724, 4.991423, 4.985418, 4.977546, 4.96772, 
    4.955954, 4.942404, 4.92739, 4.911408, 4.89511, 4.879266, 4.864686, 
    4.852138,
  // height(24,8, 0-49)
    4.922203, 4.927882, 4.933229, 4.938216, 4.942835, 4.947088, 4.95099, 
    4.954564, 4.957827, 4.960806, 4.963521, 4.965996, 4.968257, 4.970326, 
    4.972233, 4.972349, 4.97472, 4.975642, 4.976302, 4.976875, 4.977454, 
    4.979413, 4.981066, 4.982692, 4.984403, 4.986189, 4.988052, 4.989952, 
    4.991802, 4.993388, 4.994358, 4.996493, 4.998249, 4.999518, 5.000184, 
    5.000089, 4.999055, 4.996887, 4.993373, 4.988306, 4.981501, 4.972822, 
    4.962221, 4.949767, 4.935689, 4.92039, 4.904442, 4.888564, 4.873551, 
    4.860202,
  // height(24,9, 0-49)
    4.924329, 4.929885, 4.935111, 4.939977, 4.944474, 4.948607, 4.95239, 
    4.955841, 4.958982, 4.961837, 4.964429, 4.966784, 4.968927, 4.970881, 
    4.972672, 4.972748, 4.974584, 4.975426, 4.976051, 4.9766, 4.977153, 
    4.97903, 4.980568, 4.982034, 4.983612, 4.985303, 4.987132, 4.989051, 
    4.990974, 4.992595, 4.993559, 4.995654, 4.997419, 4.998772, 4.999612, 
    4.999809, 4.999207, 4.997621, 4.994853, 4.990687, 4.98492, 4.977376, 
    4.967946, 4.956625, 4.943548, 4.929025, 4.913544, 4.897759, 4.88244, 
    4.868397,
  // height(24,10, 0-49)
    4.926576, 4.931991, 4.937082, 4.941818, 4.946189, 4.950202, 4.953865, 
    4.957198, 4.960221, 4.962958, 4.965433, 4.967671, 4.969696, 4.971531, 
    4.973192, 4.97331, 4.974496, 4.975257, 4.975863, 4.976406, 4.976948, 
    4.978693, 4.980071, 4.981329, 4.982737, 4.984304, 4.98608, 4.98801, 
    4.990017, 4.99169, 4.992681, 4.994704, 4.996451, 4.997856, 4.998842, 
    4.999298, 4.999086, 4.998041, 4.995966, 4.992651, 4.98787, 4.981419, 
    4.973136, 4.962947, 4.9509, 4.937212, 4.922284, 4.906702, 4.891196, 
    4.876576,
  // height(24,11, 0-49)
    4.928943, 4.934204, 4.939147, 4.943745, 4.947984, 4.95187, 4.955413, 
    4.958628, 4.961534, 4.964156, 4.966515, 4.968637, 4.97054, 4.972244, 
    4.973755, 4.973986, 4.97442, 4.975101, 4.975702, 4.976256, 4.976806, 
    4.978368, 4.97955, 4.980563, 4.981774, 4.983195, 4.984904, 4.986845, 
    4.988947, 4.990697, 4.991765, 4.993696, 4.995408, 4.996849, 4.997957, 
    4.998643, 4.998786, 4.998235, 4.996804, 4.994276, 4.990419, 4.985002, 
    4.977817, 4.968729, 4.957708, 4.944883, 4.930571, 4.91528, 4.899696, 
    4.884621,
  // height(24,12, 0-49)
    4.931442, 4.936534, 4.941318, 4.945765, 4.949864, 4.953617, 4.957031, 
    4.960122, 4.962908, 4.965411, 4.967651, 4.969649, 4.971423, 4.972981, 
    4.974318, 4.974725, 4.974307, 4.974916, 4.975528, 4.976114, 4.976694, 
    4.978027, 4.978982, 4.979725, 4.98072, 4.981984, 4.983621, 4.985569, 
    4.98778, 4.989639, 4.990843, 4.992671, 4.994336, 4.995801, 4.997019, 
    4.997913, 4.998381, 4.998281, 4.997436, 4.995634, 4.992631, 4.988174, 
    4.982021, 4.973984, 4.963962, 4.952005, 4.938346, 4.923423, 4.907864, 
    4.892451,
  // height(24,13, 0-49)
    4.934093, 4.939003, 4.943612, 4.947893, 4.951836, 4.955441, 4.958715, 
    4.961672, 4.964326, 4.966701, 4.968812, 4.970676, 4.972308, 4.973703, 
    4.974848, 4.975464, 4.974095, 4.974648, 4.975296, 4.975943, 4.976576, 
    4.977641, 4.978346, 4.978808, 4.97958, 4.980684, 4.982246, 4.984205, 
    4.986533, 4.988531, 4.989935, 4.991654, 4.993267, 4.994752, 4.996068, 
    4.997155, 4.997918, 4.99823, 4.997921, 4.996779, 4.994556, 4.990984, 
    4.985788, 4.978738, 4.969673, 4.958571, 4.94559, 4.931089, 4.915645, 
    4.900013,
  // height(24,14, 0-49)
    4.936921, 4.94163, 4.946046, 4.950143, 4.953909, 4.957345, 4.96046, 
    4.963262, 4.96577, 4.968, 4.969966, 4.971681, 4.973152, 4.974371, 
    4.975314, 4.976134, 4.973717, 4.97424, 4.974955, 4.975695, 4.976418, 
    4.977182, 4.977629, 4.977811, 4.978366, 4.979317, 4.980805, 4.982772, 
    4.985224, 4.987384, 4.989049, 4.990658, 4.992219, 4.993719, 4.995128, 
    4.996392, 4.997429, 4.998117, 4.998294, 4.997752, 4.996239, 4.993473, 
    4.989157, 4.983024, 4.974865, 4.964593, 4.952296, 4.938266, 4.923021, 
    4.907284,
  // height(24,15, 0-49)
    4.939954, 4.944445, 4.948641, 4.952525, 4.956085, 4.959326, 4.962252, 
    4.964876, 4.967212, 4.969275, 4.971076, 4.972627, 4.973923, 4.974956, 
    4.975694, 4.976676, 4.973099, 4.973635, 4.974455, 4.975329, 4.976182, 
    4.976626, 4.976819, 4.976738, 4.977095, 4.977906, 4.979325, 4.981301, 
    4.983872, 4.986211, 4.988193, 4.98969, 4.991199, 4.992713, 4.994207, 
    4.995636, 4.996924, 4.997959, 4.998579, 4.99858, 4.99771, 4.995675, 
    4.992167, 4.986881, 4.979572, 4.970099, 4.958487, 4.944963, 4.929991, 
    4.914255,
  // height(24,16, 0-49)
    4.943211, 4.947452, 4.951399, 4.955036, 4.958356, 4.961365, 4.964069, 
    4.966485, 4.968622, 4.970495, 4.972114, 4.973482, 4.974594, 4.975438, 
    4.975983, 4.977036, 4.972176, 4.972776, 4.97375, 4.974805, 4.975837, 
    4.975954, 4.975911, 4.9756, 4.975791, 4.976484, 4.977843, 4.979822, 
    4.982503, 4.985028, 4.98737, 4.988751, 4.990204, 4.991729, 4.993303, 
    4.994886, 4.996407, 4.997757, 4.998783, 4.999278, 4.99899, 4.997621, 
    4.994846, 4.990343, 4.983829, 4.97512, 4.964186, 4.9512, 4.936568, 
    4.920935,
  // height(24,17, 0-49)
    4.946694, 4.950654, 4.95431, 4.957654, 4.960692, 4.963429, 4.965877, 
    4.968051, 4.969965, 4.971627, 4.973047, 4.974223, 4.975149, 4.97581, 
    4.976184, 4.977188, 4.970901, 4.971617, 4.972795, 4.974083, 4.975348, 
    4.975148, 4.974903, 4.974407, 4.974476, 4.975085, 4.976398, 4.978378, 
    4.981153, 4.983857, 4.986584, 4.987842, 4.989233, 4.990761, 4.992407, 
    4.994132, 4.995866, 4.997506, 4.998901, 4.999847, 5.000089, 4.999326, 
    4.997222, 4.993437, 4.987666, 4.979686, 4.969424, 4.956998, 4.942767, 
    4.927331,
  // height(24,18, 0-49)
    4.950392, 4.954015, 4.957329, 4.960334, 4.963038, 4.965462, 4.96762, 
    4.969528, 4.9712, 4.972644, 4.973861, 4.974846, 4.975591, 4.976085, 
    4.976321, 4.97714, 4.969261, 4.970144, 4.971568, 4.973141, 4.974692, 
    4.974195, 4.973797, 4.973176, 4.973178, 4.973746, 4.975035, 4.977013, 
    4.97986, 4.982726, 4.985838, 4.986964, 4.988281, 4.9898, 4.991502, 
    4.99335, 4.99528, 4.997187, 4.998922, 5.000279, 5.001005, 5.000793, 
    4.999304, 4.996184, 4.991109, 4.983826, 4.974225, 4.962378, 4.948599, 
    4.933446,
  // height(24,19, 0-49)
    4.954257, 4.957479, 4.960381, 4.962982, 4.965306, 4.967378, 4.969222, 
    4.970854, 4.972284, 4.973517, 4.974545, 4.975358, 4.975943, 4.976294, 
    4.976423, 4.976936, 4.967296, 4.968376, 4.970076, 4.971971, 4.973859, 
    4.973104, 4.972607, 4.971929, 4.971931, 4.972509, 4.973804, 4.975785, 
    4.978683, 4.981678, 4.985153, 4.986128, 4.987349, 4.988836, 4.990572, 
    4.992523, 4.994625, 4.996772, 4.998816, 5.000549, 5.001719, 5.002016, 
    5.001093, 4.99859, 4.994166, 4.98755, 4.978599, 4.967349, 4.954068, 
    4.939276,
  // height(24,20, 0-49)
    4.959174, 4.962858, 4.966164, 4.969108, 4.971708, 4.973982, 4.975949, 
    4.977625, 4.979029, 4.980179, 4.981099, 4.981818, 4.982371, 4.982801, 
    4.983164, 0, 4.964798, 4.966055, 4.967796, 4.969609, 4.971327, 4.969703, 
    4.968443, 4.967083, 4.966592, 4.9669, 4.968161, 4.970348, 4.973696, 
    4.977341, 4.981765, 4.983172, 4.984841, 4.986776, 4.988951, 4.991327, 
    4.993841, 4.996396, 4.998845, 5.000997, 5.002602, 5.003364, 5.002938, 
    5.000969, 4.997112, 4.991087, 4.982724, 4.972033, 4.959246, 4.944842,
  // height(24,21, 0-49)
    4.963408, 4.966722, 4.969628, 4.972158, 4.974346, 4.976221, 4.977811, 
    4.979146, 4.980244, 4.981132, 4.981833, 4.982378, 4.982804, 4.983163, 
    4.983527, 0, 4.959586, 4.9611, 4.963162, 4.96533, 4.967396, 4.965482, 
    4.964082, 4.96265, 4.96222, 4.962704, 4.964239, 4.966779, 4.970561, 
    4.974705, 4.979818, 4.98141, 4.983339, 4.985602, 4.98816, 4.990963, 
    4.993931, 4.996956, 4.999882, 5.002509, 5.004585, 5.00581, 5.005842, 
    5.004326, 5.000915, 4.995324, 4.987371, 4.97705, 4.964567, 4.950371,
  // height(24,22, 0-49)
    4.967702, 4.970664, 4.973182, 4.975305, 4.977076, 4.978538, 4.979732, 
    4.980693, 4.981451, 4.982034, 4.982473, 4.982803, 4.983067, 4.983329, 
    4.983677, 0, 4.955086, 4.956829, 4.959173, 4.961654, 4.964025, 4.961829, 
    4.960271, 4.958739, 4.958321, 4.95891, 4.960636, 4.963431, 4.967537, 
    4.97206, 4.977712, 4.979404, 4.981507, 4.984018, 4.986888, 4.990057, 
    4.993435, 4.9969, 5.000288, 5.003388, 5.00594, 5.007639, 5.008145, 
    5.007098, 5.004148, 4.999008, 4.99149, 4.981569, 4.969436, 4.955513,
  // height(24,23, 0-49)
    4.971951, 4.974577, 4.976721, 4.978443, 4.979802, 4.980852, 4.98164, 
    4.982214, 4.98261, 4.982863, 4.983012, 4.983098, 4.983173, 4.983312, 
    4.983619, 0, 4.951283, 4.953178, 4.955709, 4.958392, 4.960952, 4.958478, 
    4.956745, 4.95508, 4.954624, 4.955256, 4.957099, 4.960074, 4.964422, 
    4.969233, 4.975299, 4.977072, 4.979327, 4.982063, 4.985225, 4.988744, 
    4.992522, 4.996426, 5.000281, 5.003865, 5.006908, 5.009098, 5.010088, 
    5.009516, 5.007031, 5.002338, 4.995245, 4.985715, 4.973922, 4.960277,
  // height(24,24, 0-49)
    4.976042, 4.978349, 4.980137, 4.981477, 4.982438, 4.983085, 4.983476, 
    4.983662, 4.983689, 4.983603, 4.983446, 4.983268, 4.98313, 4.983118, 
    4.983349, 0, 4.948518, 4.95047, 4.953073, 4.955839, 4.958478, 4.955807, 
    4.953943, 4.952183, 4.951692, 4.952342, 4.954256, 4.957346, 4.961858, 
    4.966876, 4.973243, 4.975129, 4.977551, 4.980509, 4.98394, 4.987772, 
    4.991901, 4.996183, 5.000436, 5.004429, 5.007885, 5.010486, 5.011881, 
    5.011705, 5.009609, 5.005295, 4.998567, 4.989384, 4.97791, 4.964542,
  // height(24,25, 0-49)
    4.979859, 4.981875, 4.983335, 4.984321, 4.984909, 4.985174, 4.985183, 
    4.984993, 4.984659, 4.984231, 4.983762, 4.983307, 4.982939, 4.982748, 
    4.982862, 0, 4.94658, 4.948485, 4.951038, 4.953754, 4.956346, 4.953585, 
    4.951666, 4.949878, 4.949385, 4.95006, 4.952026, 4.955197, 4.959819, 
    4.964978, 4.971531, 4.973589, 4.976222, 4.979423, 4.983128, 4.987259, 
    4.991705, 4.996318, 5.000906, 5.005232, 5.009016, 5.011939, 5.013646, 
    5.013772, 5.011967, 5.007938, 5.00149, 4.992584, 4.981378, 4.968261,
  // height(24,26, 0-49)
    4.983298, 4.98506, 4.986228, 4.986894, 4.987146, 4.987062, 4.986718, 
    4.986174, 4.985493, 4.984731, 4.983946, 4.983204, 4.982584, 4.982186, 
    4.982136, 0, 4.945513, 4.947264, 4.949642, 4.952173, 4.954591, 4.951852, 
    4.949958, 4.948216, 4.947764, 4.948481, 4.95049, 4.953713, 4.958396, 
    4.963634, 4.970265, 4.972566, 4.975461, 4.978936, 4.982924, 4.987339, 
    4.992069, 4.996956, 5.001805, 5.006377, 5.010392, 5.013525, 5.015426, 
    5.015734, 5.014105, 5.01025, 5.003979, 4.99526, 4.984254, 4.97135,
  // height(24,27, 0-49)
    4.986259, 4.987812, 4.988739, 4.989136, 4.989098, 4.988709, 4.988045, 
    4.987175, 4.986165, 4.985077, 4.983976, 4.982936, 4.982043, 4.9814, 
    4.981136, 0, 4.94546, 4.946948, 4.949024, 4.951235, 4.95335, 4.950716, 
    4.948902, 4.947252, 4.946861, 4.947614, 4.949643, 4.952878, 4.957563, 
    4.962814, 4.969408, 4.972008, 4.975201, 4.978966, 4.983234, 4.987912, 
    4.99288, 4.997982, 5.003019, 5.007753, 5.011899, 5.015141, 5.017131, 
    5.017511, 5.015946, 5.012156, 5.005963, 4.997341, 4.986464, 4.973726,
  // height(24,28, 0-49)
    4.988665, 4.990068, 4.990814, 4.991004, 4.990735, 4.990089, 4.989146, 
    4.98798, 4.986658, 4.985248, 4.983824, 4.982468, 4.981272, 4.980346, 
    4.979819, 0, 4.946815, 4.947936, 4.949587, 4.951346, 4.953032, 4.950542, 
    4.948813, 4.947252, 4.946893, 4.947637, 4.949623, 4.952797, 4.957403, 
    4.962586, 4.969032, 4.971952, 4.975448, 4.97949, 4.984002, 4.98889, 
    4.994031, 4.999268, 5.004402, 5.0092, 5.013378, 5.016623, 5.018593, 
    5.018941, 5.017337, 5.013512, 5.007304, 4.998701, 4.987891, 4.975283,
  // height(24,29, 0-49)
    4.990462, 4.991789, 4.992432, 4.992489, 4.992052, 4.991203, 4.990024, 
    4.988585, 4.986959, 4.985222, 4.983455, 4.981752, 4.980217, 4.978965, 
    4.978124, 0, 4.949393, 4.950053, 4.951162, 4.952341, 4.953464, 4.951066, 
    4.949343, 4.947788, 4.947369, 4.948007, 4.949859, 4.952889, 4.957327, 
    4.96235, 4.968523, 4.971735, 4.9755, 4.97978, 4.984496, 4.989554, 
    4.994829, 5.000166, 5.005371, 5.010205, 5.014393, 5.01762, 5.019548, 
    5.019832, 5.018151, 5.014245, 5.007967, 4.999325, 4.988527, 4.976,
  // height(24,30, 0-49)
    4.990738, 4.99121, 4.991029, 4.990311, 4.989165, 4.987687, 4.985961, 
    4.984056, 4.982023, 4.979897, 4.977703, 4.975448, 4.973134, 4.970758, 
    4.968334, 4.967433, 4.952801, 4.952506, 4.95306, 4.954014, 4.955168, 
    4.953628, 4.952737, 4.951961, 4.952108, 4.953052, 4.954916, 4.957685, 
    4.961609, 4.965942, 4.971194, 4.974047, 4.977447, 4.981374, 4.985769, 
    4.990544, 4.995582, 5.000725, 5.005774, 5.010484, 5.014568, 5.017704, 
    5.019542, 5.019734, 5.017958, 5.013961, 5.007609, 4.998928, 4.988154, 
    4.975735,
  // height(24,31, 0-49)
    4.991224, 4.991782, 4.991659, 4.990963, 4.989799, 4.988257, 4.986423, 
    4.984369, 4.982151, 4.979816, 4.977396, 4.974913, 4.972373, 4.969775, 
    4.967119, 4.966956, 4.953699, 4.952859, 4.952815, 4.953157, 4.953729, 
    4.952262, 4.951339, 4.950546, 4.950665, 4.951616, 4.953545, 4.956422, 
    4.960444, 4.964846, 4.969977, 4.973281, 4.977116, 4.981448, 4.986209, 
    4.991305, 4.996608, 5.001957, 5.007145, 5.011923, 5.016, 5.01905, 
    5.020725, 5.020681, 5.018607, 5.014267, 5.007555, 4.998531, 4.987468, 
    4.97485,
  // height(24,32, 0-49)
    4.990952, 4.991582, 4.991526, 4.990881, 4.989748, 4.988213, 4.986357, 
    4.984251, 4.981956, 4.979523, 4.976988, 4.974381, 4.971712, 4.968981, 
    4.966177, 4.966247, 4.954534, 4.953211, 4.952619, 4.952398, 4.952437, 
    4.951101, 4.950212, 4.94947, 4.949618, 4.950622, 4.952628, 4.955601, 
    4.959674, 4.964085, 4.969033, 4.97274, 4.976955, 4.98163, 4.986691, 
    4.992035, 4.99753, 5.003008, 5.008257, 5.013021, 5.017007, 5.019885, 
    5.02131, 5.020944, 5.018488, 5.013731, 5.006595, 4.997181, 4.985804, 
    4.972989,
  // height(24,33, 0-49)
    4.989976, 4.990683, 4.990708, 4.990148, 4.98909, 4.987619, 4.985811, 
    4.983734, 4.981448, 4.979006, 4.976447, 4.973802, 4.971087, 4.968307, 
    4.965442, 4.965351, 4.955271, 4.953551, 4.952481, 4.951764, 4.95134, 
    4.950182, 4.949387, 4.948767, 4.949002, 4.950088, 4.952173, 4.955213, 
    4.959281, 4.96364, 4.968359, 4.972418, 4.976954, 4.981907, 4.987197, 
    4.992716, 4.998327, 5.003853, 5.00908, 5.013745, 5.017552, 5.020169, 
    5.021256, 5.020481, 5.017564, 5.012319, 5.004707, 4.994871, 4.983172, 
    4.970181,
  // height(24,34, 0-49)
    4.988362, 4.989154, 4.989285, 4.98884, 4.9879, 4.986543, 4.984841, 
    4.982858, 4.980649, 4.978268, 4.975753, 4.973141, 4.970451, 4.967691, 
    4.964846, 4.964324, 4.955907, 4.953883, 4.95241, 4.951271, 4.950449, 
    4.949511, 4.948865, 4.948426, 4.948793, 4.949985, 4.952144, 4.955214, 
    4.959218, 4.96347, 4.967926, 4.972286, 4.977082, 4.982247, 4.987697, 
    4.993318, 4.998965, 5.004459, 5.009578, 5.014056, 5.017594, 5.019861, 
    5.020521, 5.019255, 5.015803, 5.010012, 5.001885, 4.991614, 4.979609, 
    4.96648,
  // height(24,35, 0-49)
    4.986187, 4.987076, 4.987331, 4.987029, 4.986242, 4.985043, 4.983495, 
    4.981658, 4.979582, 4.977318, 4.974906, 4.972382, 4.969771, 4.967087, 
    4.964324, 4.963235, 4.956457, 4.954219, 4.952422, 4.950934, 4.949782, 
    4.94909, 4.948639, 4.948434, 4.94897, 4.950284, 4.952501, 4.955562, 
    4.959439, 4.963533, 4.967704, 4.972306, 4.977299, 4.98261, 4.988148, 
    4.993796, 4.9994, 5.004778, 5.009702, 5.013903, 5.017081, 5.018907, 
    5.019053, 5.017218, 5.013171, 5.006792, 4.998133, 4.987436, 4.975163, 
    4.961967,
  // height(24,36, 0-49)
    4.983537, 4.98453, 4.984925, 4.98479, 4.984187, 4.983179, 4.981824, 
    4.980174, 4.978276, 4.976174, 4.973908, 4.971516, 4.969026, 4.966462, 
    4.963827, 4.962144, 4.956951, 4.95458, 4.952532, 4.950767, 4.949354, 
    4.948923, 4.9487, 4.948773, 4.949505, 4.950946, 4.953201, 4.956208, 
    4.959899, 4.963787, 4.967659, 4.972442, 4.977566, 4.982953, 4.988503, 
    4.994096, 4.999576, 5.004749, 5.009388, 5.013221, 5.015947, 5.017244, 
    5.016798, 5.014329, 5.009636, 5.002648, 4.993464, 4.982381, 4.969909, 
    4.956739,
  // height(24,37, 0-49)
    4.980508, 4.981606, 4.982151, 4.982196, 4.981798, 4.981007, 4.979875, 
    4.978444, 4.976758, 4.974855, 4.972772, 4.970547, 4.968214, 4.965799, 
    4.963324, 4.9611, 4.957419, 4.954983, 4.952751, 4.950772, 4.949162, 
    4.949, 4.949028, 4.949411, 4.950358, 4.951927, 4.954195, 4.957103, 
    4.96055, 4.96419, 4.967753, 4.97265, 4.977834, 4.983218, 4.988704, 
    4.99416, 4.999428, 5.004307, 5.008569, 5.01194, 5.014123, 5.014809, 
    5.013699, 5.010541, 5.005176, 4.997579, 4.987903, 4.976503, 4.963933, 
    4.950914,
  // height(24,38, 0-49)
    4.977201, 4.978397, 4.979091, 4.979325, 4.979144, 4.978589, 4.977698, 
    4.976512, 4.975065, 4.97339, 4.971519, 4.969489, 4.967337, 4.965096, 
    4.962796, 4.960145, 4.957889, 4.955441, 4.953079, 4.950952, 4.949204, 
    4.949308, 4.949604, 4.950312, 4.951482, 4.953172, 4.955426, 4.958192, 
    4.96134, 4.964695, 4.967939, 4.972879, 4.978047, 4.983353, 4.988689, 
    4.993921, 4.998884, 5.003378, 5.007168, 5.009984, 5.011538, 5.011535, 
    5.0097, 5.005819, 4.999774, 4.991597, 4.981497, 4.96988, 4.957343, 
    4.944621,
  // height(24,39, 0-49)
    4.973715, 4.974999, 4.975837, 4.976258, 4.976297, 4.975984, 4.975348, 
    4.974423, 4.973234, 4.971807, 4.970172, 4.968362, 4.966412, 4.964359, 
    4.962245, 4.959305, 4.958379, 4.955961, 4.953523, 4.9513, 4.949468, 
    4.949832, 4.950396, 4.951439, 4.95283, 4.954629, 4.956837, 4.959415, 
    4.962219, 4.965253, 4.968168, 4.973073, 4.978147, 4.983289, 4.988388, 
    4.993306, 4.997871, 5.001883, 5.005105, 5.007277, 5.00812, 5.007362, 
    5.004759, 5.000136, 4.993432, 4.984732, 4.974305, 4.962605, 4.950256, 
    4.938003,
  // height(24,40, 0-49)
    4.970154, 4.971507, 4.972474, 4.973073, 4.973326, 4.973255, 4.972881, 
    4.972223, 4.971304, 4.970143, 4.968762, 4.967189, 4.965458, 4.963606, 
    4.96168, 4.958601, 4.958908, 4.956546, 4.954076, 4.951808, 4.949941, 
    4.950551, 4.951377, 4.952746, 4.95435, 4.956237, 4.958365, 4.960715, 
    4.96313, 4.96581, 4.968381, 4.973172, 4.978065, 4.982956, 4.987728, 
    4.992238, 4.996309, 4.999742, 5.002305, 5.003745, 5.003803, 5.002235, 
    4.998837, 4.993484, 4.986167, 4.977036, 4.966411, 4.954787, 4.942811, 
    4.931215,
  // height(24,41, 0-49)
    4.966611, 4.968009, 4.969085, 4.969845, 4.970301, 4.970465, 4.970348, 
    4.969962, 4.969318, 4.968431, 4.967318, 4.965998, 4.964501, 4.962861, 
    4.961126, 4.958048, 4.959484, 4.957199, 4.954734, 4.952466, 4.950603, 
    4.951441, 4.952514, 4.954194, 4.955987, 4.957934, 4.959948, 4.96203, 
    4.964015, 4.966311, 4.968513, 4.973105, 4.977732, 4.982281, 4.98663, 
    4.990634, 4.994115, 4.996872, 4.998685, 4.999315, 4.998528, 4.996117, 
    4.99192, 4.985871, 4.978022, 4.96858, 4.957916, 4.946559, 4.935153, 
    4.924411,
  // height(24,42, 0-49)
    4.963175, 4.964589, 4.965748, 4.966649, 4.96729, 4.967675, 4.967805, 
    4.967684, 4.967317, 4.966709, 4.96587, 4.964814, 4.963562, 4.962146, 
    4.960603, 4.957645, 4.960103, 4.957912, 4.955489, 4.953257, 4.951434, 
    4.952474, 4.953773, 4.955733, 4.957686, 4.959659, 4.961521, 4.963294, 
    4.964817, 4.966691, 4.968498, 4.972802, 4.977069, 4.98118, 4.985012, 
    4.988411, 4.991204, 4.993195, 4.994174, 4.993927, 4.992252, 4.988981, 
    4.984013, 4.977334, 4.969066, 4.959468, 4.948955, 4.938068, 4.927447, 
    4.917754,
  // height(24,43, 0-49)
    4.959915, 4.961318, 4.962533, 4.963548, 4.964352, 4.964938, 4.965301, 
    4.965435, 4.965337, 4.965007, 4.964446, 4.963661, 4.962666, 4.96148, 
    4.960136, 4.957391, 4.960761, 4.95868, 4.956325, 4.954162, 4.952404, 
    4.953622, 4.955115, 4.957315, 4.959389, 4.961347, 4.963018, 4.964441, 
    4.965469, 4.966885, 4.968258, 4.972181, 4.975993, 4.979571, 4.982786, 
    4.985485, 4.987495, 4.988636, 4.988711, 4.987537, 4.984951, 4.980837, 
    4.97515, 4.967946, 4.959401, 4.94983, 4.939674, 4.929479, 4.919853, 
    4.911402,
  // height(24,44, 0-49)
    4.956895, 4.958255, 4.959497, 4.960596, 4.961537, 4.962301, 4.962876, 
    4.963249, 4.963411, 4.963352, 4.963067, 4.962556, 4.961821, 4.960875, 
    4.959737, 4.957268, 4.961443, 4.959482, 4.957224, 4.955157, 4.953481, 
    4.954848, 4.956501, 4.958893, 4.961037, 4.962934, 4.964368, 4.965406, 
    4.965909, 4.966825, 4.967713, 4.971162, 4.974424, 4.97737, 4.979871, 
    4.981776, 4.98292, 4.983132, 4.98225, 4.98012, 4.976628, 4.971716, 
    4.965401, 4.957804, 4.949159, 4.93982, 4.930246, 4.920966, 4.912542, 
    4.905505,
  // height(24,45, 0-49)
    4.954153, 4.955442, 4.956679, 4.957835, 4.958883, 4.959798, 4.960562, 
    4.961154, 4.961558, 4.961758, 4.961742, 4.961503, 4.961034, 4.960333, 
    4.959406, 4.957256, 4.962121, 4.960298, 4.958159, 4.956203, 4.954621, 
    4.95611, 4.957882, 4.960408, 4.962569, 4.964353, 4.96551, 4.966124, 
    4.966069, 4.96644, 4.966787, 4.969665, 4.972278, 4.974496, 4.976191, 
    4.977215, 4.977416, 4.976646, 4.974771, 4.971683, 4.967322, 4.961689, 
    4.95487, 4.947047, 4.938503, 4.929619, 4.920855, 4.912706, 4.905671, 
    4.900196,
  // height(24,46, 0-49)
    4.951709, 4.952902, 4.954107, 4.955286, 4.956411, 4.957448, 4.958375, 
    4.959161, 4.959786, 4.960229, 4.960472, 4.960496, 4.96029, 4.959839, 
    4.959132, 4.957314, 4.962758, 4.961088, 4.95909, 4.957263, 4.955777, 
    4.957358, 4.959206, 4.961804, 4.963924, 4.965539, 4.966373, 4.966525, 
    4.965885, 4.965662, 4.965401, 4.967614, 4.969483, 4.970881, 4.971683, 
    4.97175, 4.970951, 4.969162, 4.966289, 4.962273, 4.957111, 4.950871, 
    4.943702, 4.935844, 4.927619, 4.919419, 4.911686, 4.904869, 4.899387, 
    4.895587,
  // height(24,47, 0-49)
    4.949562, 4.950633, 4.951778, 4.952954, 4.954126, 4.955256, 4.956315, 
    4.957269, 4.95809, 4.958755, 4.959237, 4.959513, 4.959562, 4.959362, 
    4.958882, 4.957393, 4.963307, 4.961806, 4.959966, 4.958274, 4.956888, 
    4.958531, 4.960414, 4.963019, 4.965039, 4.966431, 4.966897, 4.96655, 
    4.965296, 4.964425, 4.963489, 4.964943, 4.965979, 4.966473, 4.966308, 
    4.965361, 4.963523, 4.960705, 4.956856, 4.951973, 4.946115, 4.939414, 
    4.932077, 4.924395, 4.916712, 4.90942, 4.902925, 4.897609, 4.893805, 
    4.891757,
  // height(24,48, 0-49)
    4.94768, 4.948614, 4.949677, 4.950824, 4.952013, 4.953206, 4.954365, 
    4.955455, 4.956445, 4.957305, 4.958005, 4.958517, 4.958811, 4.958855, 
    4.958607, 4.95743, 4.963704, 4.962394, 4.960724, 4.959174, 4.957884, 
    4.959568, 4.961443, 4.963991, 4.965849, 4.966964, 4.967022, 4.966144, 
    4.964246, 4.962679, 4.960994, 4.961605, 4.961727, 4.961245, 4.960056, 
    4.958057, 4.95517, 4.951344, 4.946577, 4.940922, 4.934504, 4.927511, 
    4.920208, 4.912917, 4.905994, 4.899813, 4.894729, 4.891049, 4.889009, 
    4.888746,
  // height(24,49, 0-49)
    4.945692, 4.946275, 4.947063, 4.948007, 4.949056, 4.950163, 4.951286, 
    4.952384, 4.953416, 4.954346, 4.955135, 4.95574, 4.956119, 4.956212, 
    4.955952, 4.954215, 4.967573, 4.965439, 4.962609, 4.960008, 4.957872, 
    4.961558, 4.965416, 4.970356, 4.973582, 4.975026, 4.974078, 4.971011, 
    4.965668, 4.960866, 4.955824, 4.955507, 4.954542, 4.952848, 4.950368, 
    4.947054, 4.942887, 4.937885, 4.932127, 4.925748, 4.918957, 4.912019, 
    4.905252, 4.899001, 4.89361, 4.88939, 4.886611, 4.885452, 4.886003, 
    4.888259,
  // height(25,0, 0-49)
    4.925933, 4.931124, 4.936015, 4.940607, 4.944907, 4.948923, 4.952667, 
    4.956147, 4.959369, 4.962331, 4.965029, 4.967461, 4.969619, 4.971503, 
    4.973116, 4.974247, 4.975694, 4.976534, 4.977195, 4.977763, 4.978303, 
    4.97908, 4.979904, 4.98088, 4.98202, 4.983343, 4.984835, 4.986478, 
    4.988221, 4.990023, 4.991735, 4.993485, 4.994883, 4.995748, 4.995881, 
    4.995065, 4.993076, 4.989686, 4.984684, 4.977894, 4.969201, 4.95857, 
    4.946083, 4.931956, 4.916556, 4.9004, 4.884132, 4.868479, 4.854189, 
    4.841959,
  // height(25,1, 0-49)
    4.927026, 4.932236, 4.937124, 4.941692, 4.945944, 4.949895, 4.953556, 
    4.956938, 4.960046, 4.962883, 4.965448, 4.967741, 4.96976, 4.971508, 
    4.972995, 4.97379, 4.975451, 4.976137, 4.976635, 4.977072, 4.977521, 
    4.978458, 4.979441, 4.980615, 4.981967, 4.983503, 4.985191, 4.98702, 
    4.988934, 4.99092, 4.992792, 4.994941, 4.996752, 4.998055, 4.998661, 
    4.998352, 4.996904, 4.994087, 4.98968, 4.983487, 4.975367, 4.965255, 
    4.953193, 4.939358, 4.924083, 4.907857, 4.891315, 4.875189, 4.860251, 
    4.847242,
  // height(25,2, 0-49)
    4.928236, 4.933441, 4.938304, 4.942826, 4.947015, 4.950887, 4.954455, 
    4.95773, 4.960721, 4.963433, 4.965869, 4.968032, 4.969925, 4.971556, 
    4.972939, 4.973425, 4.975278, 4.975841, 4.976205, 4.97653, 4.976901, 
    4.977989, 4.979106, 4.980435, 4.981947, 4.983635, 4.985459, 4.987404, 
    4.989417, 4.991495, 4.993425, 4.995854, 4.997965, 4.999597, 5.000571, 
    5.000686, 4.999723, 4.997451, 4.993648, 4.988107, 4.980661, 4.97122, 
    4.959781, 4.946479, 4.931597, 4.91558, 4.899025, 4.882655, 4.867242, 
    4.853558,
  // height(25,3, 0-49)
    4.929566, 4.934745, 4.939562, 4.944022, 4.948135, 4.951917, 4.955383, 
    4.958548, 4.961421, 4.964013, 4.966328, 4.968372, 4.970154, 4.971688, 
    4.972991, 4.973203, 4.975204, 4.975671, 4.975931, 4.976166, 4.976469, 
    4.977692, 4.978915, 4.980353, 4.981971, 4.983752, 4.985653, 4.987656, 
    4.989704, 4.991798, 4.993697, 4.996298, 4.998598, 5.000453, 5.001705, 
    5.00216, 5.001616, 4.99985, 4.996643, 4.991779, 4.985082, 4.976425, 
    4.965772, 4.953203, 4.938946, 4.923386, 4.907069, 4.890676, 4.874971, 
    4.860731,
  // height(25,4, 0-49)
    4.931008, 4.93614, 4.940896, 4.945281, 4.949308, 4.952993, 4.956354, 
    4.959407, 4.962167, 4.964643, 4.966847, 4.968788, 4.970478, 4.971931, 
    4.973177, 4.973155, 4.975237, 4.975637, 4.975821, 4.975992, 4.976242, 
    4.977576, 4.978874, 4.98037, 4.982038, 4.983856, 4.98578, 4.987794, 
    4.98983, 4.991879, 4.993676, 4.996348, 4.998741, 5.000727, 5.002164, 
    5.002882, 5.002693, 5.001389, 4.998754, 4.994576, 4.988664, 4.980871, 
    4.971121, 4.959445, 4.946002, 4.931112, 4.915251, 4.899047, 4.883229, 
    4.868569,
  // height(25,5, 0-49)
    4.932553, 4.937619, 4.942299, 4.9466, 4.950532, 4.954118, 4.957373, 
    4.960318, 4.962967, 4.965339, 4.967442, 4.969292, 4.970905, 4.9723, 
    4.973505, 4.973295, 4.975376, 4.975733, 4.975873, 4.975999, 4.976211, 
    4.977631, 4.978968, 4.980473, 4.982137, 4.983939, 4.985843, 4.987827, 
    4.98982, 4.991777, 4.993423, 4.996082, 4.998482, 5.000516, 5.002064, 
    5.002976, 5.003079, 5.002186, 5.000093, 4.996589, 4.991478, 4.984593, 
    4.975825, 4.965151, 4.952667, 4.938615, 4.923396, 4.907567, 4.891808, 
    4.876867,
  // height(25,6, 0-49)
    4.934185, 4.93917, 4.943763, 4.94797, 4.951805, 4.955288, 4.95844, 
    4.961281, 4.963829, 4.966102, 4.968116, 4.96989, 4.97144, 4.97279, 
    4.973968, 4.973625, 4.975606, 4.975941, 4.976063, 4.97617, 4.976358, 
    4.977833, 4.979174, 4.980636, 4.982246, 4.983988, 4.985836, 4.987762, 
    4.989691, 4.991532, 4.992995, 4.995569, 4.997908, 4.999924, 5.001517, 
    5.00256, 5.002903, 5.002374, 5.000784, 4.997931, 4.993614, 4.987652, 
    4.979905, 4.970301, 4.958872, 4.945784, 4.931354, 4.916058, 4.900511, 
    4.885429,
  // height(25,7, 0-49)
    4.935893, 4.940784, 4.94528, 4.949388, 4.953124, 4.956505, 4.959556, 
    4.962297, 4.964751, 4.966934, 4.968871, 4.970577, 4.972075, 4.973391, 
    4.974547, 4.974128, 4.975905, 4.976233, 4.976362, 4.976471, 4.976653, 
    4.97815, 4.979456, 4.980828, 4.98234, 4.983981, 4.985743, 4.987593, 
    4.989452, 4.991168, 4.992439, 4.994873, 4.997096, 4.999042, 5.000629, 
    5.001756, 5.002291, 5.002082, 5.000955, 4.998718, 4.995172, 4.990123, 
    4.983405, 4.974901, 4.964583, 4.952542, 4.939005, 4.924366, 4.909166, 
    4.894073,
  // height(25,8, 0-49)
    4.937671, 4.942457, 4.946848, 4.950853, 4.954486, 4.957766, 4.960718, 
    4.963364, 4.965728, 4.96783, 4.969694, 4.971343, 4.972795, 4.974077, 
    4.975214, 4.97478, 4.976242, 4.976571, 4.97673, 4.976866, 4.977058, 
    4.97854, 4.979775, 4.981012, 4.982388, 4.983896, 4.985551, 4.987316, 
    4.98911, 4.990705, 4.991796, 4.994046, 4.996115, 4.997952, 4.999499, 
    5.00067, 5.001359, 5.001431, 5.000728, 4.999069, 4.996257, 4.992092, 
    4.986383, 4.978979, 4.969792, 4.958836, 4.946263, 4.932373, 4.91763, 
    4.902642,
  // height(25,9, 0-49)
    4.939522, 4.944192, 4.948471, 4.952366, 4.955894, 4.959072, 4.961926, 
    4.964479, 4.966755, 4.96878, 4.970574, 4.972166, 4.973575, 4.974823, 
    4.975928, 4.975544, 4.976576, 4.976916, 4.977123, 4.977306, 4.977529, 
    4.978956, 4.980087, 4.981149, 4.982355, 4.983707, 4.985243, 4.986919, 
    4.988662, 4.990154, 4.991093, 4.993133, 4.995021, 4.996726, 4.998206, 
    4.999397, 5.00021, 5.000529, 5.000213, 4.999092, 4.996973, 4.993648, 
    4.988911, 4.982576, 4.974506, 4.964649, 4.953072, 4.939991, 4.92579, 
    4.911009,
  // height(25,10, 0-49)
    4.941456, 4.945998, 4.950157, 4.953936, 4.957352, 4.960425, 4.963178, 
    4.965636, 4.967824, 4.96977, 4.971497, 4.973028, 4.974387, 4.975594, 
    4.976652, 4.976379, 4.976869, 4.977222, 4.977496, 4.977747, 4.978018, 
    4.979352, 4.980344, 4.981201, 4.982213, 4.983394, 4.984804, 4.986394, 
    4.988105, 4.989521, 4.990354, 4.992166, 4.993861, 4.99542, 4.99682, 
    4.998015, 4.998931, 4.999473, 4.999509, 4.998883, 4.997409, 4.994874, 
    4.991057, 4.985744, 4.978755, 4.969977, 4.959402, 4.947165, 4.933567, 
    4.919079,
  // height(25,11, 0-49)
    4.943488, 4.947892, 4.951918, 4.955572, 4.958869, 4.961828, 4.964473, 
    4.96683, 4.968925, 4.970785, 4.972435, 4.973901, 4.975202, 4.976351, 
    4.977344, 4.977236, 4.977071, 4.977445, 4.9778, 4.978139, 4.978481, 
    4.979679, 4.980506, 4.981133, 4.981936, 4.982936, 4.984219, 4.985733, 
    4.98743, 4.988805, 4.98959, 4.991169, 4.992666, 4.994079, 4.995396, 
    4.996587, 4.997594, 4.998336, 4.998695, 4.998528, 4.99765, 4.995848, 
    4.992891, 4.988542, 4.982579, 4.97484, 4.96525, 4.953867, 4.940912, 
    4.926785,
  // height(25,12, 0-49)
    4.94564, 4.949892, 4.953773, 4.957288, 4.960452, 4.963284, 4.965809, 
    4.968053, 4.970044, 4.971808, 4.973372, 4.974759, 4.975985, 4.977059, 
    4.97797, 4.978063, 4.977129, 4.977533, 4.97799, 4.978438, 4.978873, 
    4.979895, 4.980533, 4.980914, 4.981503, 4.982321, 4.983479, 4.984927, 
    4.986634, 4.988007, 4.988809, 4.990157, 4.991462, 4.992733, 4.993971, 
    4.995159, 4.996251, 4.997179, 4.997838, 4.998092, 4.997764, 4.996637, 
    4.994474, 4.991019, 4.986021, 4.979267, 4.970627, 4.960088, 4.947798, 
    4.934089,
  // height(25,13, 0-49)
    4.947933, 4.952016, 4.955732, 4.959089, 4.962103, 4.964792, 4.967181, 
    4.969296, 4.971166, 4.972819, 4.97428, 4.975571, 4.976707, 4.977689, 
    4.978497, 4.978809, 4.976994, 4.977444, 4.978021, 4.978601, 4.979153, 
    4.979963, 4.980396, 4.980526, 4.980901, 4.981544, 4.982584, 4.983975, 
    4.985711, 4.987123, 4.988012, 4.989138, 4.990263, 4.991405, 4.992577, 
    4.993766, 4.994943, 4.996046, 4.996986, 4.997628, 4.997803, 4.997297, 
    4.995863, 4.99323, 4.989122, 4.983292, 4.975555, 4.965837, 4.95422, 
    4.94097,
  // height(25,14, 0-49)
    4.950387, 4.954278, 4.957808, 4.960986, 4.963825, 4.966348, 4.968579, 
    4.970545, 4.972275, 4.973796, 4.975134, 4.976312, 4.977338, 4.97821, 
    4.978907, 4.979425, 4.97661, 4.97713, 4.977851, 4.978589, 4.979284, 
    4.979852, 4.980071, 4.979954, 4.980126, 4.980606, 4.981539, 4.982883, 
    4.984664, 4.98615, 4.987199, 4.988118, 4.989079, 4.990109, 4.991226, 
    4.99243, 4.993695, 4.994971, 4.996171, 4.997174, 4.99781, 4.99787, 
    4.997099, 4.995217, 4.991927, 4.98695, 4.980062, 4.971135, 4.960188, 
    4.947428,
  // height(25,15, 0-49)
    4.953012, 4.956685, 4.960002, 4.96297, 4.965608, 4.967937, 4.969985, 
    4.971778, 4.973346, 4.974717, 4.975914, 4.976958, 4.977856, 4.978607, 
    4.979187, 4.979874, 4.975935, 4.976555, 4.977448, 4.97837, 4.979236, 
    4.979536, 4.979541, 4.979192, 4.97918, 4.979517, 4.980358, 4.981665, 
    4.983503, 4.985093, 4.986369, 4.987097, 4.987914, 4.988852, 4.989933, 
    4.991162, 4.992521, 4.993965, 4.995416, 4.996754, 4.997815, 4.998388, 
    4.998218, 4.997016, 4.99447, 4.990279, 4.98418, 4.976004, 4.965717, 
    4.95347,
  // height(25,16, 0-49)
    4.955808, 4.959229, 4.9623, 4.965026, 4.967431, 4.969538, 4.971376, 
    4.972972, 4.974357, 4.975558, 4.976596, 4.97749, 4.978249, 4.978869, 
    4.979337, 4.980128, 4.974936, 4.975688, 4.976779, 4.977916, 4.978982, 
    4.978996, 4.978796, 4.978239, 4.978075, 4.978295, 4.979061, 4.980342, 
    4.982244, 4.983959, 4.98552, 4.986079, 4.986772, 4.987638, 4.9887, 
    4.989968, 4.99143, 4.993042, 4.994732, 4.996383, 4.997833, 4.998872, 
    4.999245, 4.998656, 4.996783, 4.993306, 4.987936, 4.98047, 4.970826, 
    4.959108,
  // height(25,17, 0-49)
    4.958763, 4.961892, 4.964672, 4.96712, 4.969258, 4.971113, 4.972718, 
    4.974096, 4.975282, 4.976298, 4.977165, 4.9779, 4.978511, 4.979, 
    4.979367, 4.980179, 4.9736, 4.974513, 4.975829, 4.977204, 4.978499, 
    4.97822, 4.977831, 4.977103, 4.976825, 4.976961, 4.977675, 4.978942, 
    4.980911, 4.982769, 4.984655, 4.985065, 4.985654, 4.986466, 4.987527, 
    4.988847, 4.990417, 4.992199, 4.994118, 4.99606, 4.997868, 4.99933, 
    5.000191, 5.000153, 4.998885, 4.996056, 4.991358, 4.984556, 4.975537, 
    4.964358,
  // height(25,18, 0-49)
    4.961843, 4.964629, 4.967072, 4.969197, 4.971034, 4.972611, 4.973962, 
    4.975113, 4.976092, 4.976921, 4.977616, 4.97819, 4.978654, 4.979015, 
    4.979291, 4.980046, 4.971954, 4.973047, 4.974599, 4.976233, 4.977781, 
    4.977211, 4.976659, 4.975799, 4.975451, 4.975545, 4.976236, 4.977504, 
    4.979541, 4.981548, 4.983785, 4.984062, 4.984563, 4.985336, 4.986408, 
    4.98779, 4.989474, 4.991421, 4.993559, 4.995777, 4.997911, 4.999756, 
    5.001056, 5.001511, 5.000786, 4.998543, 4.99446, 4.988282, 4.979865, 
    4.969234,
  // height(25,19, 0-49)
    4.965, 4.967378, 4.969427, 4.971184, 4.972685, 4.973964, 4.975053, 
    4.975977, 4.976758, 4.977411, 4.977946, 4.978371, 4.978695, 4.978937, 
    4.979131, 4.97977, 4.970062, 4.97134, 4.973125, 4.975019, 4.976834, 
    4.975983, 4.975299, 4.974353, 4.973983, 4.974082, 4.974786, 4.976074, 
    4.978185, 4.980337, 4.982932, 4.983087, 4.983509, 4.98425, 4.985336, 
    4.986781, 4.988577, 4.990685, 4.993031, 4.995503, 4.99794, 5.000132, 
    5.001826, 5.002723, 5.002485, 5.000772, 4.997253, 4.991659, 4.983825, 
    4.973745,
  // height(25,20, 0-49)
    4.96907, 4.971853, 4.97428, 4.976379, 4.978179, 4.979703, 4.980981, 
    4.982036, 4.982894, 4.983582, 4.984131, 4.98457, 4.984934, 4.985262, 
    4.9856, 0, 4.967362, 4.968657, 4.970433, 4.97227, 4.973977, 4.972389, 
    4.971055, 4.969516, 4.968708, 4.968553, 4.969211, 4.970665, 4.973172, 
    4.975917, 4.979388, 4.979959, 4.980811, 4.981984, 4.98349, 4.985337, 
    4.98751, 4.989974, 4.992662, 4.995465, 4.99823, 5.000757, 5.002801, 
    5.00407, 5.004237, 5.002963, 4.999919, 4.994827, 4.987511, 4.977941,
  // height(25,21, 0-49)
    4.972409, 4.974806, 4.976856, 4.978595, 4.980055, 4.981269, 4.982268, 
    4.983077, 4.983721, 4.984225, 4.984614, 4.984921, 4.985179, 4.985434, 
    4.985746, 0, 4.962254, 4.963721, 4.965726, 4.967824, 4.969792, 4.9679, 
    4.966414, 4.964807, 4.964072, 4.964111, 4.965068, 4.966903, 4.969873, 
    4.97314, 4.977301, 4.978094, 4.979231, 4.980741, 4.982622, 4.984862, 
    4.987442, 4.990312, 4.993392, 4.996568, 4.999682, 5.002536, 5.004883, 
    5.006442, 5.00689, 5.005895, 5.003135, 4.998338, 4.991322, 4.982051,
  // height(25,22, 0-49)
    4.97575, 4.977777, 4.979461, 4.980845, 4.981971, 4.982874, 4.983584, 
    4.984133, 4.984543, 4.984839, 4.985049, 4.985203, 4.985339, 4.98551, 
    4.985789, 0, 4.957802, 4.959422, 4.961627, 4.96395, 4.966136, 4.963939, 
    4.962275, 4.960557, 4.959836, 4.959994, 4.961162, 4.963283, 4.966613, 
    4.970295, 4.975018, 4.975973, 4.977332, 4.97912, 4.981323, 4.983923, 
    4.986884, 4.990145, 4.993617, 4.997175, 5.000654, 5.003854, 5.006526, 
    5.008392, 5.009137, 5.008434, 5.005967, 5.001472, 4.994767, 4.985815,
  // height(25,23, 0-49)
    4.97903, 4.9807, 4.98203, 4.983072, 4.98387, 4.984463, 4.984885, 
    4.985168, 4.985334, 4.985412, 4.985426, 4.985411, 4.985411, 4.985483, 
    4.985715, 0, 4.953951, 4.955665, 4.95799, 4.960441, 4.962743, 4.960247, 
    4.958386, 4.956528, 4.955769, 4.955982, 4.957291, 4.959627, 4.96324, 
    4.967253, 4.972426, 4.973531, 4.9751, 4.977151, 4.979666, 4.982618, 
    4.98596, 4.98962, 4.993496, 4.997456, 5.001327, 5.004899, 5.007923, 
    5.010116, 5.011169, 5.010761, 5.00858, 5.00437, 4.997954, 4.989296,
  // height(25,24, 0-49)
    4.982182, 4.983513, 4.984507, 4.985221, 4.985703, 4.985996, 4.986135, 
    4.98615, 4.98607, 4.985919, 4.985728, 4.985533, 4.98538, 4.985335, 
    4.985494, 0, 4.951048, 4.95278, 4.955128, 4.957605, 4.959929, 4.957211, 
    4.9552, 4.953234, 4.952438, 4.952682, 4.954084, 4.956569, 4.960389, 
    4.964658, 4.970174, 4.971457, 4.973247, 4.975561, 4.978374, 4.98165, 
    4.985334, 4.989345, 4.993575, 4.997882, 5.002086, 5.005975, 5.009296, 
    5.011769, 5.013084, 5.012925, 5.010993, 5.007029, 5.000869, 4.992476,
  // height(25,25, 0-49)
    4.985147, 4.986164, 4.986844, 4.98725, 4.987433, 4.987438, 4.9873, 
    4.987053, 4.986725, 4.986343, 4.985937, 4.985548, 4.985225, 4.98504, 
    4.985095, 0, 4.948891, 4.950555, 4.952825, 4.955217, 4.957455, 4.95462, 
    4.952531, 4.950522, 4.949719, 4.949996, 4.95147, 4.954067, 4.958037, 
    4.962492, 4.968243, 4.969755, 4.971803, 4.974401, 4.977515, 4.981103, 
    4.985105, 4.989431, 4.993968, 4.998568, 5.003051, 5.007197, 5.010757, 
    5.013449, 5.014969, 5.015006, 5.013266, 5.009499, 5.003544, 4.99537,
  // height(25,26, 0-49)
    4.987865, 4.9886, 4.988998, 4.98912, 4.989028, 4.98876, 4.988358, 
    4.987854, 4.987276, 4.986655, 4.986023, 4.985425, 4.98491, 4.984558, 
    4.98447, 0, 4.947531, 4.949038, 4.951124, 4.95332, 4.955368, 4.952527, 
    4.950438, 4.948456, 4.947687, 4.948007, 4.94954, 4.952215, 4.956279, 
    4.960855, 4.966729, 4.968522, 4.970867, 4.97377, 4.97719, 4.98108, 
    4.985371, 4.989972, 4.994764, 4.999599, 5.004291, 5.008625, 5.01235, 
    5.015193, 5.01685, 5.017016, 5.015405, 5.011773, 5.005966, 4.997958,
  // height(25,27, 0-49)
    4.990288, 4.990781, 4.990932, 4.990807, 4.990461, 4.989943, 4.989286, 
    4.988528, 4.987698, 4.986828, 4.985954, 4.985124, 4.984395, 4.983844, 
    4.983571, 0, 4.947104, 4.948366, 4.950164, 4.952053, 4.953806, 4.951047, 
    4.949018, 4.947112, 4.946393, 4.946748, 4.948308, 4.951011, 4.9551, 
    4.959718, 4.965595, 4.967705, 4.970366, 4.973579, 4.977294, 4.981462, 
    4.986007, 4.990837, 4.995832, 5.000842, 5.005686, 5.010149, 5.013985, 
    5.016919, 5.018657, 5.018899, 5.017364, 5.013811, 5.008099, 5.000204,
  // height(25,28, 0-49)
    4.992364, 4.99267, 4.992622, 4.992288, 4.991722, 4.990971, 4.990073, 
    4.989061, 4.987968, 4.986831, 4.985691, 4.984602, 4.983626, 4.982843, 
    4.982348, 0, 4.947995, 4.94893, 4.950346, 4.951824, 4.953187, 4.950557, 
    4.948601, 4.946773, 4.946075, 4.946415, 4.947931, 4.950579, 4.954597, 
    4.959157, 4.964909, 4.967333, 4.970298, 4.97379, 4.977762, 4.982154, 
    4.986895, 4.991891, 4.997024, 5.002145, 5.00708, 5.011614, 5.015508, 
    5.018489, 5.020265, 5.020542, 5.019038, 5.015524, 5.009858, 5.002028,
  // height(25,29, 0-49)
    4.99406, 4.994244, 4.994057, 4.993563, 4.992815, 4.991854, 4.990718, 
    4.989445, 4.98807, 4.986638, 4.985197, 4.983812, 4.982553, 4.981504, 
    4.980756, 0, 4.950003, 4.95055, 4.951498, 4.952468, 4.953333, 4.950801, 
    4.948859, 4.947036, 4.946271, 4.946498, 4.947872, 4.950364, 4.954204, 
    4.958596, 4.964083, 4.966768, 4.969983, 4.973703, 4.97788, 4.982456, 
    4.98736, 4.992499, 4.997761, 5.002997, 5.008034, 5.012661, 5.016634, 
    5.019682, 5.021515, 5.021831, 5.020354, 5.016856, 5.011202, 5.003389,
  // height(25,30, 0-49)
    4.994519, 4.993861, 4.992861, 4.991597, 4.990131, 4.988516, 4.986785, 
    4.984964, 4.983063, 4.981089, 4.979038, 4.976903, 4.974685, 4.97239, 
    4.970056, 4.968032, 4.954024, 4.95362, 4.953893, 4.954456, 4.955149, 
    4.953227, 4.951905, 4.950692, 4.950378, 4.950848, 4.952226, 4.954489, 
    4.957869, 4.961644, 4.966294, 4.968657, 4.97154, 4.974941, 4.978828, 
    4.983158, 4.987868, 4.99287, 4.998047, 5.00325, 5.008296, 5.012966, 
    5.017006, 5.020132, 5.02204, 5.022424, 5.021001, 5.017544, 5.01192, 
    5.004138,
  // height(25,31, 0-49)
    4.995345, 4.994719, 4.99372, 4.992418, 4.990875, 4.98914, 4.98725, 
    4.985236, 4.983119, 4.98091, 4.978617, 4.976248, 4.9738, 4.97128, 
    4.968707, 4.967444, 4.954495, 4.953582, 4.953315, 4.953332, 4.953514, 
    4.951689, 4.950369, 4.949167, 4.948839, 4.949316, 4.950732, 4.953062, 
    4.956487, 4.960275, 4.964766, 4.967505, 4.970757, 4.974515, 4.978742, 
    4.983388, 4.988389, 4.993653, 4.999059, 5.004455, 5.009655, 5.014433, 
    5.018531, 5.02166, 5.023511, 5.023779, 5.022181, 5.018497, 5.012614, 
    5.004563,
  // height(25,32, 0-49)
    4.995613, 4.995025, 4.99404, 4.992726, 4.991141, 4.989335, 4.987347, 
    4.985208, 4.982944, 4.980573, 4.978112, 4.975571, 4.972955, 4.970267, 
    4.967512, 4.966613, 4.954969, 4.953597, 4.952828, 4.952345, 4.952063, 
    4.950393, 4.949138, 4.948009, 4.947721, 4.948237, 4.949703, 4.952083, 
    4.955504, 4.959243, 4.96351, 4.966569, 4.97013, 4.97418, 4.978678, 
    4.983575, 4.988803, 4.994267, 4.999846, 5.005381, 5.010685, 5.015527, 
    5.019639, 5.022727, 5.024477, 5.024584, 5.022766, 5.018817, 5.01264, 
    5.00429,
  // height(25,33, 0-49)
    4.995334, 4.994799, 4.993851, 4.992554, 4.990967, 4.989133, 4.987097, 
    4.984889, 4.982537, 4.980067, 4.977499, 4.97485, 4.972124, 4.969328, 
    4.966456, 4.965581, 4.955402, 4.953644, 4.952435, 4.951514, 4.95083, 
    4.949367, 4.948236, 4.947248, 4.947051, 4.947638, 4.949155, 4.951556, 
    4.954919, 4.958547, 4.962534, 4.96586, 4.96967, 4.973946, 4.978648, 
    4.983727, 4.989114, 4.994714, 5.000402, 5.006021, 5.011372, 5.016219, 
    5.020291, 5.023284, 5.024884, 5.024779, 5.022697, 5.01844, 5.011938, 
    5.003271,
  // height(25,34, 0-49)
    4.994516, 4.994058, 4.993176, 4.991931, 4.990377, 4.98856, 4.986521, 
    4.984294, 4.981909, 4.979394, 4.976773, 4.974064, 4.971285, 4.968438, 
    4.965515, 4.964412, 4.955777, 4.953714, 4.952136, 4.950844, 4.949824, 
    4.94861, 4.947661, 4.946874, 4.946813, 4.947495, 4.949058, 4.95145, 
    4.954698, 4.95816, 4.961833, 4.965373, 4.969373, 4.97381, 4.978651, 
    4.983845, 4.989325, 4.994994, 5.000727, 5.006361, 5.011694, 5.016483, 
    5.020451, 5.02329, 5.024677, 5.024305, 5.02191, 5.017309, 5.010454, 
    5.001464,
  // height(25,35, 0-49)
    4.993182, 4.992826, 4.992038, 4.990879, 4.989397, 4.987638, 4.985642, 
    4.983441, 4.98107, 4.978556, 4.975928, 4.97321, 4.970424, 4.967576, 
    4.96466, 4.963175, 4.9561, 4.953816, 4.951942, 4.95035, 4.949063, 
    4.948124, 4.947401, 4.946869, 4.946983, 4.94778, 4.949381, 4.95173, 
    4.954807, 4.958058, 4.961395, 4.965098, 4.969231, 4.97377, 4.978685, 
    4.983928, 4.989433, 4.995101, 5.000806, 5.006383, 5.011625, 5.016284, 
    5.020075, 5.022686, 5.023796, 5.023099, 5.02034, 5.015363, 5.008144, 
    4.998838,
  // height(25,36, 0-49)
    4.99136, 4.991127, 4.990465, 4.989424, 4.988052, 4.986389, 4.984475, 
    4.982344, 4.980028, 4.97756, 4.974968, 4.972284, 4.969531, 4.966724, 
    4.963866, 4.961936, 4.956396, 4.953965, 4.951863, 4.950037, 4.948545, 
    4.947903, 4.94744, 4.947205, 4.947526, 4.948452, 4.950078, 4.95235, 
    4.955209, 4.958213, 4.961207, 4.965024, 4.969234, 4.973816, 4.978744, 
    4.983969, 4.989426, 4.995021, 5.000623, 5.006064, 5.011133, 5.01558, 
    5.019113, 5.02142, 5.022179, 5.021094, 5.017928, 5.012548, 5.004965, 
    4.995371,
  // height(25,37, 0-49)
    4.989093, 4.989005, 4.988489, 4.987594, 4.986362, 4.984831, 4.983038, 
    4.981017, 4.9788, 4.976418, 4.973905, 4.97129, 4.968606, 4.965876, 
    4.963112, 4.960749, 4.956685, 4.954175, 4.951907, 4.949906, 4.948266, 
    4.947929, 4.947752, 4.947848, 4.9484, 4.949461, 4.951101, 4.953265, 
    4.955864, 4.958595, 4.961247, 4.96513, 4.969367, 4.973936, 4.978812, 
    4.983953, 4.989293, 4.994737, 5.000153, 5.005373, 5.010181, 5.014324, 
    5.01751, 5.019426, 5.01976, 5.018228, 5.014614, 5.008818, 5.000887, 
    4.991054,
  // height(25,38, 0-49)
    4.986433, 4.986499, 4.986148, 4.985423, 4.98436, 4.982993, 4.981357, 
    4.979482, 4.977402, 4.975144, 4.972745, 4.970237, 4.967655, 4.965031, 
    4.962386, 4.959657, 4.956991, 4.954454, 4.952072, 4.949954, 4.948216, 
    4.948183, 4.948303, 4.948752, 4.949552, 4.950753, 4.952391, 4.954421, 
    4.956728, 4.959168, 4.961491, 4.965396, 4.969607, 4.974107, 4.978873, 
    4.983865, 4.989013, 4.994225, 4.999371, 5.004277, 5.008728, 5.012469, 
    5.015213, 5.016651, 5.016483, 5.014445, 5.010352, 5.00414, 4.995898, 
    4.985897,
  // height(25,39, 0-49)
    4.98344, 4.983667, 4.983495, 4.982955, 4.982084, 4.980909, 4.979459, 
    4.977764, 4.975853, 4.973757, 4.971507, 4.969138, 4.966689, 4.964193, 
    4.961687, 4.95869, 4.957332, 4.954806, 4.952355, 4.950166, 4.948378, 
    4.948637, 4.949059, 4.949871, 4.950925, 4.952264, 4.953889, 4.955763, 
    4.957753, 4.959896, 4.961904, 4.965787, 4.969928, 4.974308, 4.978906, 
    4.983677, 4.988561, 4.99346, 4.998243, 5.002738, 5.006731, 5.009968, 
    5.01217, 5.013039, 5.012294, 5.0097, 5.00511, 4.998499, 4.990002, 4.97993,
  // height(25,40, 0-49)
    4.980185, 4.980569, 4.980579, 4.980239, 4.979576, 4.978613, 4.977376, 
    4.975892, 4.974182, 4.972278, 4.970209, 4.96801, 4.96572, 4.963377, 
    4.961021, 4.957868, 4.957716, 4.955232, 4.952751, 4.950531, 4.948729, 
    4.949263, 4.949982, 4.951154, 4.952459, 4.953933, 4.955529, 4.957229, 
    4.95889, 4.960732, 4.962445, 4.966266, 4.970292, 4.974501, 4.978872, 
    4.983361, 4.987904, 4.992404, 4.996732, 5.000714, 5.004144, 5.006771, 
    5.008329, 5.008542, 5.007154, 5.003967, 4.998874, 4.9919, 4.983227, 
    4.973203,
  // height(25,41, 0-49)
    4.976741, 4.977275, 4.977466, 4.97733, 4.976886, 4.976152, 4.975149, 
    4.973896, 4.972416, 4.970734, 4.968876, 4.966875, 4.964769, 4.962596, 
    4.960401, 4.957204, 4.958153, 4.95573, 4.953249, 4.951032, 4.949247, 
    4.950036, 4.951032, 4.952551, 4.954097, 4.955692, 4.957246, 4.958759, 
    4.960083, 4.96163, 4.963066, 4.966787, 4.970655, 4.974645, 4.978733, 
    4.982875, 4.987002, 4.991017, 4.994792, 4.998161, 5.000918, 5.00283, 
    5.003649, 5.003125, 5.001037, 4.997231, 4.991654, 4.984376, 4.975628, 
    4.965791,
  // height(25,42, 0-49)
    4.973186, 4.973859, 4.974224, 4.97429, 4.974071, 4.973577, 4.972821, 
    4.971821, 4.970592, 4.969154, 4.967532, 4.965755, 4.963854, 4.96187, 
    4.959843, 4.956702, 4.958642, 4.956295, 4.953839, 4.951653, 4.949909, 
    4.950922, 4.952172, 4.954015, 4.955778, 4.957478, 4.958976, 4.96029, 
    4.961278, 4.962534, 4.963706, 4.967291, 4.970962, 4.974685, 4.978436, 
    4.982165, 4.985803, 4.989247, 4.992375, 4.995026, 4.997008, 4.998106, 
    4.998096, 4.996766, 4.993938, 4.989511, 4.983484, 4.975986, 4.967286, 
    4.957791,
  // height(25,43, 0-49)
    4.969604, 4.970394, 4.970921, 4.971184, 4.971187, 4.970936, 4.970438, 
    4.969702, 4.968741, 4.967569, 4.966205, 4.964672, 4.962998, 4.961216, 
    4.959366, 4.956364, 4.959184, 4.95692, 4.954512, 4.952376, 4.950689, 
    4.951897, 4.953369, 4.955495, 4.957449, 4.959227, 4.960651, 4.961758, 
    4.962413, 4.963387, 4.964305, 4.967716, 4.971148, 4.97456, 4.977921, 
    4.981175, 4.984247, 4.987039, 4.989427, 4.991263, 4.992372, 4.992564, 
    4.99165, 4.989461, 4.985876, 4.980847, 4.974436, 4.966821, 4.958312, 
    4.949332,
  // height(25,44, 0-49)
    4.966064, 4.966953, 4.967626, 4.968073, 4.968293, 4.968284, 4.968047, 
    4.967584, 4.966902, 4.966008, 4.964917, 4.963645, 4.962215, 4.960651, 
    4.958984, 4.956183, 4.95977, 4.9576, 4.955254, 4.953185, 4.951562, 
    4.952929, 4.954587, 4.956951, 4.959055, 4.960881, 4.962212, 4.963103, 
    4.963431, 4.964125, 4.96479, 4.967986, 4.971137, 4.974195, 4.977112, 
    4.979828, 4.982265, 4.984324, 4.98589, 4.986822, 4.986973, 4.986184, 
    4.984309, 4.981235, 4.976897, 4.971315, 4.964608, 4.957005, 4.948846, 
    4.940559,
  // height(25,45, 0-49)
    4.962638, 4.963603, 4.964401, 4.965019, 4.965446, 4.965672, 4.965693, 
    4.965505, 4.965105, 4.964497, 4.96369, 4.962691, 4.961516, 4.960183, 
    4.958711, 4.95615, 4.96039, 4.958319, 4.956052, 4.954056, 4.952502, 
    4.953992, 4.955791, 4.95834, 4.960548, 4.962384, 4.963598, 4.964264, 
    4.96427, 4.96468, 4.965085, 4.968025, 4.97085, 4.973502, 4.975922, 
    4.978043, 4.97978, 4.981034, 4.9817, 4.981656, 4.98078, 4.978958, 
    4.976094, 4.972135, 4.967084, 4.961026, 4.954139, 4.946698, 4.939058, 
    4.931637,
  // height(25,46, 0-49)
    4.959384, 4.960401, 4.961304, 4.962074, 4.962692, 4.963142, 4.963412, 
    4.963494, 4.963376, 4.963057, 4.962538, 4.961819, 4.96091, 4.959814, 
    4.958544, 4.956244, 4.961024, 4.959065, 4.956888, 4.954971, 4.95348, 
    4.955057, 4.95695, 4.959622, 4.961882, 4.963686, 4.964756, 4.965185, 
    4.964869, 4.964985, 4.965108, 4.967745, 4.970198, 4.972394, 4.974265, 
    4.975734, 4.97671, 4.977099, 4.976804, 4.975729, 4.973786, 4.970906, 
    4.967056, 4.962245, 4.956552, 4.950125, 4.9432, 4.936079, 4.92913, 
    4.922746,
  // height(25,47, 0-49)
    4.95635, 4.957393, 4.95838, 4.959281, 4.960072, 4.960729, 4.961237, 
    4.961576, 4.961733, 4.961699, 4.961466, 4.961028, 4.960386, 4.959536, 
    4.958477, 4.956443, 4.961648, 4.959813, 4.957735, 4.955901, 4.954465, 
    4.956092, 4.958033, 4.960762, 4.963014, 4.964739, 4.965635, 4.965809, 
    4.965172, 4.964973, 4.964783, 4.967062, 4.969089, 4.970776, 4.972046, 
    4.972809, 4.972975, 4.972452, 4.971157, 4.969021, 4.966, 4.962074, 
    4.957274, 4.951685, 4.945455, 4.938794, 4.931985, 4.925356, 4.919264, 
    4.914069,
  // height(25,48, 0-49)
    4.953563, 4.954612, 4.955658, 4.956668, 4.957611, 4.958456, 4.959181, 
    4.959764, 4.960183, 4.96042, 4.960465, 4.960305, 4.959929, 4.959326, 
    4.958488, 4.956709, 4.96223, 4.960528, 4.958559, 4.956808, 4.955421, 
    4.957064, 4.959004, 4.961722, 4.963907, 4.965501, 4.966192, 4.966093, 
    4.965123, 4.964581, 4.964033, 4.965894, 4.967434, 4.968557, 4.969174, 
    4.969187, 4.968502, 4.967037, 4.964726, 4.961534, 4.957456, 4.952534, 
    4.946867, 4.940608, 4.933976, 4.927238, 4.920715, 4.914744, 4.909664, 
    4.90578,
  // height(25,49, 0-49)
    4.95051, 4.9514, 4.952364, 4.953356, 4.954337, 4.95527, 4.956123, 
    4.956862, 4.957456, 4.957881, 4.95811, 4.958118, 4.957881, 4.957365, 
    4.956535, 4.954092, 4.966395, 4.963832, 4.960638, 4.957756, 4.955451, 
    4.959006, 4.962871, 4.96796, 4.971593, 4.973686, 4.973638, 4.971708, 
    4.96775, 4.964478, 4.961112, 4.962604, 4.963628, 4.964084, 4.963889, 
    4.962953, 4.961198, 4.958563, 4.95502, 4.950583, 4.945317, 4.939349, 
    4.932869, 4.926122, 4.919407, 4.91305, 4.907397, 4.902774, 4.899466, 
    4.897687,
  // height(26,0, 0-49)
    4.94, 4.944391, 4.94844, 4.952157, 4.95555, 4.958627, 4.961393, 4.963849, 
    4.965998, 4.96784, 4.969378, 4.970623, 4.97159, 4.972304, 4.9728, 
    4.972906, 4.973375, 4.973431, 4.973461, 4.973564, 4.973804, 4.974427, 
    4.975248, 4.976345, 4.977716, 4.979355, 4.981232, 4.983315, 4.985551, 
    4.987894, 4.990223, 4.992686, 4.994967, 4.996955, 4.998531, 4.999562, 
    4.999901, 4.999391, 4.997859, 4.995126, 4.991014, 4.985359, 4.978026, 
    4.968945, 4.958121, 4.945682, 4.931883, 4.917126, 4.901945, 4.886976,
  // height(26,1, 0-49)
    4.941255, 4.945621, 4.949628, 4.95329, 4.956614, 4.959611, 4.962287, 
    4.96465, 4.966698, 4.96844, 4.96988, 4.971029, 4.971907, 4.972544, 
    4.972975, 4.97282, 4.973508, 4.973464, 4.973378, 4.973377, 4.973534, 
    4.974285, 4.975206, 4.976415, 4.977892, 4.979619, 4.981553, 4.983666, 
    4.985904, 4.988244, 4.990533, 4.993175, 4.995648, 4.997859, 4.999695, 
    5.00104, 5.001753, 5.001679, 5.000646, 4.998471, 4.994966, 4.989946, 
    4.983253, 4.97478, 4.964502, 4.952498, 4.938988, 4.924335, 4.909052, 
    4.893767,
  // height(26,2, 0-49)
    4.942569, 4.946893, 4.950846, 4.954443, 4.957692, 4.960606, 4.963196, 
    4.965467, 4.967426, 4.969079, 4.970437, 4.971511, 4.972326, 4.97291, 
    4.973302, 4.972916, 4.973806, 4.973686, 4.973504, 4.973412, 4.973489, 
    4.974351, 4.975346, 4.976624, 4.978158, 4.979918, 4.981861, 4.983953, 
    4.986146, 4.988422, 4.990607, 4.993344, 4.995931, 4.998283, 5.000306, 
    5.001887, 5.002901, 5.0032, 5.002613, 5.00096, 4.998045, 4.993671, 
    4.987662, 4.979883, 4.970272, 4.958864, 4.945834, 4.931497, 4.916326, 
    4.900925,
  // height(26,3, 0-49)
    4.943935, 4.948204, 4.952092, 4.955615, 4.958785, 4.961618, 4.964122, 
    4.966311, 4.968189, 4.969768, 4.97106, 4.97208, 4.972853, 4.973409, 
    4.973786, 4.973205, 4.974256, 4.974084, 4.97383, 4.973662, 4.973668, 
    4.974619, 4.975657, 4.976962, 4.978502, 4.98025, 4.982156, 4.984193, 
    4.986302, 4.988472, 4.990499, 4.99326, 4.995889, 4.99831, 5.000443, 
    5.002193, 5.003439, 5.004045, 5.003849, 5.002671, 5.000317, 4.996583, 
    4.991277, 4.984245, 4.975389, 4.964705, 4.952313, 4.938476, 4.923614, 
    4.908288,
  // height(26,4, 0-49)
    4.945349, 4.949549, 4.953363, 4.956806, 4.959896, 4.962646, 4.96507, 
    4.967181, 4.96899, 4.970509, 4.97175, 4.972735, 4.973485, 4.974032, 
    4.974418, 4.973681, 4.974834, 4.974633, 4.974329, 4.974107, 4.97405, 
    4.975069, 4.976121, 4.977407, 4.978909, 4.980601, 4.982437, 4.984389, 
    4.986394, 4.988424, 4.990258, 4.992982, 4.995586, 4.998013, 5.000195, 
    5.002046, 5.003461, 5.004312, 5.004447, 5.003695, 5.001862, 4.998744, 
    4.994145, 4.987888, 4.979846, 4.969979, 4.958351, 4.945166, 4.930783, 
    4.915707,
  // height(26,5, 0-49)
    4.946802, 4.950924, 4.954657, 4.958016, 4.961022, 4.96369, 4.966037, 
    4.968078, 4.969824, 4.971294, 4.9725, 4.973464, 4.974208, 4.974766, 
    4.975174, 4.974328, 4.975505, 4.975296, 4.974972, 4.974713, 4.974607, 
    4.97567, 4.976707, 4.977932, 4.979356, 4.980954, 4.982691, 4.984538, 
    4.986431, 4.988306, 4.989924, 4.992555, 4.995082, 4.997459, 4.999632, 
    5.001528, 5.003053, 5.004092, 5.004505, 5.004128, 5.002773, 5.000243, 
    4.996334, 4.99086, 4.983668, 4.974679, 4.963905, 4.951492, 4.937729, 
    4.923054,
  // height(26,6, 0-49)
    4.948296, 4.952331, 4.955975, 4.959248, 4.962167, 4.964754, 4.967025, 
    4.969, 4.97069, 4.972117, 4.973296, 4.974251, 4.975002, 4.975583, 
    4.976024, 4.975116, 4.97623, 4.976032, 4.975711, 4.975441, 4.975303, 
    4.976385, 4.977377, 4.978502, 4.979811, 4.981283, 4.982903, 4.984636, 
    4.986417, 4.988131, 4.989528, 4.992019, 4.994424, 4.996704, 4.998821, 
    5.000714, 5.002299, 5.003477, 5.004117, 5.004066, 5.00315, 5.001173, 
    4.997931, 4.99323, 4.986898, 4.978821, 4.968964, 4.957409, 4.944374, 
    4.930231,
  // height(26,7, 0-49)
    4.949835, 4.953774, 4.957324, 4.960505, 4.963335, 4.965837, 4.968033, 
    4.96994, 4.971579, 4.972966, 4.974124, 4.975074, 4.97584, 4.976448, 
    4.976927, 4.976012, 4.976964, 4.976792, 4.976501, 4.976244, 4.976095, 
    4.977169, 4.97809, 4.97908, 4.980241, 4.981565, 4.983052, 4.984669, 
    4.986344, 4.987903, 4.98909, 4.991405, 4.993648, 4.995795, 4.997818, 
    4.999667, 5.001273, 5.002547, 5.003373, 5.003607, 5.003088, 5.001628, 
    4.999024, 4.995079, 4.989602, 4.982448, 4.97354, 4.962898, 4.950672, 
    4.93716,
  // height(26,8, 0-49)
    4.951429, 4.955265, 4.958713, 4.961794, 4.96453, 4.966943, 4.969059, 
    4.970898, 4.97248, 4.97383, 4.974967, 4.975914, 4.976696, 4.977333, 
    4.977845, 4.976974, 4.97766, 4.977527, 4.977291, 4.977073, 4.976935, 
    4.977974, 4.978799, 4.979623, 4.980614, 4.98177, 4.983119, 4.98462, 
    4.986207, 4.987626, 4.988623, 4.99073, 4.992783, 4.994769, 4.996668, 
    4.998445, 5.000041, 5.001379, 5.002355, 5.002841, 5.002684, 5.001705, 
    4.99971, 4.99649, 4.991849, 4.985611, 4.97766, 4.967961, 4.956597, 
    4.943792,
  // height(26,9, 0-49)
    4.953088, 4.956812, 4.96015, 4.963123, 4.965757, 4.968074, 4.970102, 
    4.971866, 4.973389, 4.974695, 4.975805, 4.976745, 4.977537, 4.978196, 
    4.978734, 4.97796, 4.97827, 4.978189, 4.978033, 4.97788, 4.97778, 
    4.978755, 4.97946, 4.980095, 4.980895, 4.981874, 4.98308, 4.984471, 
    4.985987, 4.987292, 4.988131, 4.990008, 4.991851, 4.993655, 4.995411, 
    4.997094, 4.998659, 5.000037, 5.00114, 5.001849, 5.002026, 5.001497, 
    5.000074, 4.99755, 4.993714, 4.988372, 4.981369, 4.972619, 4.962144, 
    4.950095,
  // height(26,10, 0-49)
    4.954827, 4.958428, 4.961646, 4.964502, 4.967022, 4.969234, 4.971165, 
    4.972841, 4.974293, 4.975544, 4.97662, 4.977544, 4.978334, 4.979006, 
    4.979555, 4.97893, 4.97875, 4.978733, 4.978679, 4.978618, 4.978583, 
    4.979466, 4.980032, 4.980456, 4.981056, 4.981851, 4.982915, 4.984207, 
    4.985671, 4.986889, 4.987614, 4.989247, 4.990867, 4.992477, 4.99408, 
    4.995658, 4.997178, 4.998582, 4.999794, 5.000707, 5.001192, 5.001086, 
    5.000204, 4.998339, 4.995272, 4.990792, 4.98471, 4.976898, 4.967317, 
    4.956054,
  // height(26,11, 0-49)
    4.956657, 4.960123, 4.963208, 4.965933, 4.968327, 4.970419, 4.972239, 
    4.973818, 4.975185, 4.976367, 4.977395, 4.978288, 4.979064, 4.97973, 
    4.980277, 4.979839, 4.979058, 4.979119, 4.979188, 4.979247, 4.979304, 
    4.980065, 4.980476, 4.980678, 4.981071, 4.981682, 4.982608, 4.983808, 
    4.985242, 4.986406, 4.987069, 4.98845, 4.989841, 4.991255, 4.992701, 
    4.994172, 4.995643, 4.997068, 4.998378, 4.99948, 5.000252, 5.000543, 
    5.00017, 4.998927, 4.996589, 4.992929, 4.987732, 4.98083, 4.972133, 
    4.961664,
  // height(26,12, 0-49)
    4.958586, 4.961901, 4.964838, 4.967417, 4.96967, 4.971628, 4.973322, 
    4.974786, 4.976053, 4.977152, 4.978113, 4.978957, 4.9797, 4.980344, 
    4.98087, 4.980648, 4.979154, 4.979307, 4.979526, 4.97973, 4.979906, 
    4.980518, 4.980759, 4.980734, 4.980921, 4.981354, 4.982149, 4.983266, 
    4.984689, 4.985831, 4.986491, 4.987618, 4.988783, 4.990006, 4.9913, 
    4.992667, 4.994092, 4.995536, 4.996943, 4.998224, 4.99927, 4.999934, 
    5.000038, 4.999378, 4.997725, 4.994837, 4.990478, 4.984446, 4.976607, 
    4.966925,
  // height(26,13, 0-49)
    4.960617, 4.963764, 4.966533, 4.968949, 4.971044, 4.97285, 4.974402, 
    4.975734, 4.976882, 4.97788, 4.978757, 4.979533, 4.980224, 4.980828, 
    4.981322, 4.981328, 4.979001, 4.979272, 4.979662, 4.980037, 4.98036, 
    4.980793, 4.980856, 4.980605, 4.980595, 4.980857, 4.981531, 4.982577, 
    4.984003, 4.985156, 4.985874, 4.986757, 4.987704, 4.988744, 4.989898, 
    4.991172, 4.992559, 4.994028, 4.99553, 4.996988, 4.998293, 4.999307, 
    4.999858, 4.999741, 4.998724, 4.996556, 4.992984, 4.987775, 4.980757, 
    4.971845,
  // height(26,14, 0-49)
    4.962743, 4.965701, 4.968283, 4.970517, 4.972435, 4.974072, 4.975463, 
    4.976647, 4.977662, 4.978541, 4.979313, 4.980003, 4.980623, 4.981172, 
    4.981625, 4.981853, 4.978575, 4.978984, 4.97957, 4.980143, 4.980638, 
    4.980866, 4.980747, 4.980277, 4.980084, 4.980192, 4.980755, 4.98174, 
    4.983183, 4.984377, 4.985216, 4.985863, 4.986608, 4.987482, 4.988513, 
    4.989711, 4.991073, 4.992577, 4.994179, 4.995807, 4.99736, 4.998702, 
    4.999669, 5.000055, 4.999626, 4.998124, 4.995279, 4.99084, 4.984598, 
    4.976427,
  // height(26,15, 0-49)
    4.96495, 4.967693, 4.970068, 4.972099, 4.973822, 4.975271, 4.976488, 
    4.977509, 4.978373, 4.979118, 4.979771, 4.980357, 4.980891, 4.98137, 
    4.981779, 4.982203, 4.977856, 4.978431, 4.979234, 4.980026, 4.980718, 
    4.98072, 4.98042, 4.979746, 4.97939, 4.979363, 4.979831, 4.980763, 
    4.982235, 4.983498, 4.984517, 4.984947, 4.985507, 4.986237, 4.987163, 
    4.988302, 4.989655, 4.991206, 4.992913, 4.99471, 4.996499, 4.998151, 
    4.999502, 5.000349, 5.000455, 4.999561, 4.997384, 4.993657, 4.98814, 
    4.980677,
  // height(26,16, 0-49)
    4.967216, 4.969719, 4.971859, 4.973665, 4.975173, 4.97642, 4.977448, 
    4.978295, 4.979, 4.979597, 4.98012, 4.98059, 4.981026, 4.981429, 4.98179, 
    4.98237, 4.976842, 4.977604, 4.978645, 4.979676, 4.980588, 4.980343, 
    4.979868, 4.979012, 4.978518, 4.978383, 4.978773, 4.979663, 4.981173, 
    4.982527, 4.983779, 4.984013, 4.984412, 4.98502, 4.985863, 4.986963, 
    4.988326, 4.989933, 4.991749, 4.993711, 4.995725, 4.997665, 4.999369, 
    5.000635, 5.001229, 5.000884, 4.999315, 4.996238, 4.991397, 4.984601,
  // height(26,17, 0-49)
    4.969512, 4.97174, 4.973618, 4.975176, 4.976452, 4.977484, 4.978314, 
    4.97898, 4.979518, 4.979966, 4.980352, 4.980701, 4.981031, 4.981352, 
    4.981671, 4.982362, 4.975548, 4.976512, 4.977801, 4.979086, 4.980233, 
    4.979731, 4.979088, 4.978076, 4.977477, 4.977263, 4.977597, 4.978462, 
    4.980017, 4.981482, 4.98301, 4.983071, 4.983333, 4.983841, 4.984626, 
    4.985706, 4.987091, 4.988766, 4.990695, 4.99282, 4.995048, 4.997253, 
    4.999278, 5.000922, 5.001952, 5.002101, 5.001079, 4.998593, 4.994374, 
    4.988206,
  // height(26,18, 0-49)
    4.971802, 4.973717, 4.975297, 4.976582, 4.977609, 4.978417, 4.979047, 
    4.979535, 4.979914, 4.980217, 4.98047, 4.980698, 4.980921, 4.981159, 
    4.981435, 4.982197, 4.974019, 4.975191, 4.976727, 4.978267, 4.979657, 
    4.978886, 4.978089, 4.97695, 4.976281, 4.976023, 4.97633, 4.977189, 
    4.978799, 4.980386, 4.982221, 4.982135, 4.982282, 4.982712, 4.983455, 
    4.984532, 4.985951, 4.9877, 4.989746, 4.992026, 4.994454, 4.996904, 
    4.999218, 5.001203, 5.002622, 5.003211, 5.00268, 5.00073, 4.99708, 
    4.991498,
  // height(26,19, 0-49)
    4.974044, 4.975593, 4.976839, 4.977823, 4.978588, 4.979169, 4.979604, 
    4.979926, 4.980161, 4.980335, 4.98047, 4.980588, 4.98071, 4.980864, 
    4.981096, 4.981905, 4.972337, 4.973706, 4.975469, 4.977249, 4.978876, 
    4.977831, 4.976893, 4.975658, 4.974956, 4.974691, 4.975004, 4.975879, 
    4.977556, 4.979274, 4.981433, 4.981222, 4.981273, 4.981641, 4.982354, 
    4.983438, 4.984897, 4.986722, 4.98888, 4.991309, 4.993922, 4.996593, 
    4.999171, 5.001457, 5.003224, 5.004207, 5.004115, 5.00265, 4.999523, 
    4.994492,
  // height(26,20, 0-49)
    4.977043, 4.979004, 4.980653, 4.982024, 4.983145, 4.984046, 4.984755, 
    4.985302, 4.985719, 4.986032, 4.986275, 4.986479, 4.986677, 4.986904, 
    4.987205, 0, 4.969875, 4.971127, 4.972816, 4.974531, 4.976083, 4.974407, 
    4.972915, 4.971169, 4.97008, 4.969584, 4.969836, 4.970838, 4.972848, 
    4.975082, 4.978014, 4.978158, 4.978577, 4.979314, 4.980385, 4.981804, 
    4.983576, 4.985689, 4.988112, 4.990792, 4.993645, 4.996556, 4.999379, 
    5.001928, 5.003983, 5.005283, 5.005549, 5.004485, 5.001798, 4.997241,
  // height(26,21, 0-49)
    4.97925, 4.980883, 4.98223, 4.983332, 4.984216, 4.984912, 4.985448, 
    4.985849, 4.986141, 4.98635, 4.9865, 4.986621, 4.986745, 4.986916, 
    4.987184, 0, 4.965111, 4.966493, 4.968369, 4.970301, 4.97207, 4.970103, 
    4.968467, 4.966664, 4.965661, 4.965364, 4.965918, 4.967295, 4.969753, 
    4.972483, 4.976055, 4.976404, 4.977072, 4.978096, 4.979475, 4.981217, 
    4.983313, 4.985742, 4.988464, 4.991421, 4.994527, 4.997666, 5.000692, 
    5.003428, 5.005657, 5.007132, 5.007581, 5.006714, 5.004252, 4.999951,
  // height(26,22, 0-49)
    4.981404, 4.982722, 4.983783, 4.984627, 4.985284, 4.985783, 4.986148, 
    4.986403, 4.986568, 4.986663, 4.986715, 4.986749, 4.986797, 4.986908, 
    4.98714, 0, 4.96099, 4.962482, 4.964514, 4.966624, 4.968567, 4.966304, 
    4.964496, 4.962591, 4.961608, 4.961434, 4.962199, 4.963859, 4.966667, 
    4.969792, 4.973887, 4.974385, 4.975251, 4.976512, 4.978163, 4.980196, 
    4.982597, 4.985335, 4.988364, 4.991613, 4.994995, 4.998389, 5.00165, 
    5.004604, 5.007035, 5.008707, 5.009351, 5.008693, 5.006459, 5.002415,
  // height(26,23, 0-49)
    4.983479, 4.984495, 4.985284, 4.985883, 4.986323, 4.986632, 4.986832, 
    4.98694, 4.986977, 4.986959, 4.986909, 4.98685, 4.986816, 4.986859, 
    4.987047, 0, 4.957404, 4.958957, 4.961073, 4.96328, 4.965307, 4.962757, 
    4.96076, 4.958724, 4.957712, 4.957599, 4.958509, 4.960382, 4.963464, 
    4.966908, 4.971419, 4.972058, 4.973106, 4.974591, 4.9765, 4.978821, 
    4.981529, 4.984586, 4.987936, 4.991505, 4.995192, 4.998876, 5.002409, 
    5.00561, 5.008269, 5.010154, 5.011004, 5.010548, 5.008529, 5.004719,
  // height(26,24, 0-49)
    4.985459, 4.986189, 4.98672, 4.987087, 4.98732, 4.987445, 4.987481, 
    4.987444, 4.987351, 4.987216, 4.987059, 4.986901, 4.986779, 4.986742, 
    4.986866, 0, 4.954684, 4.956232, 4.958356, 4.960571, 4.962602, 4.959841, 
    4.957701, 4.955566, 4.954525, 4.954449, 4.955456, 4.957479, 4.960763, 
    4.964447, 4.969274, 4.970074, 4.971316, 4.973023, 4.975178, 4.977761, 
    4.980742, 4.984078, 4.98771, 4.991553, 4.995505, 4.999441, 5.003209, 
    5.006629, 5.009492, 5.011566, 5.012599, 5.012326, 5.010496, 5.006893,
  // height(26,25, 0-49)
    4.987332, 4.987795, 4.988081, 4.988227, 4.98826, 4.988207, 4.988082, 
    4.987899, 4.987672, 4.987413, 4.98714, 4.986873, 4.986648, 4.986516, 
    4.986553, 0, 4.952617, 4.954093, 4.956138, 4.958269, 4.960216, 4.957344, 
    4.955132, 4.95296, 4.95192, 4.951881, 4.952963, 4.955096, 4.958523, 
    4.962382, 4.96742, 4.968424, 4.96989, 4.971837, 4.974241, 4.977078, 
    4.980317, 4.983906, 4.987782, 4.991862, 4.996039, 5.000186, 5.004151, 
    5.007753, 5.010787, 5.013021, 5.014207, 5.014087, 5.012415, 5.008984,
  // height(26,26, 0-49)
    4.989085, 4.989303, 4.989362, 4.989299, 4.989142, 4.988912, 4.988623, 
    4.988289, 4.987917, 4.98752, 4.987116, 4.986723, 4.986379, 4.986131, 
    4.986053, 0, 4.951242, 4.952576, 4.954455, 4.95641, 4.958189, 4.955317, 
    4.953111, 4.950973, 4.949968, 4.949975, 4.951116, 4.953321, 4.956832, 
    4.960795, 4.965936, 4.967187, 4.96891, 4.971114, 4.973774, 4.976858, 
    4.980333, 4.984146, 4.988233, 4.992505, 4.996861, 5.001172, 5.005288, 
    5.009029, 5.012194, 5.014551, 5.015856, 5.015856, 5.014309, 5.011011,
  // height(26,27, 0-49)
    4.990705, 4.990705, 4.990558, 4.990302, 4.989961, 4.989553, 4.989096, 
    4.988595, 4.988062, 4.987507, 4.986948, 4.986408, 4.985921, 4.985535, 
    4.985317, 0, 4.950675, 4.9518, 4.953434, 4.955128, 4.956655, 4.953875, 
    4.951737, 4.949679, 4.948724, 4.948766, 4.949928, 4.952152, 4.955673, 
    4.959657, 4.964782, 4.966302, 4.968293, 4.970756, 4.97366, 4.976973, 
    4.980659, 4.984664, 4.988923, 4.993354, 4.997853, 5.002294, 5.00653, 
    5.010384, 5.013654, 5.016113, 5.017517, 5.017615, 5.016166, 5.012967,
  // height(26,28, 0-49)
    4.992178, 4.991997, 4.991673, 4.991239, 4.990721, 4.990136, 4.989495, 
    4.988809, 4.988087, 4.987344, 4.9866, 4.985881, 4.985225, 4.984678, 
    4.984301, 0, 4.951277, 4.95214, 4.953459, 4.954813, 4.956015, 4.953386, 
    4.95134, 4.949368, 4.948436, 4.948458, 4.949565, 4.951716, 4.955142, 
    4.959041, 4.964017, 4.965793, 4.968029, 4.970719, 4.973828, 4.977328, 
    4.981176, 4.985326, 4.989712, 4.994259, 4.998865, 5.003407, 5.007742, 
    5.011695, 5.015062, 5.017617, 5.019115, 5.019303, 5.017936, 5.014811,
  // height(26,29, 0-49)
    4.993492, 4.993173, 4.992706, 4.992117, 4.991431, 4.990662, 4.989821, 
    4.98892, 4.987972, 4.987, 4.986029, 4.985097, 4.984242, 4.98352, 
    4.982977, 0, 4.952824, 4.953395, 4.954348, 4.955293, 4.95609, 4.953598, 
    4.951597, 4.949647, 4.948653, 4.948557, 4.949506, 4.951476, 4.95469, 
    4.958384, 4.963066, 4.965036, 4.967458, 4.970321, 4.97359, 4.977238, 
    4.981226, 4.985511, 4.990031, 4.994714, 4.999458, 5.004147, 5.00863, 
    5.012733, 5.016247, 5.018942, 5.020564, 5.020856, 5.019571, 5.016503,
  // height(26,30, 0-49)
    4.99386, 4.992723, 4.991463, 4.990121, 4.988725, 4.987293, 4.985828, 
    4.984329, 4.982784, 4.98118, 4.979504, 4.977741, 4.975895, 4.973988, 
    4.972077, 4.969747, 4.956999, 4.956827, 4.957161, 4.957656, 4.958186, 
    4.95614, 4.954606, 4.953129, 4.952481, 4.952558, 4.953475, 4.955208, 
    4.957977, 4.961077, 4.964963, 4.966609, 4.968697, 4.971236, 4.974212, 
    4.977611, 4.981407, 4.985562, 4.990018, 4.994699, 4.999503, 5.004301, 
    5.008934, 5.013212, 5.016919, 5.019805, 5.021607, 5.022055, 5.020894, 
    5.017915,
  // height(26,31, 0-49)
    4.994776, 4.99362, 4.992315, 4.990895, 4.989389, 4.987814, 4.986178, 
    4.984484, 4.982728, 4.980905, 4.979011, 4.977039, 4.974996, 4.972894, 
    4.97077, 4.969105, 4.957089, 4.956472, 4.956341, 4.956375, 4.956476, 
    4.954564, 4.953073, 4.951636, 4.950986, 4.951061, 4.95199, 4.953743, 
    4.956496, 4.959546, 4.963222, 4.965158, 4.96754, 4.970372, 4.973639, 
    4.977323, 4.981398, 4.985823, 4.99054, 4.995468, 5.000506, 5.005515, 
    5.010334, 5.014765, 5.01858, 5.021528, 5.023334, 5.023723, 5.022443, 
    5.01929,
  // height(26,32, 0-49)
    4.995375, 4.994205, 4.99286, 4.991376, 4.989777, 4.988082, 4.986303, 
    4.984447, 4.982514, 4.980509, 4.978431, 4.976282, 4.974068, 4.971794, 
    4.969482, 4.968209, 4.95724, 4.956205, 4.955632, 4.955235, 4.954943, 
    4.953212, 4.951815, 4.950471, 4.949865, 4.949964, 4.950908, 4.952662, 
    4.955353, 4.958293, 4.961698, 4.963876, 4.966497, 4.969563, 4.973063, 
    4.976978, 4.981282, 4.985934, 4.990874, 4.996023, 5.001267, 5.006473, 
    5.011462, 5.016034, 5.019948, 5.022943, 5.024738, 5.025053, 5.023633, 
    5.020279,
  // height(26,33, 0-49)
    4.995639, 4.99447, 4.9931, 4.991568, 4.989897, 4.988105, 4.98621, 
    4.984221, 4.982143, 4.979988, 4.97776, 4.975465, 4.973111, 4.970702, 
    4.968242, 4.967098, 4.957392, 4.955994, 4.955024, 4.954244, 4.95361, 
    4.952107, 4.950858, 4.949664, 4.949143, 4.949293, 4.950252, 4.951982, 
    4.954559, 4.957333, 4.960416, 4.962787, 4.965594, 4.96884, 4.972515, 
    4.976605, 4.981087, 4.985918, 4.991039, 4.996368, 5.001789, 5.007158, 
    5.012293, 5.01698, 5.020972, 5.023992, 5.025752, 5.025967, 5.02438, 
    5.020803,
  // height(26,34, 0-49)
    4.995543, 4.994396, 4.993027, 4.99147, 4.98975, 4.98789, 4.985905, 
    4.983811, 4.98162, 4.979345, 4.976997, 4.97459, 4.97213, 4.969624, 
    4.967066, 4.965834, 4.957517, 4.955821, 4.954513, 4.953405, 4.952485, 
    4.951245, 4.95019, 4.9492, 4.948807, 4.949031, 4.950005, 4.951681, 
    4.954097, 4.956656, 4.959386, 4.961906, 4.964849, 4.968222, 4.972019, 
    4.97623, 4.980836, 4.985796, 4.991051, 4.996513, 5.002068, 5.007562, 
    5.012805, 5.017571, 5.021602, 5.024612, 5.026301, 5.026382, 5.024599, 
    5.020772,
  // height(26,35, 0-49)
    4.995066, 4.99397, 4.992628, 4.991074, 4.989336, 4.987434, 4.985391, 
    4.983224, 4.98095, 4.978586, 4.976151, 4.97366, 4.971129, 4.968563, 
    4.965956, 4.964484, 4.957617, 4.955689, 4.954103, 4.952727, 4.951577, 
    4.950626, 4.949806, 4.949069, 4.948839, 4.949157, 4.950138, 4.951736, 
    4.953943, 4.956252, 4.958614, 4.961243, 4.964278, 4.967728, 4.971596, 
    4.975876, 4.980554, 4.985588, 4.990923, 4.996468, 5.002102, 5.007667, 
    5.012964, 5.017759, 5.02178, 5.024729, 5.026304, 5.026208, 5.024194, 
    5.02009,
  // height(26,36, 0-49)
    4.99419, 4.993175, 4.991889, 4.99037, 4.988643, 4.986734, 4.984667, 
    4.98246, 4.980136, 4.977716, 4.975226, 4.972688, 4.970117, 4.967527, 
    4.964915, 4.96312, 4.957703, 4.95561, 4.953803, 4.952217, 4.950887, 
    4.950241, 4.949687, 4.949242, 4.949209, 4.949636, 4.95062, 4.952115, 
    4.954077, 4.95611, 4.958105, 4.960808, 4.963894, 4.967376, 4.971268, 
    4.975566, 4.98026, 4.985313, 4.990666, 4.996232, 5.001882, 5.007453, 
    5.012741, 5.017495, 5.021441, 5.024268, 5.025669, 5.02535, 5.023067, 
    5.018667,
  // height(26,37, 0-49)
    4.992908, 4.991998, 4.9908, 4.989348, 4.987668, 4.985786, 4.983728, 
    4.981519, 4.979182, 4.976744, 4.974233, 4.971678, 4.969099, 4.966518, 
    4.963937, 4.961798, 4.957793, 4.955594, 4.953619, 4.951871, 4.950411, 
    4.950073, 4.949806, 4.949687, 4.949876, 4.950426, 4.951407, 4.952781, 
    4.954471, 4.956215, 4.957856, 4.9606, 4.963703, 4.967181, 4.971049, 
    4.975317, 4.979972, 4.984982, 4.990291, 4.995806, 5.001399, 5.006898, 
    5.012094, 5.01673, 5.020518, 5.023149, 5.024311, 5.023713, 5.021127, 
    5.016415,
  // height(26,38, 0-49)
    4.991222, 4.990443, 4.98936, 4.988006, 4.986406, 4.984589, 4.98258, 
    4.980407, 4.978095, 4.975675, 4.97318, 4.970641, 4.968087, 4.965544, 
    4.963021, 4.960566, 4.957904, 4.955646, 4.953547, 4.951684, 4.950138, 
    4.950104, 4.950134, 4.950362, 4.950793, 4.951478, 4.952455, 4.953692, 
    4.955092, 4.956546, 4.957858, 4.960621, 4.96371, 4.967146, 4.970952, 
    4.975142, 4.979702, 4.98461, 4.989802, 4.995189, 5.000639, 5.005978, 
    5.010987, 5.015409, 5.01895, 5.021299, 5.022146, 5.021213, 5.018287, 
    5.013258,
  // height(26,39, 0-49)
    4.989146, 4.988517, 4.987576, 4.98635, 4.984865, 4.983149, 4.981227, 
    4.979128, 4.976882, 4.974522, 4.972079, 4.969591, 4.967091, 4.96461, 
    4.962165, 4.959454, 4.95805, 4.955768, 4.953585, 4.951646, 4.950048, 
    4.950306, 4.950636, 4.951224, 4.951909, 4.952735, 4.953708, 4.954801, 
    4.955904, 4.957078, 4.958095, 4.960857, 4.963908, 4.967274, 4.970981, 
    4.975045, 4.979459, 4.984196, 4.9892, 4.994374, 4.999588, 5.004664, 
    5.009383, 5.013483, 5.016672, 5.018644, 5.019099, 5.017773, 5.014479, 
    5.009132,
  // height(26,40, 0-49)
    4.986707, 4.986245, 4.985466, 4.984396, 4.983058, 4.981478, 4.979682, 
    4.977698, 4.975558, 4.973294, 4.970941, 4.968537, 4.966121, 4.963724, 
    4.961371, 4.958483, 4.95824, 4.95596, 4.953722, 4.951737, 4.950122, 
    4.950653, 4.951275, 4.952221, 4.953166, 4.954142, 4.955109, 4.956059, 
    4.956869, 4.957781, 4.958541, 4.961287, 4.964283, 4.967553, 4.97113, 
    4.975026, 4.979239, 4.983742, 4.988476, 4.993349, 4.998224, 5.002929, 
    5.007241, 5.010903, 5.013631, 5.015126, 5.015107, 5.013333, 5.009647, 
    5.004004,
  // height(26,41, 0-49)
    4.983946, 4.983662, 4.983064, 4.982172, 4.981009, 4.979598, 4.977962, 
    4.976132, 4.974137, 4.972007, 4.969779, 4.967493, 4.965187, 4.962894, 
    4.960647, 4.957664, 4.958471, 4.956212, 4.953946, 4.951943, 4.950333, 
    4.951114, 4.952014, 4.953312, 4.954513, 4.955637, 4.9566, 4.957409, 
    4.957942, 4.95862, 4.959163, 4.961884, 4.964809, 4.967964, 4.97138, 
    4.97507, 4.97903, 4.983232, 4.987618, 4.992094, 4.996525, 5.000741, 
    5.004525, 5.007628, 5.009777, 5.010693, 5.010121, 5.007853, 5.003766, 
    4.997855,
  // height(26,42, 0-49)
    4.980917, 4.980814, 4.98041, 4.979715, 4.978751, 4.977537, 4.976097, 
    4.974453, 4.972636, 4.970678, 4.968611, 4.966472, 4.964302, 4.962132, 
    4.959999, 4.957001, 4.958748, 4.95652, 4.954246, 4.952245, 4.950657, 
    4.95166, 4.952818, 4.954448, 4.955894, 4.957162, 4.958123, 4.958803, 
    4.95908, 4.959553, 4.959918, 4.962606, 4.965451, 4.968475, 4.971704, 
    4.97515, 4.978807, 4.982642, 4.986598, 4.990582, 4.994461, 4.998068, 
    5.0012, 5.003619, 5.005074, 5.005314, 5.004117, 5.001315, 4.996832, 
    4.990704,
  // height(26,43, 0-49)
    4.977679, 4.97776, 4.977554, 4.977072, 4.976327, 4.975336, 4.974116, 
    4.972692, 4.971086, 4.969328, 4.967451, 4.965489, 4.963478, 4.961449, 
    4.959437, 4.956493, 4.959065, 4.956875, 4.954607, 4.952624, 4.951071, 
    4.952264, 4.953651, 4.955585, 4.95726, 4.958661, 4.959623, 4.960185, 
    4.960233, 4.960534, 4.960759, 4.963408, 4.966163, 4.96904, 4.97206, 
    4.975228, 4.978531, 4.981936, 4.985381, 4.988777, 4.991995, 4.994875, 
    4.99723, 4.998845, 4.999496, 4.998971, 4.997089, 4.993732, 4.988872, 
    4.982594,
  // height(26,44, 0-49)
    4.974301, 4.974561, 4.974557, 4.974297, 4.973784, 4.973035, 4.972059, 
    4.970877, 4.96951, 4.967981, 4.966322, 4.964559, 4.962726, 4.960854, 
    4.958971, 4.956134, 4.959414, 4.957269, 4.955017, 4.953065, 4.951551, 
    4.952901, 4.954484, 4.956686, 4.958561, 4.960083, 4.961043, 4.961501, 
    4.961351, 4.961507, 4.961627, 4.964231, 4.966889, 4.969604, 4.972392, 
    4.975247, 4.97815, 4.981063, 4.983919, 4.986634, 4.989085, 4.991127, 
    4.992589, 4.993289, 4.99304, 4.991673, 4.989062, 4.985146, 4.979949, 
    4.973607,
  // height(26,45, 0-49)
    4.970855, 4.971286, 4.971483, 4.971446, 4.971176, 4.970679, 4.969965, 
    4.969045, 4.967938, 4.96666, 4.965239, 4.963696, 4.962062, 4.960358, 
    4.958611, 4.955917, 4.95979, 4.957693, 4.955468, 4.95355, 4.952076, 
    4.95355, 4.955291, 4.957713, 4.959756, 4.961379, 4.962333, 4.9627, 
    4.962382, 4.962423, 4.96246, 4.965011, 4.967559, 4.970098, 4.972632, 
    4.97514, 4.977598, 4.979958, 4.982154, 4.984101, 4.985687, 4.986785, 
    4.987253, 4.986942, 4.985713, 4.983451, 4.980091, 4.975633, 4.970161, 
    4.963855,
  // height(26,46, 0-49)
    4.967414, 4.968003, 4.968394, 4.968578, 4.968554, 4.968318, 4.967876, 
    4.967232, 4.9664, 4.96539, 4.964222, 4.962915, 4.961491, 4.959968, 
    4.958365, 4.955836, 4.960183, 4.95814, 4.955951, 4.954069, 4.952631, 
    4.954192, 4.956049, 4.95864, 4.960809, 4.962502, 4.963447, 4.963733, 
    4.963276, 4.963221, 4.963187, 4.965672, 4.968098, 4.970442, 4.972695, 
    4.974825, 4.976792, 4.978544, 4.980013, 4.981115, 4.981754, 4.981822, 
    4.98121, 4.979815, 4.977552, 4.974366, 4.970264, 4.965308, 4.959643, 
    4.953489,
  // height(26,47, 0-49)
    4.964046, 4.964777, 4.965352, 4.965752, 4.96597, 4.965997, 4.965829, 
    4.96547, 4.96492, 4.964187, 4.963284, 4.962223, 4.961019, 4.959685, 
    4.958235, 4.955878, 4.960584, 4.958601, 4.956454, 4.954607, 4.953197, 
    4.954808, 4.956738, 4.959435, 4.961684, 4.963416, 4.964339, 4.964552, 
    4.96398, 4.963842, 4.963738, 4.966136, 4.968418, 4.970546, 4.972489, 
    4.974205, 4.975642, 4.976735, 4.977419, 4.977613, 4.977237, 4.976211, 
    4.974462, 4.97194, 4.968619, 4.964515, 4.959707, 4.954324, 4.948567, 
    4.942689,
  // height(26,48, 0-49)
    4.96081, 4.961668, 4.962411, 4.963017, 4.963469, 4.963753, 4.96386, 
    4.963782, 4.963516, 4.963064, 4.962431, 4.961621, 4.960644, 4.959507, 
    4.958216, 4.956029, 4.960979, 4.959066, 4.956965, 4.955151, 4.953761, 
    4.955386, 4.957339, 4.960083, 4.962356, 4.964089, 4.964973, 4.965117, 
    4.964446, 4.964223, 4.964039, 4.966322, 4.968429, 4.970309, 4.971912, 
    4.973177, 4.974042, 4.974437, 4.974288, 4.973528, 4.972093, 4.969935, 
    4.967025, 4.963368, 4.959004, 4.954024, 4.948578, 4.942863, 4.937129, 
    4.93166,
  // height(26,49, 0-49)
    4.957191, 4.958059, 4.958873, 4.959602, 4.960219, 4.9607, 4.961027, 
    4.961179, 4.961144, 4.960912, 4.960473, 4.959821, 4.95895, 4.957851, 
    4.956515, 4.953525, 4.964903, 4.962058, 4.958658, 4.955644, 4.953284, 
    4.956749, 4.960586, 4.965696, 4.969499, 4.971891, 4.972278, 4.970906, 
    4.967642, 4.965106, 4.962541, 4.964893, 4.966942, 4.968615, 4.969858, 
    4.970594, 4.970757, 4.97027, 4.969067, 4.967099, 4.964337, 4.960783, 
    4.956475, 4.951499, 4.945994, 4.940145, 4.934196, 4.928425, 4.923135, 
    4.918625,
  // height(27,0, 0-49)
    4.952485, 4.956017, 4.95919, 4.962013, 4.964487, 4.966623, 4.968421, 
    4.969888, 4.971034, 4.971874, 4.972427, 4.972726, 4.972806, 4.972714, 
    4.972504, 4.972033, 4.971988, 4.9717, 4.971503, 4.971475, 4.971662, 
    4.97227, 4.973104, 4.974205, 4.975557, 4.977133, 4.978898, 4.980816, 
    4.982846, 4.984953, 4.987058, 4.989343, 4.991569, 4.993695, 4.995677, 
    4.997463, 4.998989, 5.00017, 5.000906, 5.001068, 5.000506, 4.999043, 
    4.996487, 4.992639, 4.987311, 4.98035, 4.971671, 4.961278, 4.9493, 
    4.936006,
  // height(27,1, 0-49)
    4.953785, 4.957267, 4.960383, 4.963142, 4.965549, 4.967614, 4.969344, 
    4.970743, 4.971827, 4.97261, 4.973116, 4.973373, 4.973421, 4.973308, 
    4.973083, 4.972408, 4.972571, 4.972211, 4.971914, 4.971784, 4.971873, 
    4.97256, 4.97343, 4.974563, 4.975933, 4.977504, 4.979235, 4.981091, 
    4.983034, 4.985042, 4.987011, 4.989357, 4.991658, 4.993884, 4.995999, 
    4.997962, 4.999713, 5.001177, 5.002253, 5.002817, 5.002716, 5.001765, 
    4.999763, 4.996496, 4.991755, 4.985361, 4.977194, 4.967225, 4.955546, 
    4.942395,
  // height(27,2, 0-49)
    4.9551, 4.958522, 4.961576, 4.964267, 4.96661, 4.96861, 4.970279, 
    4.971625, 4.97266, 4.973405, 4.97388, 4.974118, 4.974155, 4.974039, 
    4.97382, 4.972966, 4.973311, 4.972891, 4.972506, 4.972278, 4.972264, 
    4.973009, 4.97389, 4.975019, 4.976368, 4.9779, 4.979566, 4.981339, 
    4.983176, 4.985064, 4.98687, 4.989237, 4.991573, 4.993855, 4.996058, 
    4.998144, 5.000066, 5.00175, 5.003102, 5.003998, 5.004288, 5.003786, 
    5.002285, 4.999563, 4.995397, 4.989588, 4.981988, 4.972539, 4.961292, 
    4.948447,
  // height(27,3, 0-49)
    4.956424, 4.959782, 4.962767, 4.965392, 4.967669, 4.969612, 4.971227, 
    4.972527, 4.973528, 4.974247, 4.97471, 4.974946, 4.974991, 4.974892, 
    4.974695, 4.973688, 4.974173, 4.973708, 4.973245, 4.972928, 4.972816, 
    4.973597, 4.974463, 4.975552, 4.976844, 4.978302, 4.979884, 4.981561, 
    4.983288, 4.985043, 4.986671, 4.989024, 4.991359, 4.993658, 4.995905, 
    4.99807, 5.000108, 5.001954, 5.003517, 5.004678, 5.00529, 5.005171, 
    5.004114, 5.001892, 4.998278, 4.993056, 4.986063, 4.977203, 4.966496, 
    4.9541,
  // height(27,4, 0-49)
    4.957763, 4.961049, 4.963962, 4.966518, 4.968731, 4.970614, 4.97218, 
    4.973444, 4.974419, 4.975125, 4.975588, 4.975837, 4.975906, 4.975838, 
    4.975676, 4.974549, 4.975114, 4.974617, 4.974098, 4.973704, 4.973499, 
    4.974296, 4.97512, 4.976135, 4.977338, 4.978698, 4.980179, 4.981754, 
    4.983374, 4.984993, 4.986437, 4.988748, 4.991049, 4.993332, 4.995584, 
    4.997785, 4.999891, 5.001845, 5.003561, 5.004924, 5.005792, 5.005991, 
    5.00532, 5.003553, 5.000459, 4.995819, 4.98945, 4.981233, 4.971154, 
    4.959323,
  // height(27,5, 0-49)
    4.959124, 4.96233, 4.965165, 4.967649, 4.969796, 4.971621, 4.973139, 
    4.974367, 4.975321, 4.976024, 4.976496, 4.976768, 4.976871, 4.976844, 
    4.976726, 4.975518, 4.976087, 4.975574, 4.975018, 4.974565, 4.97428, 
    4.975071, 4.975831, 4.976738, 4.977826, 4.979064, 4.980437, 4.981911, 
    4.983433, 4.984925, 4.986189, 4.988428, 4.990667, 4.992902, 4.995128, 
    4.997325, 4.999457, 5.001471, 5.003284, 5.004794, 5.005862, 5.006324, 
    5.005984, 5.004626, 5.002022, 4.997947, 4.992211, 4.984674, 4.975287, 
    4.964118,
  // height(27,6, 0-49)
    4.960515, 4.963633, 4.966385, 4.96879, 4.970866, 4.972629, 4.974098, 
    4.975291, 4.976225, 4.976924, 4.97741, 4.977711, 4.977855, 4.977876, 
    4.977808, 4.976558, 4.977046, 4.976531, 4.97596, 4.975471, 4.975124, 
    4.975888, 4.976562, 4.977334, 4.978279, 4.979381, 4.980637, 4.982016, 
    4.983459, 4.984834, 4.985934, 4.988077, 4.990227, 4.992387, 4.994555, 
    4.996716, 4.998837, 5.000868, 5.002738, 5.004347, 5.005566, 5.006243, 
    5.006188, 5.005199, 5.003053, 4.999527, 4.994426, 4.987591, 4.978942, 
    4.968504,
  // height(27,7, 0-49)
    4.961944, 4.964969, 4.96763, 4.969948, 4.971945, 4.97364, 4.975054, 
    4.976207, 4.977119, 4.977812, 4.978312, 4.978641, 4.978827, 4.978899, 
    4.97888, 4.977633, 4.977947, 4.977446, 4.976884, 4.976382, 4.975995, 
    4.976711, 4.97728, 4.977891, 4.978675, 4.97963, 4.980768, 4.982057, 
    4.98344, 4.984717, 4.985673, 4.987694, 4.989734, 4.991795, 4.99388, 
    4.995977, 4.998057, 5.000075, 5.001965, 5.003634, 5.004968, 5.005818, 
    5.006014, 5.00536, 5.003646, 5.000652, 4.996178, 4.990054, 4.982172, 
    4.972516,
  // height(27,8, 0-49)
    4.96342, 4.966343, 4.968904, 4.971127, 4.973035, 4.974654, 4.976002, 
    4.977108, 4.977989, 4.978671, 4.979177, 4.979532, 4.979758, 4.979877, 
    4.979905, 4.978708, 4.978746, 4.978274, 4.97775, 4.977262, 4.976861, 
    4.977507, 4.977953, 4.978384, 4.978992, 4.979788, 4.980811, 4.982022, 
    4.983364, 4.984567, 4.985405, 4.987285, 4.989192, 4.991133, 4.993113, 
    4.995123, 4.997139, 4.999117, 5.001001, 5.002707, 5.004125, 5.005124, 
    5.005543, 5.005198, 5.003892, 5.001414, 4.997559, 4.992144, 4.985043, 
    4.976196,
  // height(27,9, 0-49)
    4.964952, 4.967762, 4.970212, 4.972329, 4.974138, 4.975667, 4.976941, 
    4.977984, 4.978825, 4.979486, 4.97999, 4.980362, 4.98062, 4.980781, 
    4.980847, 4.979746, 4.979405, 4.97898, 4.978518, 4.978075, 4.977688, 
    4.978245, 4.978553, 4.978786, 4.97921, 4.979844, 4.980752, 4.981893, 
    4.983215, 4.984366, 4.985122, 4.98684, 4.988597, 4.990402, 4.992261, 
    4.994167, 4.9961, 4.998025, 4.999886, 5.001608, 5.003094, 5.004222, 
    5.004846, 5.004794, 5.003879, 5.001898, 4.998647, 4.993936, 4.987614, 
    4.979589,
  // height(27,10, 0-49)
    4.966544, 4.969228, 4.971554, 4.973551, 4.975248, 4.976675, 4.977859, 
    4.97883, 4.979616, 4.980243, 4.980734, 4.981112, 4.98139, 4.981582, 
    4.981678, 4.980717, 4.979891, 4.979529, 4.979159, 4.978791, 4.978449, 
    4.978896, 4.979054, 4.97908, 4.979313, 4.979784, 4.980581, 4.981661, 
    4.982981, 4.984105, 4.984818, 4.986358, 4.987952, 4.989606, 4.991331, 
    4.993123, 4.994964, 4.996823, 4.998651, 5.000382, 5.001927, 5.003174, 
    5.003991, 5.00422, 5.003681, 5.002182, 4.999519, 4.995496, 4.989943, 
    4.982737,
  // height(27,11, 0-49)
    4.968184, 4.970732, 4.972922, 4.974787, 4.976358, 4.97767, 4.978752, 
    4.979636, 4.980354, 4.980931, 4.981393, 4.981763, 4.982052, 4.982261, 
    4.982378, 4.981594, 4.980174, 4.979899, 4.979648, 4.979387, 4.979123, 
    4.979436, 4.979437, 4.979248, 4.979291, 4.979603, 4.980292, 4.981318, 
    4.98265, 4.983774, 4.984485, 4.985836, 4.987253, 4.988749, 4.990333, 
    4.992004, 4.993749, 4.995539, 4.997333, 4.99907, 5.000671, 5.002034, 
    5.00304, 5.00354, 5.003365, 5.00233, 5.000237, 4.996881, 4.992076, 
    4.985673,
  // height(27,12, 0-49)
    4.969869, 4.972264, 4.974305, 4.976025, 4.977458, 4.978641, 4.979606, 
    4.98039, 4.981024, 4.981538, 4.981959, 4.982306, 4.982589, 4.982803, 
    4.982933, 4.982355, 4.980234, 4.98007, 4.979968, 4.979845, 4.979689, 
    4.97985, 4.979685, 4.979283, 4.979139, 4.979298, 4.979885, 4.980863, 
    4.982218, 4.983363, 4.984119, 4.985269, 4.986504, 4.987836, 4.989278, 
    4.990828, 4.992476, 4.9942, 4.995962, 4.997709, 4.999368, 5.000849, 
    5.002039, 5.002804, 5.002984, 5.002398, 5.00085, 4.998134, 4.99405, 
    4.988423,
  // height(27,13, 0-49)
    4.971578, 4.973805, 4.975684, 4.977247, 4.978529, 4.979571, 4.980408, 
    4.98108, 4.981618, 4.982056, 4.982419, 4.982728, 4.982991, 4.983199, 
    4.983337, 4.982982, 4.980053, 4.980028, 4.980104, 4.980148, 4.980134, 
    4.980123, 4.97979, 4.979178, 4.978858, 4.978872, 4.979362, 4.980295, 
    4.981681, 4.982868, 4.983716, 4.984661, 4.98571, 4.986878, 4.988178, 
    4.989611, 4.991169, 4.992833, 4.994571, 4.996334, 4.998056, 4.999658, 
    5.001034, 5.002057, 5.002578, 5.002422, 5.001395, 4.999288, 4.995888, 
    4.991003,
  // height(27,14, 0-49)
    4.973285, 4.975332, 4.977035, 4.978428, 4.979551, 4.980443, 4.981143, 
    4.981692, 4.982125, 4.982474, 4.982768, 4.983025, 4.983253, 4.983449, 
    4.983591, 4.983465, 4.979623, 4.979764, 4.980047, 4.980291, 4.980448, 
    4.980245, 4.979743, 4.978934, 4.978452, 4.978334, 4.978735, 4.979624, 
    4.981044, 4.98229, 4.983274, 4.984014, 4.98488, 4.985888, 4.987052, 
    4.988374, 4.98985, 4.991462, 4.993183, 4.994971, 4.996765, 4.998491, 
    5.000052, 5.001328, 5.002178, 5.002431, 5.001897, 5.000363, 4.99761, 
    4.993423,
  // height(27,15, 0-49)
    4.974969, 4.976818, 4.97833, 4.979544, 4.980499, 4.981234, 4.981791, 
    4.982209, 4.982529, 4.98278, 4.982994, 4.983189, 4.983375, 4.983549, 
    4.983696, 4.983794, 4.978942, 4.979278, 4.979795, 4.980265, 4.98062, 
    4.980211, 4.979545, 4.978554, 4.977929, 4.977694, 4.978014, 4.978863, 
    4.980318, 4.981638, 4.982798, 4.983336, 4.984023, 4.984879, 4.985915, 
    4.987135, 4.988539, 4.990111, 4.991827, 4.993648, 4.99552, 4.997373, 
    4.999117, 5.000638, 5.001802, 5.002442, 5.002368, 5.00137, 4.999219, 
    4.995688,
  // height(27,16, 0-49)
    4.9766, 4.978232, 4.979541, 4.980565, 4.981343, 4.981917, 4.982327, 
    4.982615, 4.982817, 4.982967, 4.983095, 4.98322, 4.983356, 4.983504, 
    4.983661, 4.983968, 4.978021, 4.978576, 4.979346, 4.980065, 4.980643, 
    4.980015, 4.979194, 4.97804, 4.977294, 4.976964, 4.977215, 4.978029, 
    4.979517, 4.980919, 4.982292, 4.982636, 4.983153, 4.983865, 4.984783, 
    4.985914, 4.987255, 4.988797, 4.990517, 4.992379, 4.994334, 4.996316, 
    4.99824, 4.999999, 5.001459, 5.002461, 5.002818, 5.002316, 5.000722, 
    4.997799,
  // height(27,17, 0-49)
    4.97815, 4.979545, 4.980634, 4.981458, 4.982053, 4.982463, 4.982728, 
    4.982884, 4.982973, 4.983024, 4.983063, 4.983118, 4.983199, 4.983321, 
    4.983489, 4.983988, 4.976887, 4.977677, 4.978717, 4.979698, 4.980515, 
    4.97966, 4.978692, 4.977397, 4.976559, 4.976156, 4.976355, 4.977139, 
    4.97866, 4.980151, 4.981763, 4.981924, 4.982281, 4.982859, 4.983669, 
    4.98472, 4.986009, 4.987531, 4.989263, 4.991172, 4.993215, 4.995326, 
    4.997425, 4.999409, 5.001151, 5.00249, 5.003245, 5.0032, 5.002119, 
    4.999754,
  // height(27,18, 0-49)
    4.979592, 4.980724, 4.981576, 4.982186, 4.982595, 4.982841, 4.982964, 
    4.983, 4.982983, 4.982941, 4.9829, 4.982886, 4.982915, 4.983007, 
    4.983186, 4.983865, 4.975588, 4.976619, 4.977927, 4.979177, 4.980241, 
    4.979152, 4.978045, 4.976635, 4.97573, 4.975284, 4.975449, 4.976212, 
    4.977769, 4.979352, 4.981221, 4.981211, 4.981418, 4.981871, 4.982583, 
    4.983562, 4.984807, 4.986314, 4.988064, 4.990025, 4.992156, 4.994394, 
    4.996664, 4.998864, 5.000867, 5.002522, 5.003644, 5.004018, 5.003407, 
    5.001557,
  // height(27,19, 0-49)
    4.980903, 4.98174, 4.98233, 4.982714, 4.982932, 4.983019, 4.98301, 
    4.982938, 4.982831, 4.982711, 4.982603, 4.982526, 4.982506, 4.982572, 
    4.982763, 4.983617, 4.9742, 4.975467, 4.977031, 4.978539, 4.979841, 
    4.978513, 4.97728, 4.975773, 4.974828, 4.974364, 4.974518, 4.975278, 
    4.976873, 4.978549, 4.980679, 4.98051, 4.980577, 4.980914, 4.981531, 
    4.982439, 4.983643, 4.985138, 4.986907, 4.988921, 4.991139, 4.993503, 
    4.995936, 4.998341, 5.000593, 5.002542, 5.004004, 5.004765, 5.004586, 
    5.00321,
  // height(27,20, 0-49)
    4.982862, 4.984146, 4.985185, 4.986007, 4.98664, 4.987111, 4.987448, 
    4.987677, 4.987826, 4.987921, 4.987986, 4.988048, 4.988135, 4.988278, 
    4.988526, 0, 4.972143, 4.973258, 4.97473, 4.976183, 4.977445, 4.975578, 
    4.973876, 4.971932, 4.970649, 4.969963, 4.970038, 4.970872, 4.97272, 
    4.974809, 4.977582, 4.977671, 4.978006, 4.978611, 4.979485, 4.980634, 
    4.982059, 4.983755, 4.985709, 4.987898, 4.990287, 4.992825, 4.995441, 
    4.998047, 5.000524, 5.002726, 5.004475, 5.005559, 5.005739, 5.004762,
  // height(27,21, 0-49)
    4.984021, 4.985055, 4.985878, 4.986519, 4.987, 4.98735, 4.987592, 
    4.987746, 4.987836, 4.987881, 4.987903, 4.987926, 4.987977, 4.98809, 
    4.988317, 0, 4.96787, 4.969113, 4.970778, 4.972454, 4.973938, 4.971829, 
    4.970017, 4.96804, 4.966849, 4.966359, 4.966709, 4.967876, 4.970111, 
    4.97262, 4.975931, 4.976147, 4.976643, 4.977433, 4.978511, 4.979876, 
    4.981517, 4.983426, 4.985584, 4.987966, 4.990533, 4.993235, 4.996002, 
    4.998747, 5.001359, 5.003693, 5.005579, 5.006813, 5.007162, 5.006378,
  // height(27,22, 0-49)
    4.9851, 4.985905, 4.986529, 4.987001, 4.987345, 4.987583, 4.987735, 
    4.987818, 4.987849, 4.987846, 4.987824, 4.987807, 4.987818, 4.987895, 
    4.988095, 0, 4.96427, 4.965615, 4.967438, 4.969296, 4.970961, 4.968601, 
    4.96665, 4.964593, 4.963428, 4.963049, 4.963583, 4.964988, 4.96751, 
    4.970334, 4.974064, 4.974349, 4.974948, 4.975873, 4.977114, 4.978661, 
    4.980502, 4.982621, 4.984995, 4.987593, 4.990371, 4.993275, 4.996236, 
    4.999167, 5.001956, 5.004463, 5.006518, 5.007926, 5.008459, 5.007876,
  // height(27,23, 0-49)
    4.986108, 4.986693, 4.987132, 4.98745, 4.987665, 4.987799, 4.987868, 
    4.987884, 4.987857, 4.987806, 4.987741, 4.98768, 4.987649, 4.987686, 
    4.987846, 0, 4.961174, 4.962575, 4.964491, 4.966458, 4.968225, 4.965626, 
    4.963521, 4.961361, 4.960176, 4.959849, 4.960501, 4.962069, 4.964801, 
    4.96786, 4.971903, 4.972238, 4.972919, 4.973962, 4.97535, 4.977074, 
    4.979115, 4.981455, 4.984063, 4.986903, 4.989927, 4.993075, 4.996275, 
    4.999434, 5.00244, 5.005151, 5.007399, 5.008994, 5.009711, 5.00932,
  // height(27,24, 0-49)
    4.987052, 4.987432, 4.987696, 4.987866, 4.987962, 4.987997, 4.987984, 
    4.987933, 4.987851, 4.98775, 4.987639, 4.987533, 4.987454, 4.987441, 
    4.987548, 0, 4.958886, 4.960289, 4.962229, 4.964231, 4.966028, 4.963264, 
    4.961052, 4.958817, 4.957613, 4.957313, 4.958032, 4.959703, 4.962571, 
    4.965787, 4.970043, 4.970445, 4.971216, 4.972371, 4.973891, 4.975769, 
    4.977979, 4.980506, 4.983313, 4.986362, 4.989601, 4.992966, 4.996381, 
    4.99975, 5.002959, 5.005866, 5.0083, 5.010072, 5.010966, 5.010753,
  // height(27,25, 0-49)
    4.987951, 4.988135, 4.988231, 4.988259, 4.988237, 4.988174, 4.98808, 
    4.987959, 4.987818, 4.987662, 4.987497, 4.987339, 4.987206, 4.987133, 
    4.987175, 0, 4.957164, 4.958512, 4.960404, 4.962363, 4.964118, 4.961286, 
    4.959035, 4.956786, 4.955588, 4.955317, 4.956082, 4.957819, 4.960765, 
    4.964076, 4.968446, 4.968953, 4.969841, 4.971123, 4.972783, 4.974807, 
    4.977177, 4.979869, 4.98285, 4.986078, 4.989499, 4.993052, 4.996652, 
    5.000207, 5.003596, 5.006678, 5.009283, 5.011218, 5.01227, 5.012215,
  // height(27,26, 0-49)
    4.988813, 4.988812, 4.98875, 4.988639, 4.9885, 4.988336, 4.988153, 
    4.987953, 4.987741, 4.987518, 4.98729, 4.987069, 4.986872, 4.986731, 
    4.986691, 0, 4.956017, 4.957257, 4.959034, 4.960871, 4.962512, 4.95972, 
    4.957509, 4.955312, 4.954154, 4.953917, 4.954714, 4.956479, 4.959447, 
    4.962788, 4.967175, 4.967828, 4.968863, 4.970294, 4.972103, 4.974275, 
    4.976792, 4.979629, 4.982756, 4.986129, 4.989699, 4.9934, 4.997152, 
    5.000857, 5.004397, 5.007628, 5.010381, 5.01246, 5.013651, 5.013734,
  // height(27,27, 0-49)
    4.98965, 4.989479, 4.989264, 4.98902, 4.988759, 4.988484, 4.9882, 
    4.987906, 4.987603, 4.987295, 4.986986, 4.986688, 4.986415, 4.986197, 
    4.986067, 0, 4.955529, 4.956617, 4.958216, 4.959864, 4.961324, 4.958663, 
    4.956551, 4.954452, 4.95335, 4.953136, 4.95393, 4.955672, 4.958594, 
    4.961887, 4.966184, 4.967004, 4.968203, 4.969788, 4.971744, 4.974054, 
    4.976701, 4.979663, 4.98291, 4.986403, 4.990092, 4.993917, 4.997795, 
    5.001633, 5.005309, 5.008677, 5.011567, 5.013782, 5.015105, 5.01531,
  // height(27,28, 0-49)
    4.990469, 4.990145, 4.989788, 4.989411, 4.989022, 4.988625, 4.988218, 
    4.987805, 4.987385, 4.986967, 4.986554, 4.98616, 4.985801, 4.9855, 
    4.985283, 0, 4.956028, 4.956934, 4.958307, 4.959707, 4.96093, 4.958463, 
    4.956476, 4.954484, 4.953412, 4.953169, 4.953884, 4.955516, 4.958292, 
    4.961439, 4.965523, 4.966502, 4.967848, 4.969568, 4.971642, 4.974057, 
    4.976798, 4.979848, 4.983181, 4.986762, 4.990545, 4.994473, 4.998466, 
    5.002428, 5.006239, 5.009749, 5.012783, 5.015139, 5.016596, 5.016923,
  // height(27,29, 0-49)
    4.991272, 4.99082, 4.990334, 4.989828, 4.989304, 4.988763, 4.988209, 
    4.987643, 4.987072, 4.986504, 4.985958, 4.985448, 4.984994, 4.984619, 
    4.984338, 0, 4.957261, 4.957983, 4.959101, 4.960205, 4.96113, 4.958851, 
    4.956955, 4.955013, 4.953891, 4.953528, 4.954064, 4.955482, 4.958002, 
    4.960886, 4.964627, 4.965713, 4.967158, 4.968967, 4.971126, 4.973623, 
    4.976449, 4.979589, 4.983022, 4.986718, 4.990633, 4.994709, 4.998869, 
    5.003012, 5.00701, 5.010713, 5.013935, 5.016467, 5.018081, 5.018536,
  // height(27,30, 0-49)
    4.991342, 4.990104, 4.98886, 4.987627, 4.986415, 4.985223, 4.984044, 
    4.982868, 4.981678, 4.980457, 4.979197, 4.977892, 4.976555, 4.975228, 
    4.973989, 4.972118, 4.961142, 4.961493, 4.962195, 4.962931, 4.963588, 
    4.961671, 4.96014, 4.958567, 4.957699, 4.957439, 4.957901, 4.95906, 
    4.961126, 4.963423, 4.966387, 4.96713, 4.968222, 4.969685, 4.971525, 
    4.973748, 4.976355, 4.979339, 4.982685, 4.986363, 4.990328, 4.994513, 
    4.998833, 5.003178, 5.007408, 5.011355, 5.014824, 5.017593, 5.019419, 
    5.020052,
  // height(27,31, 0-49)
    4.992085, 4.990796, 4.989485, 4.988165, 4.986845, 4.985525, 4.9842, 
    4.982865, 4.981511, 4.980129, 4.978714, 4.977267, 4.975796, 4.974329, 
    4.972923, 4.971511, 4.96095, 4.960932, 4.961246, 4.961601, 4.961905, 
    4.960153, 4.958697, 4.957186, 4.956329, 4.956063, 4.956516, 4.957662, 
    4.959669, 4.961869, 4.964588, 4.965552, 4.966871, 4.968566, 4.970642, 
    4.973103, 4.975951, 4.979178, 4.982767, 4.986686, 4.990888, 4.995302, 
    4.99984, 5.004383, 5.008787, 5.012877, 5.016449, 5.019275, 5.021107, 
    5.021693,
  // height(27,32, 0-49)
    4.992704, 4.991362, 4.989981, 4.988571, 4.987143, 4.985699, 4.984235, 
    4.982752, 4.981244, 4.979711, 4.978148, 4.976559, 4.974949, 4.97334, 
    4.971759, 4.970668, 4.96088, 4.960486, 4.96041, 4.960387, 4.96035, 
    4.958791, 4.957444, 4.956033, 4.955215, 4.954963, 4.95541, 4.956527, 
    4.958438, 4.960497, 4.962925, 4.964082, 4.965597, 4.967487, 4.969763, 
    4.972429, 4.975488, 4.97893, 4.982742, 4.986887, 4.991313, 4.995951, 
    5.000702, 5.005444, 5.010021, 5.014254, 5.017927, 5.020806, 5.022637, 
    5.023165,
  // height(27,33, 0-49)
    4.993176, 4.991786, 4.990337, 4.988843, 4.987313, 4.98575, 4.984156, 
    4.982533, 4.980882, 4.979203, 4.977501, 4.975778, 4.97404, 4.972296, 
    4.97056, 4.969613, 4.960853, 4.960111, 4.959667, 4.95929, 4.95894, 
    4.957603, 4.956401, 4.955134, 4.954391, 4.954172, 4.954613, 4.955681, 
    4.957458, 4.959333, 4.961436, 4.962754, 4.964429, 4.966482, 4.968922, 
    4.971757, 4.974994, 4.978625, 4.982632, 4.986979, 4.991614, 4.996459, 
    5.001411, 5.006339, 5.011081, 5.015445, 5.019209, 5.022128, 5.023943, 
    5.024394,
  // height(27,34, 0-49)
    4.993468, 4.992046, 4.990543, 4.988973, 4.98735, 4.985679, 4.983964, 
    4.982211, 4.980426, 4.978615, 4.976783, 4.974936, 4.973081, 4.971223, 
    4.96936, 4.968389, 4.960826, 4.959777, 4.958998, 4.958305, 4.957679, 
    4.956588, 4.955568, 4.954486, 4.953852, 4.953686, 4.95412, 4.955118, 
    4.956721, 4.958376, 4.960136, 4.961588, 4.963395, 4.965575, 4.968145, 
    4.971118, 4.974501, 4.978288, 4.98246, 4.986983, 4.9918, 4.996827, 
    5.001957, 5.00705, 5.011934, 5.016407, 5.020238, 5.023174, 5.024948, 
    5.025294,
  // height(27,35, 0-49)
    4.993543, 4.992109, 4.990572, 4.988945, 4.987246, 4.98548, 4.983659, 
    4.98179, 4.979885, 4.977952, 4.976004, 4.97405, 4.972095, 4.970143, 
    4.968186, 4.967057, 4.960784, 4.959477, 4.958406, 4.957438, 4.956577, 
    4.955748, 4.954938, 4.954085, 4.953589, 4.953495, 4.953919, 4.954828, 
    4.956221, 4.957632, 4.959045, 4.960607, 4.962515, 4.964794, 4.967463, 
    4.970541, 4.974034, 4.977944, 4.982249, 4.986913, 4.991876, 4.997052, 
    5.002326, 5.007547, 5.012538, 5.017087, 5.020951, 5.023866, 5.025561, 
    5.025771,
  // height(27,36, 0-49)
    4.993363, 4.991943, 4.990395, 4.988733, 4.986978, 4.985139, 4.983231, 
    4.981265, 4.979257, 4.977222, 4.975175, 4.973129, 4.971095, 4.969073, 
    4.967054, 4.965679, 4.960728, 4.959213, 4.957893, 4.956695, 4.95564, 
    4.955082, 4.954507, 4.953914, 4.953588, 4.953581, 4.953995, 4.954797, 
    4.955952, 4.957104, 4.958177, 4.959828, 4.961814, 4.964163, 4.966903, 
    4.970053, 4.973625, 4.977619, 4.982017, 4.986782, 4.991848, 4.997127, 
    5.002496, 5.007801, 5.012851, 5.017424, 5.021269, 5.024117, 5.025689, 
    5.025723,
  // height(27,37, 0-49)
    4.992894, 4.991515, 4.989983, 4.988314, 4.986529, 4.984643, 4.982672, 
    4.980633, 4.978547, 4.97643, 4.974305, 4.972188, 4.970094, 4.968026, 
    4.965975, 4.964311, 4.960664, 4.958989, 4.957465, 4.956078, 4.95487, 
    4.954582, 4.954257, 4.953956, 4.953823, 4.953918, 4.954322, 4.955003, 
    4.955902, 4.956789, 4.957542, 4.959267, 4.961312, 4.963708, 4.96649, 
    4.969682, 4.973296, 4.977336, 4.981783, 4.986598, 4.991717, 4.997042, 
    5.00245, 5.007774, 5.01282, 5.017355, 5.021121, 5.02384, 5.025236, 
    5.025045,
  // height(27,38, 0-49)
    4.992102, 4.990796, 4.989309, 4.987664, 4.985879, 4.983975, 4.981972, 
    4.979889, 4.977752, 4.97558, 4.973402, 4.971236, 4.969102, 4.967009, 
    4.964951, 4.962999, 4.960605, 4.958811, 4.957121, 4.955583, 4.954257, 
    4.954235, 4.954173, 4.954182, 4.954263, 4.954476, 4.954871, 4.955422, 
    4.956054, 4.956684, 4.957149, 4.958934, 4.961021, 4.963445, 4.966245, 
    4.969447, 4.97307, 4.977113, 4.981561, 4.986373, 4.991481, 4.996788, 
    5.002161, 5.007431, 5.012395, 5.016815, 5.020426, 5.022949, 5.024106, 
    5.023642,
  // height(27,39, 0-49)
    4.990971, 4.989764, 4.988355, 4.986764, 4.985014, 4.983126, 4.981123, 
    4.97903, 4.976871, 4.974676, 4.97247, 4.970282, 4.968132, 4.966033, 
    4.963985, 4.961775, 4.960558, 4.95868, 4.956858, 4.955204, 4.953793, 
    4.954025, 4.954226, 4.954561, 4.954874, 4.955217, 4.955606, 4.956029, 
    4.956393, 4.956779, 4.956996, 4.958832, 4.960948, 4.963384, 4.966179, 
    4.969365, 4.972958, 4.976961, 4.981358, 4.986107, 4.991138, 4.99635, 
    5.001607, 5.006737, 5.011529, 5.015744, 5.019113, 5.021358, 5.022209, 
    5.021421,
  // height(27,40, 0-49)
    4.989492, 4.988411, 4.987108, 4.985605, 4.983923, 4.982087, 4.980121, 
    4.978053, 4.975909, 4.973721, 4.971519, 4.969333, 4.96719, 4.965103, 
    4.963079, 4.960662, 4.960529, 4.958594, 4.956668, 4.954926, 4.953461, 
    4.953931, 4.954395, 4.955062, 4.955615, 4.956097, 4.956487, 4.956788, 
    4.956896, 4.957064, 4.957074, 4.958955, 4.961094, 4.963527, 4.966299, 
    4.96944, 4.972969, 4.976889, 4.98118, 4.9858, 4.990678, 4.995711, 
    5.000761, 5.005651, 5.010171, 5.01408, 5.017112, 5.018996, 5.019468, 
    5.018303,
  // height(27,41, 0-49)
    4.98767, 4.986738, 4.98557, 4.984185, 4.982606, 4.98086, 4.978968, 
    4.97696, 4.974867, 4.972721, 4.970555, 4.9684, 4.966283, 4.964226, 
    4.962235, 4.959669, 4.96052, 4.958544, 4.956538, 4.954738, 4.95324, 
    4.953933, 4.95465, 4.955646, 4.956444, 4.957076, 4.957476, 4.957663, 
    4.957536, 4.957518, 4.957366, 4.959292, 4.961448, 4.963868, 4.9666, 
    4.969671, 4.973102, 4.976892, 4.98102, 4.985444, 4.99009, 4.994852, 
    4.999594, 5.004138, 5.008276, 5.01177, 5.014363, 5.015793, 5.015814, 
    5.014226,
  // height(27,42, 0-49)
    4.985522, 4.98476, 4.983753, 4.982516, 4.981074, 4.97945, 4.977669, 
    4.975759, 4.973754, 4.971684, 4.969582, 4.967484, 4.965418, 4.963405, 
    4.961457, 4.958804, 4.960528, 4.958524, 4.956461, 4.954623, 4.953115, 
    4.954007, 4.954963, 4.956277, 4.957321, 4.958108, 4.958529, 4.958621, 
    4.958286, 4.958118, 4.957849, 4.959821, 4.961989, 4.96439, 4.967066, 
    4.970046, 4.973344, 4.976959, 4.980868, 4.985023, 4.989351, 4.993749, 
    4.998077, 5.002162, 5.005802, 5.008768, 5.010814, 5.011698, 5.011199, 
    5.009146,
  // height(27,43, 0-49)
    4.983078, 4.982504, 4.981679, 4.980618, 4.979343, 4.977874, 4.976239, 
    4.974464, 4.972579, 4.970617, 4.968614, 4.966598, 4.964602, 4.962647, 
    4.96075, 4.958064, 4.960546, 4.958526, 4.956423, 4.954565, 4.953062, 
    4.954131, 4.955307, 4.956923, 4.958204, 4.959147, 4.959601, 4.959621, 
    4.959113, 4.958833, 4.958492, 4.960511, 4.962692, 4.965067, 4.967675, 
    4.97054, 4.973672, 4.977067, 4.980697, 4.984512, 4.988438, 4.992373, 
    4.996177, 4.999687, 5.00271, 5.00503, 5.006423, 5.006673, 5.005592, 
    5.003043,
  // height(27,44, 0-49)
    4.980382, 4.980007, 4.979383, 4.978521, 4.97744, 4.976157, 4.974699, 
    4.973089, 4.971357, 4.969535, 4.967654, 4.965747, 4.963842, 4.961959, 
    4.960116, 4.957444, 4.96057, 4.958542, 4.956412, 4.954548, 4.953062, 
    4.954283, 4.955656, 4.957548, 4.959053, 4.960151, 4.960651, 4.960621, 
    4.959981, 4.95963, 4.959256, 4.961325, 4.963518, 4.965861, 4.968388, 
    4.971116, 4.974051, 4.97718, 4.980473, 4.983876, 4.987314, 4.990685, 
    4.993859, 4.996679, 4.998967, 5.000529, 5.001168, 5.000703, 4.998985, 
    4.995923,
  // height(27,45, 0-49)
    4.977487, 4.977318, 4.976908, 4.976263, 4.975397, 4.974328, 4.973073, 
    4.971658, 4.970108, 4.968452, 4.96672, 4.964941, 4.963143, 4.961346, 
    4.959565, 4.956938, 4.960594, 4.958564, 4.956421, 4.954561, 4.953098, 
    4.954445, 4.955987, 4.958123, 4.959834, 4.961078, 4.961632, 4.961581, 
    4.960852, 4.960466, 4.960093, 4.962214, 4.964419, 4.966725, 4.969159, 
    4.971728, 4.974432, 4.977252, 4.980149, 4.983069, 4.985935, 4.988648, 
    4.991086, 4.993104, 4.994545, 4.995243, 4.995037, 4.993789, 4.991396, 
    4.987819,
  // height(27,46, 0-49)
    4.974452, 4.974493, 4.974304, 4.97389, 4.973258, 4.972421, 4.971393, 
    4.970196, 4.968852, 4.967385, 4.965823, 4.964191, 4.962515, 4.960814, 
    4.959103, 4.956544, 4.960613, 4.958589, 4.956441, 4.954591, 4.953156, 
    4.954598, 4.956281, 4.95862, 4.960506, 4.961886, 4.962506, 4.96246, 
    4.961684, 4.961299, 4.960954, 4.963126, 4.965339, 4.9676, 4.969926, 
    4.972314, 4.974755, 4.97722, 4.979667, 4.982036, 4.98425, 4.986214, 
    4.987817, 4.988932, 4.989427, 4.989168, 4.988042, 4.98596, 4.982873, 
    4.9788,
  // height(27,47, 0-49)
    4.971342, 4.971589, 4.971627, 4.971451, 4.971065, 4.970476, 4.969693, 
    4.968733, 4.967612, 4.966353, 4.964977, 4.963507, 4.961967, 4.960371, 
    4.958735, 4.956259, 4.960622, 4.95861, 4.956469, 4.954632, 4.953219, 
    4.954731, 4.956517, 4.959014, 4.961045, 4.962544, 4.963233, 4.963216, 
    4.962434, 4.962078, 4.961781, 4.963998, 4.966213, 4.96842, 4.970622, 
    4.972805, 4.974948, 4.977016, 4.978959, 4.98071, 4.982198, 4.983331, 
    4.98401, 4.984134, 4.9836, 4.982316, 4.980217, 4.977271, 4.973495, 
    4.968967,
  // height(27,48, 0-49)
    4.968221, 4.96867, 4.968932, 4.968997, 4.968864, 4.968532, 4.968005, 
    4.967294, 4.966412, 4.965373, 4.964195, 4.962899, 4.961504, 4.960023, 
    4.958469, 4.956077, 4.960622, 4.958631, 4.9565, 4.954679, 4.953285, 
    4.954834, 4.956685, 4.959286, 4.961421, 4.963017, 4.963776, 4.963808, 
    4.963056, 4.96275, 4.962512, 4.964767, 4.96697, 4.969106, 4.971163, 
    4.973114, 4.974928, 4.976556, 4.977943, 4.97902, 4.979716, 4.979949, 
    4.979635, 4.978698, 4.977073, 4.974717, 4.971618, 4.96781, 4.963374, 
    4.958452,
  // height(27,49, 0-49)
    4.964688, 4.965261, 4.965686, 4.965944, 4.966022, 4.965912, 4.965609, 
    4.96511, 4.964419, 4.963542, 4.962485, 4.96126, 4.959875, 4.958338, 
    4.95665, 4.953324, 4.963948, 4.960972, 4.957505, 4.954463, 4.952101, 
    4.95546, 4.959188, 4.964164, 4.967905, 4.970287, 4.97073, 4.969472, 
    4.966397, 4.964046, 4.961688, 4.964251, 4.966651, 4.968855, 4.970845, 
    4.972581, 4.974022, 4.975112, 4.975787, 4.975982, 4.975631, 4.974669, 
    4.973047, 4.97073, 4.967712, 4.964019, 4.959729, 4.954966, 4.949904, 
    4.944765,
  // height(28,0, 0-49)
    4.963037, 4.965694, 4.96799, 4.96993, 4.971521, 4.972774, 4.973701, 
    4.974322, 4.97466, 4.974749, 4.974625, 4.974331, 4.973917, 4.973434, 
    4.972936, 4.972286, 4.972091, 4.971761, 4.971567, 4.971555, 4.971744, 
    4.972298, 4.973012, 4.97391, 4.974973, 4.97617, 4.977477, 4.978871, 
    4.980332, 4.981852, 4.983389, 4.985156, 4.986973, 4.988846, 4.990781, 
    4.992773, 4.99481, 4.99686, 4.998869, 5.000762, 5.002431, 5.003738, 
    5.00451, 5.00454, 5.003603, 5.00145, 4.997844, 4.992567, 4.985462, 
    4.976461,
  // height(28,1, 0-49)
    4.964329, 4.966931, 4.969166, 4.971049, 4.972588, 4.973791, 4.974676, 
    4.975263, 4.975576, 4.975647, 4.975512, 4.975218, 4.974807, 4.97433, 
    4.973841, 4.973016, 4.97299, 4.972588, 4.972288, 4.972158, 4.972225, 
    4.97281, 4.973512, 4.974387, 4.975416, 4.976565, 4.977803, 4.979111, 
    4.980468, 4.981872, 4.983257, 4.985047, 4.986896, 4.988817, 4.990819, 
    4.992906, 4.995065, 4.997271, 4.999474, 5.001599, 5.003541, 5.005161, 
    5.006287, 5.006708, 5.006192, 5.004486, 5.001334, 4.996506, 4.989824, 
    4.981192,
  // height(28,2, 0-49)
    4.965621, 4.968162, 4.970339, 4.972167, 4.973656, 4.974818, 4.975669, 
    4.976233, 4.976532, 4.976597, 4.976467, 4.976181, 4.975784, 4.975326, 
    4.974851, 4.973862, 4.973973, 4.973501, 4.973098, 4.972849, 4.972789, 
    4.973388, 4.974058, 4.974888, 4.97586, 4.976943, 4.978105, 4.979328, 
    4.98059, 4.981882, 4.983115, 4.984918, 4.986787, 4.988737, 4.990783, 
    4.992933, 4.995179, 4.997493, 4.999833, 5.002124, 5.004266, 5.00612, 
    5.007517, 5.00825, 5.008084, 5.006764, 5.004031, 4.999646, 4.993412, 
    4.985214,
  // height(28,3, 0-49)
    4.966917, 4.969394, 4.971512, 4.973285, 4.974725, 4.975849, 4.976673, 
    4.977219, 4.97751, 4.977582, 4.977464, 4.977196, 4.976823, 4.976389, 
    4.975935, 4.974799, 4.974998, 4.974462, 4.973961, 4.973601, 4.973414, 
    4.97401, 4.974627, 4.975387, 4.976283, 4.977287, 4.978371, 4.979517, 
    4.980698, 4.981891, 4.98298, 4.984787, 4.986662, 4.988626, 4.990697, 
    4.992883, 4.995177, 4.997558, 4.999983, 5.002381, 5.004653, 5.00667, 
    5.008263, 5.009232, 5.009345, 5.008354, 5.006002, 5.002043, 4.996274, 
    4.988564,
  // height(28,4, 0-49)
    4.968223, 4.970632, 4.972686, 4.974402, 4.975794, 4.97688, 4.977679, 
    4.97821, 4.978501, 4.97858, 4.978481, 4.97824, 4.977897, 4.977489, 
    4.97706, 4.975801, 4.976025, 4.975429, 4.974844, 4.97438, 4.974075, 
    4.974649, 4.975199, 4.975864, 4.976665, 4.977577, 4.978583, 4.979664, 
    4.980787, 4.981899, 4.982858, 4.984657, 4.986529, 4.988494, 4.99057, 
    4.992767, 4.99508, 4.997489, 4.999952, 5.002404, 5.004749, 5.006863, 
    5.008582, 5.00972, 5.010053, 5.009339, 5.007329, 5.00378, 4.998486, 
    4.991301,
  // height(28,5, 0-49)
    4.969545, 4.971881, 4.973867, 4.975522, 4.976862, 4.977907, 4.978678, 
    4.979195, 4.979484, 4.979575, 4.979497, 4.979285, 4.978973, 4.978598, 
    4.978193, 4.976839, 4.977013, 4.976367, 4.975714, 4.975161, 4.97475, 
    4.975285, 4.975749, 4.976297, 4.976986, 4.977798, 4.978731, 4.979761, 
    4.980849, 4.981899, 4.982753, 4.984535, 4.986391, 4.988342, 4.990406, 
    4.992593, 4.994897, 4.997301, 4.999764, 5.002223, 5.00459, 5.006744, 
    5.008537, 5.009789, 5.010285, 5.009804, 5.008102, 5.004949, 5.000133, 
    4.993503,
  // height(28,6, 0-49)
    4.970886, 4.97314, 4.975051, 4.976639, 4.977922, 4.978922, 4.979661, 
    4.98016, 4.980445, 4.980545, 4.980488, 4.980305, 4.980027, 4.979684, 
    4.979302, 4.977885, 4.977926, 4.977243, 4.97654, 4.975917, 4.975418, 
    4.975897, 4.97626, 4.976669, 4.977231, 4.977938, 4.978801, 4.979794, 
    4.980872, 4.981885, 4.982657, 4.984412, 4.986242, 4.988164, 4.990201, 
    4.992358, 4.994633, 4.997004, 4.999434, 5.001863, 5.00421, 5.006363, 
    5.008183, 5.0095, 5.010123, 5.009836, 5.008419, 5.005644, 5.001309, 
    4.995253,
  // height(28,7, 0-49)
    4.97225, 4.974414, 4.976242, 4.977755, 4.978972, 4.979918, 4.980618, 
    4.981094, 4.98137, 4.981475, 4.981435, 4.981279, 4.981033, 4.980721, 
    4.98036, 4.978918, 4.978734, 4.978028, 4.977297, 4.976627, 4.976062, 
    4.976467, 4.976714, 4.976967, 4.977389, 4.977985, 4.978783, 4.979753, 
    4.980847, 4.981849, 4.982569, 4.984282, 4.986072, 4.987955, 4.989949, 
    4.992061, 4.994284, 4.996599, 4.998971, 5.001343, 5.003639, 5.005757, 
    5.007569, 5.008923, 5.00964, 5.009525, 5.00837, 5.005964, 5.002109, 
    4.996638,
  // height(28,8, 0-49)
    4.973632, 4.975698, 4.977432, 4.978859, 4.980003, 4.980888, 4.981541, 
    4.981984, 4.982244, 4.982347, 4.98232, 4.982186, 4.981969, 4.981684, 
    4.98134, 4.979915, 4.979413, 4.978697, 4.977963, 4.977275, 4.97667, 
    4.976981, 4.977097, 4.97718, 4.977454, 4.977934, 4.978669, 4.97963, 
    4.980763, 4.981778, 4.982479, 4.984136, 4.985872, 4.987704, 4.989642, 
    4.991693, 4.99385, 4.996092, 4.998385, 5.00068, 5.002903, 5.004966, 
    5.006748, 5.008116, 5.00891, 5.00895, 5.008045, 5.005998, 5.00262, 
    4.997739,
  // height(28,9, 0-49)
    4.975026, 4.976983, 4.978614, 4.979947, 4.981006, 4.98182, 4.982415, 
    4.982818, 4.983053, 4.983148, 4.983126, 4.983008, 4.982814, 4.982553, 
    4.982228, 4.980858, 4.979939, 4.979236, 4.978528, 4.977848, 4.977229, 
    4.97743, 4.977406, 4.977305, 4.977422, 4.977784, 4.978463, 4.979421, 
    4.980612, 4.981666, 4.98238, 4.983967, 4.985638, 4.987401, 4.989273, 
    4.991251, 4.993327, 4.995483, 4.997686, 4.999889, 5.002028, 5.004021, 
    5.005765, 5.007137, 5.007996, 5.008182, 5.00752, 5.005828, 5.002922, 
    4.998632,
  // height(28,10, 0-49)
    4.976417, 4.978255, 4.979773, 4.981001, 4.981967, 4.9827, 4.98323, 
    4.983584, 4.983787, 4.983865, 4.98384, 4.983733, 4.983557, 4.983315, 
    4.983003, 4.981734, 4.980297, 4.979631, 4.978978, 4.97834, 4.977737, 
    4.977809, 4.977633, 4.977343, 4.9773, 4.977544, 4.978166, 4.979129, 
    4.980392, 4.981504, 4.982268, 4.983768, 4.985357, 4.987044, 4.988835, 
    4.990729, 4.992716, 4.994777, 4.996881, 4.998987, 5.001035, 5.002955, 
    5.004656, 5.00603, 5.006954, 5.007286, 5.006864, 5.005523, 5.003084, 
    4.999376,
  // height(28,11, 0-49)
    4.977788, 4.979498, 4.980894, 4.982008, 4.982872, 4.983517, 4.983973, 
    4.984268, 4.984429, 4.984483, 4.984451, 4.984347, 4.984181, 4.983957, 
    4.983658, 4.98253, 4.980477, 4.979874, 4.979309, 4.978745, 4.978193, 
    4.978118, 4.977784, 4.977296, 4.977094, 4.977222, 4.97779, 4.978761, 
    4.980103, 4.981291, 4.982141, 4.983537, 4.985031, 4.986626, 4.988327, 
    4.990128, 4.992017, 4.993978, 4.995981, 4.997988, 4.999948, 5.001796, 
    5.00346, 5.004842, 5.005836, 5.006314, 5.006134, 5.005139, 5.003159, 
    5.000023,
  // height(28,12, 0-49)
    4.979121, 4.98069, 4.981956, 4.982948, 4.983704, 4.984252, 4.984627, 
    4.984859, 4.984973, 4.984995, 4.984945, 4.984837, 4.984681, 4.984471, 
    4.984189, 4.983234, 4.980469, 4.979962, 4.979518, 4.979064, 4.978595, 
    4.978358, 4.977861, 4.977178, 4.976821, 4.976835, 4.97735, 4.978325, 
    4.979751, 4.981029, 4.981995, 4.983273, 4.984656, 4.986147, 4.987747, 
    4.989446, 4.991234, 4.993092, 4.994994, 4.996906, 4.998783, 5.000571, 
    5.002206, 5.003607, 5.004677, 5.00531, 5.005374, 5.004723, 5.003193, 
    5.000611,
  // height(28,13, 0-49)
    4.980392, 4.981812, 4.982938, 4.983803, 4.984443, 4.98489, 4.985179, 
    4.985341, 4.985403, 4.985387, 4.985314, 4.985199, 4.985044, 4.984848, 
    4.984589, 4.983837, 4.980271, 4.979891, 4.979608, 4.979298, 4.978949, 
    4.978534, 4.977874, 4.977001, 4.976495, 4.976401, 4.976861, 4.977839, 
    4.979345, 4.980719, 4.981833, 4.982975, 4.984235, 4.98561, 4.987098, 
    4.988689, 4.990372, 4.992128, 4.993932, 4.995756, 4.997561, 4.999301, 
    5.00092, 5.002353, 5.003514, 5.00431, 5.004621, 5.004309, 5.003215, 
    5.001168,
  // height(28,14, 0-49)
    4.981575, 4.982839, 4.983819, 4.984552, 4.985072, 4.985415, 4.985616, 
    4.985703, 4.985707, 4.98565, 4.98555, 4.985421, 4.985268, 4.985085, 
    4.984856, 4.98433, 4.97988, 4.979667, 4.979576, 4.979448, 4.979251, 
    4.97865, 4.977829, 4.976778, 4.976137, 4.975942, 4.976348, 4.97732, 
    4.978895, 4.98037, 4.981659, 4.982649, 4.98377, 4.985018, 4.986386, 
    4.987864, 4.989438, 4.991094, 4.992805, 4.99455, 4.996294, 4.998002, 
    4.999622, 5.001102, 5.002368, 5.003336, 5.003896, 5.003918, 5.003249, 
    5.001713,
  // height(28,15, 0-49)
    4.982654, 4.983751, 4.984578, 4.985173, 4.985571, 4.985808, 4.985918, 
    4.98593, 4.985873, 4.985772, 4.985643, 4.985499, 4.985344, 4.985178, 
    4.984991, 4.984704, 4.979304, 4.979292, 4.979429, 4.979517, 4.979506, 
    4.978709, 4.977736, 4.976521, 4.975759, 4.975474, 4.975827, 4.976785, 
    4.978418, 4.979989, 4.981472, 4.982297, 4.983266, 4.984376, 4.985615, 
    4.986974, 4.988441, 4.989997, 4.991624, 4.993299, 4.994998, 4.996687, 
    4.998328, 4.999872, 5.001257, 5.002406, 5.003217, 5.003567, 5.003305, 
    5.002254,
  // height(28,16, 0-49)
    4.983608, 4.984528, 4.985196, 4.98565, 4.985922, 4.986052, 4.98607, 
    4.986007, 4.98589, 4.985743, 4.985583, 4.985423, 4.985268, 4.985124, 
    4.984986, 4.984951, 4.978553, 4.978775, 4.979172, 4.979506, 4.979712, 
    4.978718, 4.977604, 4.976244, 4.975379, 4.975018, 4.975318, 4.976254, 
    4.977931, 4.979589, 4.981279, 4.981926, 4.98273, 4.983689, 4.984793, 
    4.986029, 4.987384, 4.988845, 4.990394, 4.992012, 4.993679, 4.995368, 
    4.997046, 4.998671, 5.000189, 5.001527, 5.002593, 5.003264, 5.003393, 
    5.002801,
  // height(28,17, 0-49)
    4.984422, 4.985153, 4.985654, 4.985961, 4.986106, 4.986128, 4.986056, 
    4.985919, 4.985743, 4.985553, 4.985363, 4.985186, 4.985034, 4.984914, 
    4.984838, 4.985061, 4.977653, 4.978134, 4.978813, 4.97942, 4.979869, 
    4.978677, 4.977434, 4.975953, 4.975008, 4.974584, 4.974835, 4.975744, 
    4.977448, 4.979182, 4.981081, 4.981539, 4.982168, 4.982968, 4.983927, 
    4.985033, 4.986276, 4.987643, 4.98912, 4.990694, 4.992342, 4.994048, 
    4.995781, 4.997505, 4.999168, 5.000705, 5.002026, 5.00301, 5.003512, 
    5.003355,
  // height(28,18, 0-49)
    4.985089, 4.985617, 4.985938, 4.98609, 4.986105, 4.986018, 4.985858, 
    4.985652, 4.985424, 4.985193, 4.984977, 4.984787, 4.98464, 4.984551, 
    4.984545, 4.985033, 4.976648, 4.977406, 4.978383, 4.979276, 4.979985, 
    4.978594, 4.977239, 4.975657, 4.97465, 4.974179, 4.974391, 4.975267, 
    4.976982, 4.978776, 4.980881, 4.981141, 4.981584, 4.982214, 4.98302, 
    4.983992, 4.985119, 4.986394, 4.987806, 4.989342, 4.990986, 4.992723, 
    4.994529, 4.996365, 4.998188, 4.999933, 5.00151, 5.002803, 5.003664, 
    5.003913,
  // height(28,19, 0-49)
    4.985601, 4.985903, 4.986029, 4.986017, 4.985898, 4.985704, 4.985462, 
    4.985194, 4.98492, 4.984657, 4.984419, 4.984222, 4.984084, 4.984033, 
    4.984104, 4.984866, 4.975602, 4.976647, 4.977926, 4.979109, 4.980078, 
    4.978496, 4.977036, 4.975368, 4.974319, 4.973816, 4.973994, 4.974836, 
    4.976551, 4.978387, 4.980682, 4.980737, 4.980986, 4.981435, 4.982077, 
    4.982903, 4.983911, 4.985092, 4.986441, 4.987948, 4.989601, 4.991385, 
    4.993277, 4.995243, 4.997238, 4.999198, 5.001037, 5.002635, 5.003841, 
    5.004478,
  // height(28,20, 0-49)
    4.986712, 4.987498, 4.98811, 4.988571, 4.988906, 4.989136, 4.989282, 
    4.98936, 4.98939, 4.989389, 4.989371, 4.989356, 4.989365, 4.989432, 
    4.989607, 0, 4.973971, 4.974906, 4.976127, 4.977295, 4.978267, 4.976232, 
    4.974376, 4.972327, 4.970971, 4.970251, 4.970322, 4.971179, 4.973058, 
    4.975195, 4.977999, 4.978202, 4.978607, 4.979215, 4.980005, 4.980972, 
    4.982105, 4.983404, 4.984862, 4.986478, 4.988243, 4.990149, 4.992177, 
    4.994302, 4.996484, 4.998657, 5.000737, 5.002606, 5.004115, 5.005083,
  // height(28,21, 0-49)
    4.987054, 4.987665, 4.988129, 4.988471, 4.988711, 4.988868, 4.988958, 
    4.989, 4.989004, 4.988986, 4.988958, 4.988937, 4.988944, 4.989013, 
    4.989195, 0, 4.970282, 4.971366, 4.97281, 4.974231, 4.975453, 4.973234, 
    4.971309, 4.969253, 4.967992, 4.967446, 4.967751, 4.968876, 4.971061, 
    4.973518, 4.976734, 4.976965, 4.977419, 4.978096, 4.978973, 4.980039, 
    4.981282, 4.982694, 4.984271, 4.986003, 4.987885, 4.989907, 4.992052, 
    4.994292, 4.996589, 4.998882, 5.001087, 5.003087, 5.004737, 5.00586,
  // height(28,22, 0-49)
    4.987328, 4.98778, 4.988113, 4.988348, 4.988502, 4.988594, 4.988635, 
    4.98864, 4.988618, 4.988581, 4.988539, 4.988505, 4.988502, 4.988559, 
    4.988728, 0, 4.967324, 4.968526, 4.970151, 4.971785, 4.973213, 4.970802, 
    4.968777, 4.96666, 4.965425, 4.964967, 4.965406, 4.966697, 4.969078, 
    4.97174, 4.975243, 4.975431, 4.975869, 4.976557, 4.977474, 4.978605, 
    4.979939, 4.981463, 4.98317, 4.985048, 4.987089, 4.989276, 4.991593, 
    4.994008, 4.996481, 4.99895, 5.001328, 5.003502, 5.005326, 5.006629,
  // height(28,23, 0-49)
    4.987549, 4.987857, 4.98807, 4.988206, 4.988283, 4.988314, 4.98831, 
    4.988281, 4.988234, 4.988175, 4.988117, 4.988068, 4.988048, 4.988085, 
    4.988226, 0, 4.964871, 4.966145, 4.967893, 4.969668, 4.971232, 4.968641, 
    4.966502, 4.964304, 4.963049, 4.962618, 4.963121, 4.964503, 4.966997, 
    4.96978, 4.973461, 4.973578, 4.97397, 4.974645, 4.975582, 4.976766, 
    4.978186, 4.979832, 4.981688, 4.983741, 4.985978, 4.988378, 4.990917, 
    4.993559, 4.996259, 4.998947, 5.001537, 5.003915, 5.005933, 5.007423,
  // height(28,24, 0-49)
    4.98774, 4.98791, 4.988009, 4.988055, 4.98806, 4.988034, 4.987987, 
    4.987925, 4.987851, 4.987772, 4.987696, 4.987629, 4.987588, 4.987599, 
    4.987702, 0, 4.963188, 4.964485, 4.966293, 4.968147, 4.969785, 4.967083, 
    4.964877, 4.962627, 4.961349, 4.960917, 4.961437, 4.962847, 4.965379, 
    4.968204, 4.971961, 4.972018, 4.972366, 4.973018, 4.973957, 4.975173, 
    4.976654, 4.97839, 4.980366, 4.982566, 4.984974, 4.987565, 4.990309, 
    4.993167, 4.996087, 4.998994, 5.001799, 5.004381, 5.006594, 5.00827,
  // height(28,25, 0-49)
    4.987918, 4.987956, 4.987947, 4.987906, 4.98784, 4.98776, 4.987669, 
    4.987572, 4.98747, 4.98737, 4.987273, 4.987188, 4.987124, 4.987105, 
    4.987164, 0, 4.961998, 4.963271, 4.96508, 4.966942, 4.96859, 4.965873, 
    4.963664, 4.961417, 4.960142, 4.95971, 4.960229, 4.96163, 4.964145, 
    4.966951, 4.9707, 4.97073, 4.971062, 4.971709, 4.972658, 4.973903, 
    4.975436, 4.977246, 4.979321, 4.981645, 4.984196, 4.986951, 4.989874, 
    4.992926, 4.996044, 4.999156, 5.002161, 5.00494, 5.007341, 5.009192,
  // height(28,26, 0-49)
    4.988102, 4.988014, 4.9879, 4.98777, 4.987633, 4.987494, 4.987355, 
    4.987218, 4.987085, 4.986959, 4.98684, 4.986735, 4.98665, 4.986601, 
    4.986614, 0, 4.96127, 4.962483, 4.964233, 4.96604, 4.967638, 4.965005, 
    4.962867, 4.960688, 4.95945, 4.959028, 4.95953, 4.960891, 4.963342, 
    4.966077, 4.969729, 4.969779, 4.970129, 4.970798, 4.971775, 4.973054, 
    4.974634, 4.976504, 4.978654, 4.98107, 4.983733, 4.986615, 4.989684, 
    4.992893, 4.996181, 4.99947, 5.002655, 5.005613, 5.008188, 5.010205,
  // height(28,27, 0-49)
    4.988311, 4.988101, 4.987882, 4.987662, 4.987448, 4.987243, 4.987047, 
    4.986861, 4.986687, 4.986527, 4.986381, 4.986256, 4.986153, 4.986082, 
    4.986058, 0, 4.961052, 4.962173, 4.963817, 4.96551, 4.967003, 4.964544, 
    4.962538, 4.960472, 4.959287, 4.958868, 4.959324, 4.960605, 4.962934, 
    4.965534, 4.969001, 4.969101, 4.969494, 4.970201, 4.971213, 4.972528, 
    4.974146, 4.97606, 4.978265, 4.980749, 4.983495, 4.986478, 4.989666, 
    4.993008, 4.996446, 4.999894, 5.003249, 5.006377, 5.009121, 5.011301,
  // height(28,28, 0-49)
    4.988558, 4.98823, 4.987906, 4.987594, 4.987296, 4.987011, 4.986745, 
    4.986495, 4.986266, 4.986061, 4.985881, 4.985734, 4.98562, 4.985543, 
    4.985505, 0, 4.961629, 4.962648, 4.964153, 4.965688, 4.967029, 4.964806, 
    4.962961, 4.961018, 4.959865, 4.959403, 4.959753, 4.960879, 4.963003, 
    4.965382, 4.968564, 4.968718, 4.969153, 4.969889, 4.97092, 4.97225, 
    4.973881, 4.975813, 4.978045, 4.980568, 4.983372, 4.986431, 4.989717, 
    4.993181, 4.996759, 5.000366, 5.003891, 5.007196, 5.010116, 5.012463,
  // height(28,29, 0-49)
    4.988853, 4.988415, 4.987991, 4.98758, 4.987185, 4.986807, 4.986447, 
    4.986111, 4.985805, 4.985536, 4.985315, 4.985149, 4.985041, 4.984988, 
    4.984979, 0, 4.96272, 4.963651, 4.965005, 4.966348, 4.967486, 4.965503, 
    4.96379, 4.961924, 4.960732, 4.960146, 4.960302, 4.961183, 4.963007, 
    4.965075, 4.967861, 4.968034, 4.96848, 4.969221, 4.970254, 4.97159, 
    4.973233, 4.975191, 4.977465, 4.980054, 4.982945, 4.986122, 4.989549, 
    4.993178, 4.996941, 5.000747, 5.004481, 5.007996, 5.01112, 5.013654,
  // height(28,30, 0-49)
    4.98853, 4.987349, 4.986206, 4.985108, 4.984058, 4.983053, 4.98209, 
    4.981159, 4.980254, 4.979371, 4.978508, 4.977676, 4.976903, 4.976246, 
    4.975795, 4.974938, 4.965952, 4.966966, 4.968203, 4.969349, 4.970299, 
    4.968656, 4.967254, 4.965686, 4.964678, 4.964137, 4.964175, 4.964772, 
    4.966136, 4.967617, 4.969641, 4.969453, 4.969526, 4.969896, 4.970581, 
    4.971605, 4.972989, 4.974744, 4.976882, 4.979402, 4.982292, 4.98553, 
    4.989075, 4.992872, 4.996842, 5.000887, 5.004877, 5.008653, 5.012033, 
    5.014809,
  // height(28,31, 0-49)
    4.988934, 4.987695, 4.986489, 4.98532, 4.98419, 4.983098, 4.982041, 
    4.981017, 4.980021, 4.979056, 4.978122, 4.977229, 4.976397, 4.975665, 
    4.975098, 4.974432, 4.965597, 4.966311, 4.967228, 4.96806, 4.968717, 
    4.96726, 4.965956, 4.96447, 4.963483, 4.962937, 4.96296, 4.963528, 
    4.964809, 4.96617, 4.967934, 4.96792, 4.968172, 4.968722, 4.969593, 
    4.970803, 4.972375, 4.97432, 4.976649, 4.979359, 4.982438, 4.985861, 
    4.989586, 4.993555, 4.997685, 5.001874, 5.005987, 5.009863, 5.013318, 
    5.016133,
  // height(28,32, 0-49)
    4.989329, 4.988023, 4.986743, 4.985494, 4.984277, 4.983092, 4.98194, 
    4.980819, 4.979729, 4.978675, 4.977658, 4.976685, 4.97577, 4.974939, 
    4.974227, 4.97373, 4.965408, 4.965789, 4.966353, 4.966842, 4.96719, 
    4.965924, 4.964731, 4.963346, 4.9624, 4.961866, 4.961875, 4.962408, 
    4.963588, 4.964805, 4.966289, 4.966444, 4.96687, 4.967595, 4.96864, 
    4.970027, 4.971777, 4.973903, 4.976413, 4.979305, 4.982565, 4.986166, 
    4.990065, 4.994201, 4.998487, 5.002816, 5.007049, 5.011023, 5.014543, 
    5.017394,
  // height(28,33, 0-49)
    4.989703, 4.988327, 4.986968, 4.985633, 4.984324, 4.983045, 4.981792, 
    4.980573, 4.979386, 4.978236, 4.977127, 4.976064, 4.975055, 4.974112, 
    4.973249, 4.97283, 4.965299, 4.96534, 4.965545, 4.96569, 4.965733, 
    4.964666, 4.963603, 4.962349, 4.961465, 4.960958, 4.96096, 4.961446, 
    4.962501, 4.963549, 4.96474, 4.96506, 4.965649, 4.966537, 4.967746, 
    4.969299, 4.971216, 4.973511, 4.976191, 4.979255, 4.982684, 4.986455, 
    4.990518, 4.994809, 4.99924, 5.003698, 5.008042, 5.0121, 5.015676, 
    5.018547,
  // height(28,34, 0-49)
    4.990031, 4.988589, 4.987155, 4.985735, 4.984336, 4.982958, 4.981607, 
    4.980285, 4.978996, 4.977746, 4.976541, 4.975382, 4.974274, 4.973217, 
    4.972211, 4.971758, 4.965207, 4.964923, 4.964778, 4.964593, 4.964345, 
    4.963485, 4.962573, 4.961481, 4.960687, 4.960222, 4.960217, 4.960645, 
    4.961547, 4.962411, 4.963303, 4.963782, 4.964528, 4.965569, 4.966932, 
    4.96864, 4.970713, 4.973166, 4.976003, 4.979225, 4.982812, 4.986735, 
    4.990946, 4.995378, 4.999937, 5.004506, 5.008938, 5.013061, 5.01667, 
    5.019539,
  // height(28,35, 0-49)
    4.990283, 4.988789, 4.987288, 4.985792, 4.984304, 4.982832, 4.981381, 
    4.979957, 4.978567, 4.977216, 4.97591, 4.974653, 4.973446, 4.97228, 
    4.971144, 4.970554, 4.965104, 4.964519, 4.964046, 4.963553, 4.96304, 
    4.962392, 4.96165, 4.960749, 4.960071, 4.959666, 4.959654, 4.960008, 
    4.960733, 4.961397, 4.961999, 4.96263, 4.963524, 4.964712, 4.966218, 
    4.96807, 4.970286, 4.972882, 4.975864, 4.979228, 4.982954, 4.987012, 
    4.991352, 4.995899, 5.000561, 5.005215, 5.009709, 5.013865, 5.017476, 
    5.020309,
  // height(28,36, 0-49)
    4.990426, 4.988896, 4.987345, 4.985782, 4.984218, 4.982658, 4.981112, 
    4.97959, 4.9781, 4.976649, 4.975245, 4.973891, 4.972588, 4.971323, 
    4.970076, 4.969267, 4.964972, 4.964121, 4.963349, 4.962579, 4.961828, 
    4.961393, 4.960837, 4.960156, 4.959619, 4.959288, 4.959268, 4.959536, 
    4.960064, 4.96052, 4.960848, 4.961624, 4.962659, 4.963984, 4.965623, 
    4.967606, 4.969953, 4.972678, 4.975785, 4.979272, 4.983116, 4.987284, 
    4.991723, 4.996358, 5.001091, 5.005792, 5.010311, 5.014461, 5.01803, 
    5.020787,
  // height(28,37, 0-49)
    4.99042, 4.988878, 4.987295, 4.985683, 4.984055, 4.98242, 4.980792, 
    4.97918, 4.977595, 4.97605, 4.974551, 4.973106, 4.971712, 4.970358, 
    4.969019, 4.967945, 4.964811, 4.963729, 4.962691, 4.961675, 4.960719, 
    4.960494, 4.960138, 4.959701, 4.959327, 4.959084, 4.959058, 4.959228, 
    4.959541, 4.959791, 4.959871, 4.960784, 4.961951, 4.963401, 4.965164, 
    4.967265, 4.969728, 4.972565, 4.975777, 4.979362, 4.983298, 4.987546, 
    4.992053, 4.996737, 5.001498, 5.006205, 5.0107, 5.014793, 5.018272, 5.0209,
  // height(28,38, 0-49)
    4.99023, 4.988701, 4.987109, 4.98547, 4.983797, 4.982105, 4.980407, 
    4.978717, 4.977051, 4.97542, 4.973835, 4.972305, 4.97083, 4.969398, 
    4.967984, 4.966624, 4.964621, 4.963344, 4.962071, 4.960845, 4.959713, 
    4.959695, 4.959548, 4.959376, 4.959183, 4.959043, 4.959011, 4.959078, 
    4.959167, 4.959216, 4.959079, 4.960124, 4.961415, 4.962979, 4.964853, 
    4.967059, 4.969621, 4.972549, 4.975846, 4.979504, 4.983499, 4.98779, 
    4.992322, 4.997014, 5.001755, 5.006413, 5.010828, 5.014806, 5.018132, 
    5.020571,
  // height(28,39, 0-49)
    4.98982, 4.988333, 4.986758, 4.985115, 4.983422, 4.981692, 4.979945, 
    4.978195, 4.976461, 4.974759, 4.973101, 4.971496, 4.969948, 4.968448, 
    4.966973, 4.965341, 4.964407, 4.962965, 4.961492, 4.960084, 4.958814, 
    4.958994, 4.959059, 4.959167, 4.959174, 4.959148, 4.959116, 4.959077, 
    4.958942, 4.958804, 4.958484, 4.959653, 4.96106, 4.962731, 4.964701, 
    4.966998, 4.96964, 4.972637, 4.975991, 4.979691, 4.983709, 4.988005, 
    4.992517, 4.997162, 5.001826, 5.006374, 5.010642, 5.014437, 5.017542, 
    5.019726,
  // height(28,40, 0-49)
    4.989163, 4.987743, 4.986215, 4.984596, 4.982908, 4.981167, 4.979392, 
    4.977604, 4.975822, 4.974064, 4.972347, 4.970681, 4.969072, 4.967516, 
    4.965992, 4.964116, 4.964172, 4.962595, 4.960951, 4.959398, 4.958017, 
    4.958385, 4.958663, 4.959061, 4.959281, 4.959382, 4.959355, 4.959212, 
    4.958863, 4.958557, 4.95809, 4.959379, 4.960891, 4.962658, 4.964714, 
    4.967083, 4.969785, 4.972829, 4.97621, 4.979917, 4.983921, 4.988175, 
    4.992615, 4.997153, 5.001677, 5.006044, 5.010092, 5.013627, 5.016435, 
    5.018291,
  // height(28,41, 0-49)
    4.988236, 4.986912, 4.985459, 4.983894, 4.982239, 4.980513, 4.978737, 
    4.976935, 4.975128, 4.973335, 4.971576, 4.969865, 4.968209, 4.966607, 
    4.965042, 4.962963, 4.963916, 4.962226, 4.960443, 4.958775, 4.957313, 
    4.957856, 4.958346, 4.959037, 4.959479, 4.959718, 4.959705, 4.959471, 
    4.958921, 4.958473, 4.957899, 4.959299, 4.96091, 4.962762, 4.96489, 
    4.967316, 4.970056, 4.973118, 4.976497, 4.980174, 4.984117, 4.988278, 
    4.992589, 4.996957, 5.001267, 5.005378, 5.009124, 5.012317, 5.014746, 
    5.016197,
  // height(28,42, 0-49)
    4.98703, 4.98583, 4.984478, 4.982997, 4.981404, 4.979722, 4.977974, 
    4.976183, 4.974374, 4.97257, 4.97079, 4.96905, 4.96736, 4.965723, 
    4.964126, 4.961891, 4.963639, 4.961859, 4.95996, 4.958206, 4.956691, 
    4.957398, 4.958096, 4.959077, 4.959745, 4.96013, 4.960144, 4.959831, 
    4.959105, 4.958547, 4.957901, 4.959409, 4.961112, 4.963038, 4.965222, 
    4.967688, 4.970444, 4.973498, 4.976838, 4.980443, 4.98428, 4.988293, 
    4.992411, 4.996538, 5.000558, 5.00433, 5.007689, 5.010449, 5.012415, 
    5.013385,
  // height(28,43, 0-49)
    4.98554, 4.984489, 4.983268, 4.981898, 4.980398, 4.978789, 4.977099, 
    4.975349, 4.973565, 4.971771, 4.96999, 4.96824, 4.96653, 4.964868, 
    4.963245, 4.9609, 4.963339, 4.961486, 4.959499, 4.957683, 4.956139, 
    4.956997, 4.957892, 4.959154, 4.960049, 4.960588, 4.96064, 4.960272, 
    4.959402, 4.958764, 4.958083, 4.959694, 4.961483, 4.963474, 4.965702, 
    4.968185, 4.970934, 4.973947, 4.977213, 4.980706, 4.984384, 4.988188, 
    4.992046, 4.99586, 4.999508, 5.002852, 5.005733, 5.007973, 5.009391, 
    5.009803,
  // height(28,44, 0-49)
    4.983782, 4.982901, 4.981836, 4.980603, 4.979224, 4.977719, 4.976113, 
    4.974431, 4.972697, 4.970939, 4.969179, 4.967435, 4.965723, 4.964047, 
    4.962406, 4.959991, 4.963014, 4.961103, 4.959048, 4.957194, 4.955643, 
    4.956639, 4.95772, 4.959247, 4.960364, 4.961061, 4.961168, 4.960768, 
    4.95979, 4.959107, 4.958425, 4.960135, 4.962002, 4.964049, 4.966306, 
    4.968788, 4.971504, 4.974445, 4.977598, 4.980931, 4.984395, 4.987931, 
    4.991458, 4.994877, 4.99807, 5.000897, 5.003209, 5.00484, 5.005627, 
    5.005414,
  // height(28,45, 0-49)
    4.981774, 4.981083, 4.980196, 4.979126, 4.977894, 4.97652, 4.975028, 
    4.973438, 4.971782, 4.970082, 4.968363, 4.966645, 4.964943, 4.963265, 
    4.961613, 4.959162, 4.962658, 4.960703, 4.958603, 4.956729, 4.955187, 
    4.956307, 4.957557, 4.959331, 4.960659, 4.961514, 4.961693, 4.961289, 
    4.960246, 4.959553, 4.958898, 4.960707, 4.962646, 4.964738, 4.967009, 
    4.969471, 4.972126, 4.974962, 4.977961, 4.981081, 4.984278, 4.987478, 
    4.990602, 4.993547, 4.996198, 4.998419, 5.000072, 5.001008, 5.001089, 
    5.000189,
  // height(28,46, 0-49)
    4.979548, 4.979063, 4.978371, 4.977488, 4.976427, 4.975208, 4.973854, 
    4.972385, 4.970828, 4.969208, 4.96755, 4.965873, 4.964198, 4.96253, 
    4.960874, 4.958412, 4.962271, 4.960286, 4.958158, 4.95628, 4.95476, 
    4.955986, 4.957387, 4.959378, 4.960902, 4.961915, 4.96218, 4.961805, 
    4.96074, 4.960072, 4.959472, 4.961374, 4.96338, 4.965507, 4.967777, 
    4.970197, 4.972763, 4.975461, 4.978261, 4.981122, 4.983987, 4.986786, 
    4.989431, 4.991823, 4.993845, 4.995374, 4.996282, 4.996446, 4.995755, 
    4.994122,
  // height(28,47, 0-49)
    4.977147, 4.976876, 4.976397, 4.975716, 4.974848, 4.973806, 4.972611, 
    4.971286, 4.96985, 4.968332, 4.966752, 4.965134, 4.963496, 4.961848, 
    4.960196, 4.957739, 4.96185, 4.959847, 4.957707, 4.955839, 4.95435, 
    4.955663, 4.957192, 4.959366, 4.961065, 4.962229, 4.962596, 4.962281, 
    4.96124, 4.96063, 4.960107, 4.962099, 4.964166, 4.966316, 4.96857, 
    4.970924, 4.973373, 4.975894, 4.978453, 4.981, 4.983474, 4.985802, 
    4.987894, 4.98965, 4.990963, 4.991716, 4.991806, 4.991132, 4.989618, 
    4.987222,
  // height(28,48, 0-49)
    4.974618, 4.974567, 4.974308, 4.973845, 4.973186, 4.972341, 4.971326, 
    4.970162, 4.968867, 4.967466, 4.965981, 4.964435, 4.962846, 4.961228, 
    4.959587, 4.957145, 4.961398, 4.959391, 4.957252, 4.9554, 4.953947, 
    4.955328, 4.956959, 4.959277, 4.961123, 4.962427, 4.962908, 4.962682, 
    4.96171, 4.961189, 4.960761, 4.962839, 4.964956, 4.967119, 4.969338, 
    4.971605, 4.973905, 4.976213, 4.978484, 4.980662, 4.982685, 4.984473, 
    4.98594, 4.986984, 4.987511, 4.987416, 4.986622, 4.985056, 4.982687, 
    4.979521,
  // height(28,49, 0-49)
    4.971751, 4.97187, 4.971794, 4.971513, 4.971032, 4.970352, 4.969482, 
    4.968434, 4.96722, 4.965861, 4.964369, 4.962768, 4.961073, 4.959293, 
    4.957433, 4.953966, 4.963982, 4.960976, 4.957507, 4.954463, 4.952083, 
    4.955269, 4.95878, 4.963472, 4.966963, 4.969119, 4.969381, 4.967987, 
    4.964842, 4.962405, 4.959975, 4.962437, 4.964849, 4.967206, 4.969516, 
    4.971771, 4.973949, 4.976017, 4.977924, 4.979613, 4.981015, 4.982051, 
    4.98264, 4.982693, 4.982131, 4.980882, 4.978908, 4.976194, 4.972773, 
    4.968725,
  // height(29,0, 0-49)
    4.971556, 4.973361, 4.974815, 4.975937, 4.976742, 4.97725, 4.977488, 
    4.977488, 4.977288, 4.976929, 4.976456, 4.97591, 4.975338, 4.97478, 
    4.974274, 4.973676, 4.973505, 4.973238, 4.973083, 4.97306, 4.973165, 
    4.973533, 4.973971, 4.974497, 4.975105, 4.975779, 4.976512, 4.977307, 
    4.978165, 4.979098, 4.980094, 4.981372, 4.982794, 4.984384, 4.986169, 
    4.988163, 4.99037, 4.992781, 4.995366, 4.998078, 5.000845, 5.003565, 
    5.00611, 5.008316, 5.009995, 5.010931, 5.010883, 5.009605, 5.006854, 
    5.002412,
  // height(29,1, 0-49)
    4.97285, 4.9746, 4.976003, 4.977079, 4.977844, 4.97832, 4.978535, 
    4.978521, 4.978314, 4.977955, 4.977486, 4.976948, 4.976385, 4.975832, 
    4.975327, 4.974553, 4.974493, 4.974136, 4.97386, 4.973703, 4.973669, 
    4.97404, 4.974442, 4.974925, 4.975485, 4.976109, 4.976785, 4.977513, 
    4.978296, 4.979141, 4.980009, 4.981315, 4.982766, 4.984389, 4.986212, 
    4.988253, 4.990514, 4.992992, 4.995659, 4.998469, 5.001352, 5.00421, 
    5.006918, 5.009318, 5.011222, 5.012416, 5.012663, 5.011715, 5.009322, 
    5.005255,
  // height(29,2, 0-49)
    4.974152, 4.975846, 4.977199, 4.978231, 4.97896, 4.979407, 4.979604, 
    4.979578, 4.979369, 4.979012, 4.978549, 4.978021, 4.977464, 4.976915, 
    4.976405, 4.97546, 4.975474, 4.975027, 4.974627, 4.974336, 4.974163, 
    4.974525, 4.97488, 4.975307, 4.975816, 4.976388, 4.977014, 4.977693, 
    4.978423, 4.979195, 4.979949, 4.981287, 4.982766, 4.984417, 4.986269, 
    4.988337, 4.990631, 4.993144, 4.995852, 4.998711, 5.001653, 5.004588, 
    5.007389, 5.009909, 5.011964, 5.013349, 5.013828, 5.013155, 5.011086, 
    5.007389,
  // height(29,3, 0-49)
    4.975455, 4.977093, 4.978398, 4.979385, 4.98008, 4.980501, 4.980679, 
    4.980646, 4.980434, 4.980083, 4.979627, 4.979106, 4.978555, 4.978006, 
    4.977489, 4.976379, 4.976416, 4.975876, 4.975358, 4.974937, 4.97463, 
    4.974973, 4.975272, 4.975631, 4.976077, 4.976596, 4.977183, 4.977833, 
    4.978536, 4.979261, 4.979921, 4.981289, 4.982796, 4.98447, 4.98634, 
    4.988424, 4.990729, 4.993248, 4.995963, 4.998829, 5.001781, 5.004733, 
    5.007569, 5.010144, 5.012286, 5.013795, 5.014449, 5.014008, 5.01223, 
    5.008885,
  // height(29,4, 0-49)
    4.976765, 4.978344, 4.979596, 4.980538, 4.981195, 4.981589, 4.981749, 
    4.981706, 4.981493, 4.981143, 4.980695, 4.980181, 4.979634, 4.979084, 
    4.978553, 4.977294, 4.977292, 4.976662, 4.976037, 4.975495, 4.975061, 
    4.975371, 4.975604, 4.975881, 4.976256, 4.976723, 4.97728, 4.97792, 
    4.978625, 4.979328, 4.979919, 4.98132, 4.982853, 4.984545, 4.986426, 
    4.988512, 4.990811, 4.993315, 4.996003, 4.99884, 5.00176, 5.004683, 
    5.0075, 5.010075, 5.012246, 5.013824, 5.0146, 5.014348, 5.012831, 5.009826,
  // height(29,5, 0-49)
    4.978075, 4.97959, 4.980784, 4.981678, 4.982295, 4.98266, 4.9828, 
    4.982745, 4.982529, 4.982182, 4.981737, 4.981228, 4.980682, 4.980126, 
    4.979578, 4.978192, 4.978077, 4.977365, 4.976644, 4.975996, 4.975449, 
    4.975712, 4.975867, 4.976048, 4.976345, 4.976757, 4.977293, 4.977944, 
    4.978681, 4.97939, 4.979939, 4.981371, 4.982926, 4.984634, 4.986518, 
    4.988595, 4.990872, 4.99334, 4.995981, 4.998755, 5.001609, 5.004463, 
    5.007217, 5.009746, 5.0119, 5.013502, 5.014358, 5.014255, 5.012973, 
    5.010293,
  // height(29,6, 0-49)
    4.979375, 4.980821, 4.981953, 4.982794, 4.983367, 4.983699, 4.983816, 
    4.983747, 4.983525, 4.983177, 4.982736, 4.982229, 4.981682, 4.981119, 
    4.980551, 4.979065, 4.978755, 4.977969, 4.97717, 4.976434, 4.975792, 
    4.975995, 4.976058, 4.976129, 4.976338, 4.976693, 4.977218, 4.977898, 
    4.978695, 4.979438, 4.979978, 4.981435, 4.98301, 4.984728, 4.986608, 
    4.988667, 4.990908, 4.993323, 4.995894, 4.998584, 5.00134, 5.004094, 
    5.006751, 5.009197, 5.011295, 5.012885, 5.013788, 5.013808, 5.012739, 
    5.010373,
  // height(29,7, 0-49)
    4.980656, 4.982026, 4.983089, 4.983871, 4.984396, 4.98469, 4.984782, 
    4.984697, 4.984466, 4.984116, 4.983675, 4.98317, 4.982621, 4.982047, 
    4.981458, 4.979904, 4.979315, 4.978468, 4.977612, 4.976809, 4.976092, 
    4.976218, 4.97618, 4.976123, 4.976236, 4.976532, 4.977053, 4.977777, 
    4.978659, 4.979466, 4.980029, 4.981503, 4.983092, 4.984814, 4.986686, 
    4.988718, 4.99091, 4.993259, 4.995742, 4.998327, 5.000965, 5.003592, 
    5.006126, 5.008463, 5.010478, 5.012031, 5.012955, 5.013077, 5.012204, 
    5.010143,
  // height(29,8, 0-49)
    4.981897, 4.983184, 4.984174, 4.984893, 4.985365, 4.98562, 4.985681, 
    4.985578, 4.985337, 4.984982, 4.984541, 4.984036, 4.983485, 4.982903, 
    4.982292, 4.980708, 4.979747, 4.978858, 4.977969, 4.977125, 4.976357, 
    4.976388, 4.976235, 4.976039, 4.976047, 4.976282, 4.976804, 4.977584, 
    4.978576, 4.979469, 4.980087, 4.981573, 4.983167, 4.984883, 4.986736, 
    4.988731, 4.990869, 4.993138, 4.99552, 4.997984, 5.000488, 5.002973, 
    5.005363, 5.007573, 5.009488, 5.010984, 5.011919, 5.012128, 5.011442, 
    5.009677,
  // height(29,9, 0-49)
    4.983086, 4.984283, 4.985192, 4.985842, 4.986258, 4.986469, 4.986499, 
    4.986375, 4.986122, 4.985764, 4.985322, 4.984818, 4.984266, 4.983675, 
    4.983043, 4.981473, 4.980051, 4.97914, 4.978247, 4.977389, 4.976596, 
    4.976516, 4.976236, 4.97589, 4.975786, 4.975957, 4.976483, 4.977327, 
    4.978443, 4.979445, 4.980153, 4.981635, 4.983224, 4.984926, 4.986752, 
    4.988701, 4.990771, 4.992952, 4.995222, 4.997556, 4.999913, 5.002243, 
    5.004482, 5.006552, 5.008358, 5.009792, 5.010726, 5.011018, 5.010513, 
    5.009043,
  // height(29,10, 0-49)
    4.984201, 4.9853, 4.986125, 4.986701, 4.987059, 4.987222, 4.987219, 
    4.987072, 4.986808, 4.986445, 4.986005, 4.985502, 4.984953, 4.984358, 
    4.983712, 4.982196, 4.980223, 4.979319, 4.978451, 4.977612, 4.976825, 
    4.976614, 4.976199, 4.975692, 4.975474, 4.975579, 4.976107, 4.977016, 
    4.978267, 4.979397, 4.980227, 4.981689, 4.983257, 4.984932, 4.986719, 
    4.988612, 4.990606, 4.992688, 4.99484, 4.997035, 4.99924, 5.001411, 
    5.003496, 5.005424, 5.007121, 5.008492, 5.009428, 5.009802, 5.009476, 
    5.008297,
  // height(29,11, 0-49)
    4.985221, 4.986217, 4.986951, 4.987451, 4.987747, 4.987863, 4.987825, 
    4.987659, 4.987381, 4.987016, 4.986578, 4.986081, 4.985535, 4.984943, 
    4.984293, 4.982874, 4.980265, 4.979398, 4.978592, 4.977806, 4.977054, 
    4.9767, 4.976141, 4.975471, 4.975133, 4.975172, 4.9757, 4.976673, 
    4.978061, 4.979329, 4.980305, 4.981731, 4.983263, 4.984897, 4.98663, 
    4.988455, 4.990363, 4.992339, 4.994365, 4.996418, 4.998469, 5.000483, 
    5.002415, 5.004209, 5.005803, 5.007117, 5.008061, 5.008524, 5.008382, 
    5.00749,
  // height(29,12, 0-49)
    4.986129, 4.987016, 4.987657, 4.988077, 4.98831, 4.988379, 4.988306, 
    4.988117, 4.987829, 4.987461, 4.98703, 4.986541, 4.986005, 4.985423, 
    4.984781, 4.983505, 4.980176, 4.979388, 4.978679, 4.977983, 4.977303, 
    4.976789, 4.976083, 4.975247, 4.974793, 4.974764, 4.975285, 4.976314, 
    4.977836, 4.979246, 4.980394, 4.981762, 4.983236, 4.98481, 4.986475, 
    4.98822, 4.99003, 4.991893, 4.99379, 4.9957, 4.997602, 4.999462, 5.00125, 
    5.002921, 5.004425, 5.005697, 5.00666, 5.007222, 5.007267, 5.006666,
  // height(29,13, 0-49)
    4.98691, 4.987683, 4.988225, 4.988565, 4.988734, 4.988751, 4.988646, 
    4.988435, 4.988138, 4.98777, 4.987345, 4.98687, 4.986352, 4.985789, 
    4.985172, 4.984077, 4.97996, 4.979289, 4.978722, 4.978153, 4.97758, 
    4.976897, 4.976046, 4.975048, 4.974481, 4.974383, 4.974892, 4.975965, 
    4.977607, 4.979157, 4.980497, 4.98178, 4.983175, 4.984669, 4.986247, 
    4.987896, 4.989599, 4.991342, 4.993107, 4.994876, 4.996633, 4.998353, 
    5.000012, 5.001576, 5.003008, 5.004256, 5.005257, 5.005929, 5.00617, 
    5.005861,
  // height(29,14, 0-49)
    4.987552, 4.988207, 4.988649, 4.988905, 4.989006, 4.988974, 4.988832, 
    4.988601, 4.988295, 4.987929, 4.987513, 4.987056, 4.986562, 4.986031, 
    4.985457, 4.984582, 4.97962, 4.979108, 4.978724, 4.978326, 4.977896, 
    4.977039, 4.976047, 4.974896, 4.974222, 4.974059, 4.974547, 4.975648, 
    4.977391, 4.979072, 4.980613, 4.981785, 4.983075, 4.984465, 4.985938, 
    4.987476, 4.989061, 4.990677, 4.992309, 4.993942, 4.995565, 4.997159, 
    4.998707, 5.000188, 5.001571, 5.002817, 5.003875, 5.004673, 5.00512, 
    5.005102,
  // height(29,15, 0-49)
    4.988047, 4.988579, 4.988916, 4.989087, 4.989118, 4.989033, 4.988854, 
    4.988601, 4.988286, 4.987922, 4.98752, 4.987084, 4.986623, 4.986136, 
    4.985628, 4.985004, 4.979161, 4.978853, 4.978694, 4.978505, 4.978258, 
    4.977225, 4.976098, 4.97481, 4.974041, 4.973814, 4.974275, 4.975384, 
    4.977204, 4.978997, 4.980742, 4.981776, 4.982933, 4.984197, 4.985542, 
    4.986952, 4.988406, 4.989891, 4.991391, 4.992896, 4.994396, 4.995882, 
    4.997343, 4.998764, 5.000125, 5.001397, 5.002533, 5.003475, 5.004138, 
    5.004411,
  // height(29,16, 0-49)
    4.988392, 4.988796, 4.989022, 4.989101, 4.98906, 4.98892, 4.988703, 
    4.988425, 4.988101, 4.987741, 4.987353, 4.986944, 4.986523, 4.986093, 
    4.985668, 4.985326, 4.978594, 4.978531, 4.978637, 4.978697, 4.978667, 
    4.977459, 4.976213, 4.974801, 4.973953, 4.973667, 4.974092, 4.975191, 
    4.977059, 4.978941, 4.980883, 4.98175, 4.982749, 4.983858, 4.985055, 
    4.986319, 4.987631, 4.988978, 4.990348, 4.991733, 4.993127, 4.994525, 
    4.995924, 4.997314, 4.998682, 5.000005, 5.001247, 5.002351, 5.00324, 
    5.003806,
  // height(29,17, 0-49)
    4.988588, 4.988854, 4.988962, 4.988945, 4.988825, 4.988625, 4.988366, 
    4.988063, 4.987727, 4.98737, 4.986999, 4.986622, 4.986247, 4.985889, 
    4.985566, 4.98553, 4.977942, 4.97816, 4.978563, 4.978907, 4.979125, 
    4.977752, 4.9764, 4.974884, 4.973968, 4.973629, 4.97401, 4.97508, 
    4.976967, 4.978909, 4.981034, 4.981708, 4.982517, 4.983448, 4.984474, 
    4.985574, 4.986732, 4.987938, 4.98918, 4.990454, 4.991757, 4.99309, 
    4.994452, 4.995841, 4.997247, 4.998652, 5.000022, 5.001309, 5.002435, 
    5.003295,
  // height(29,18, 0-49)
    4.988639, 4.988755, 4.988736, 4.98861, 4.988406, 4.988142, 4.987838, 
    4.987507, 4.987159, 4.986805, 4.986453, 4.986112, 4.985792, 4.985513, 
    4.98531, 4.985602, 4.977243, 4.977769, 4.978495, 4.979146, 4.979639, 
    4.978107, 4.976663, 4.97506, 4.974088, 4.973702, 4.974034, 4.975058, 
    4.976934, 4.978906, 4.981187, 4.981641, 4.982238, 4.982964, 4.983794, 
    4.984714, 4.985708, 4.986764, 4.987881, 4.989054, 4.990283, 4.991574, 
    4.992928, 4.994346, 4.995821, 4.997337, 4.998865, 5.000354, 5.001728, 
    5.002884,
  // height(29,19, 0-49)
    4.98855, 4.988499, 4.988338, 4.988094, 4.987796, 4.987462, 4.987109, 
    4.986747, 4.986388, 4.986039, 4.985707, 4.985406, 4.985149, 4.984963, 
    4.984892, 4.98553, 4.976555, 4.977411, 4.978475, 4.979445, 4.980222, 
    4.978542, 4.977019, 4.975341, 4.974323, 4.973892, 4.974168, 4.975128, 
    4.976965, 4.978934, 4.981341, 4.981552, 4.981909, 4.982407, 4.983021, 
    4.98374, 4.984555, 4.985459, 4.98645, 4.98753, 4.988702, 4.989972, 
    4.991343, 4.99282, 4.994395, 4.996053, 4.997765, 4.999477, 5.001114, 
    5.002572,
  // height(29,20, 0-49)
    4.989048, 4.989503, 4.989847, 4.990098, 4.99027, 4.990378, 4.990433, 
    4.990442, 4.990415, 4.99036, 4.990286, 4.990209, 4.990146, 4.990134, 
    4.990227, 0, 4.975359, 4.976153, 4.977207, 4.978203, 4.979018, 4.976952, 
    4.975087, 4.973069, 4.971763, 4.971109, 4.97125, 4.972173, 4.974099, 
    4.976275, 4.979077, 4.979346, 4.979769, 4.980332, 4.98101, 4.981788, 
    4.982655, 4.983606, 4.984644, 4.985774, 4.987006, 4.988348, 4.98981, 
    4.991399, 4.993111, 4.994935, 4.996837, 4.99877, 5.000656, 5.002386,
  // height(29,21, 0-49)
    4.988827, 4.98916, 4.989402, 4.98957, 4.989676, 4.989734, 4.989754, 
    4.989744, 4.989711, 4.98966, 4.9896, 4.989542, 4.989507, 4.989525, 
    4.989647, 0, 4.972302, 4.973264, 4.974558, 4.975825, 4.976907, 4.974704, 
    4.972797, 4.970784, 4.969567, 4.96906, 4.969389, 4.970522, 4.972679, 
    4.975086, 4.978195, 4.978409, 4.978792, 4.979332, 4.980003, 4.980789, 
    4.981676, 4.98266, 4.983741, 4.984922, 4.986211, 4.987618, 4.989153, 
    4.990819, 4.992617, 4.994532, 4.996534, 4.998575, 5.000577, 5.002439,
  // height(29,22, 0-49)
    4.988561, 4.988786, 4.988936, 4.989029, 4.989077, 4.989089, 4.989075, 
    4.989043, 4.988997, 4.988944, 4.988889, 4.988842, 4.988819, 4.988848, 
    4.988978, 0, 4.970036, 4.971129, 4.972622, 4.974118, 4.975419, 4.973063, 
    4.971076, 4.969011, 4.967807, 4.967357, 4.967772, 4.969004, 4.971275, 
    4.973795, 4.977079, 4.977161, 4.977431, 4.977885, 4.978497, 4.979252, 
    4.980139, 4.981151, 4.982288, 4.983549, 4.98494, 4.986465, 4.988132, 
    4.989944, 4.991897, 4.993972, 4.996139, 4.998345, 5.000515, 5.002546,
  // height(29,23, 0-49)
    4.988266, 4.988394, 4.988463, 4.988487, 4.988479, 4.988449, 4.988403, 
    4.988348, 4.988288, 4.988229, 4.988175, 4.988132, 4.988114, 4.988146, 
    4.988268, 0, 4.968285, 4.969466, 4.971102, 4.972762, 4.974215, 4.971715, 
    4.969638, 4.967495, 4.966257, 4.9658, 4.966229, 4.967482, 4.969783, 
    4.972326, 4.975673, 4.975587, 4.97571, 4.976046, 4.976573, 4.977282, 
    4.978163, 4.979208, 4.980416, 4.981785, 4.983315, 4.985008, 4.986862, 
    4.988875, 4.991038, 4.993327, 4.995707, 4.998123, 5.000495, 5.002719,
  // height(29,24, 0-49)
    4.987961, 4.987996, 4.987988, 4.98795, 4.987892, 4.987821, 4.987746, 
    4.98767, 4.987597, 4.987533, 4.987478, 4.987438, 4.987423, 4.987453, 
    4.987559, 0, 4.967278, 4.968503, 4.970228, 4.971992, 4.973543, 4.970967, 
    4.968838, 4.966646, 4.96537, 4.964878, 4.96527, 4.966482, 4.968736, 
    4.971223, 4.974539, 4.974289, 4.974264, 4.97447, 4.974896, 4.975535, 
    4.976382, 4.977432, 4.978685, 4.980134, 4.981779, 4.98362, 4.985648, 
    4.987854, 4.990224, 4.992731, 4.995331, 4.997964, 5.000548, 5.002974,
  // height(29,25, 0-49)
    4.98766, 4.987607, 4.987528, 4.98743, 4.987325, 4.987216, 4.987114, 
    4.987021, 4.986938, 4.986869, 4.986818, 4.986785, 4.986776, 4.986806, 
    4.986895, 0, 4.966704, 4.967937, 4.969695, 4.971504, 4.973098, 4.970532, 
    4.968414, 4.966226, 4.964935, 4.964411, 4.964749, 4.965886, 4.968045, 
    4.970422, 4.973626, 4.973247, 4.973096, 4.973194, 4.973528, 4.974099, 
    4.974905, 4.975947, 4.977223, 4.97873, 4.980465, 4.982426, 4.984601, 
    4.986979, 4.989538, 4.992245, 4.995053, 4.997897, 5.000687, 5.003313,
  // height(29,26, 0-49)
    4.987382, 4.987242, 4.987093, 4.986938, 4.986787, 4.986643, 4.986514, 
    4.986403, 4.986313, 4.986247, 4.986204, 4.986186, 4.986193, 4.986231, 
    4.986312, 0, 4.966497, 4.967708, 4.969454, 4.971251, 4.972836, 4.970378, 
    4.968344, 4.96622, 4.96495, 4.964405, 4.96468, 4.965718, 4.967741, 
    4.969964, 4.972982, 4.972522, 4.972288, 4.972305, 4.972567, 4.97308, 
    4.973845, 4.974867, 4.976147, 4.977685, 4.979478, 4.981522, 4.983808, 
    4.986319, 4.989032, 4.991911, 4.994902, 4.997937, 5.000921, 5.003737,
  // height(29,27, 0-49)
    4.987139, 4.986915, 4.986696, 4.986484, 4.986285, 4.986104, 4.98595, 
    4.985823, 4.985728, 4.985668, 4.985642, 4.98565, 4.985687, 4.985753, 
    4.985845, 0, 4.966663, 4.967835, 4.969529, 4.971269, 4.972798, 4.970535, 
    4.968647, 4.966635, 4.965405, 4.964836, 4.965031, 4.96594, 4.967781, 
    4.969799, 4.972559, 4.972056, 4.971772, 4.971733, 4.971939, 4.972399, 
    4.97312, 4.974112, 4.975377, 4.97692, 4.978742, 4.980838, 4.983202, 
    4.985818, 4.98866, 4.991688, 4.994846, 4.998058, 5.001228, 5.00423,
  // height(29,28, 0-49)
    4.986944, 4.986639, 4.986349, 4.986075, 4.985826, 4.985606, 4.985421, 
    4.985277, 4.985176, 4.985127, 4.985129, 4.985179, 4.985272, 4.985394, 
    4.985533, 0, 4.967456, 4.968589, 4.970207, 4.971852, 4.973289, 4.971285, 
    4.969576, 4.967695, 4.966493, 4.965866, 4.965929, 4.966646, 4.968236, 
    4.969983, 4.972405, 4.971874, 4.97155, 4.971457, 4.971603, 4.971999, 
    4.97266, 4.973596, 4.97482, 4.976341, 4.978161, 4.980283, 4.982701, 
    4.985398, 4.98835, 4.991515, 4.994833, 4.998222, 5.001579, 5.004774,
  // height(29,29, 0-49)
    4.986812, 4.986425, 4.986062, 4.985725, 4.98542, 4.985151, 4.984928, 
    4.984759, 4.984652, 4.984617, 4.984658, 4.984773, 4.984951, 4.985173, 
    4.985413, 0, 4.968573, 4.969682, 4.971219, 4.972744, 4.974048, 4.972317, 
    4.970768, 4.968982, 4.967752, 4.967, 4.966858, 4.967312, 4.968576, 
    4.969975, 4.971971, 4.971394, 4.971013, 4.970857, 4.970938, 4.971271, 
    4.971876, 4.97277, 4.97397, 4.975489, 4.977334, 4.979512, 4.982013, 
    4.984826, 4.987921, 4.991253, 4.994759, 4.998352, 5.001921, 5.005327,
  // height(29,30, 0-49)
    4.986113, 4.985028, 4.983992, 4.98301, 4.982088, 4.981229, 4.980436, 
    4.979713, 4.979061, 4.978491, 4.978013, 4.977649, 4.977439, 4.977439, 
    4.97774, 4.978108, 4.970986, 4.972597, 4.974332, 4.975877, 4.977121, 
    4.975759, 4.974507, 4.972983, 4.97189, 4.971142, 4.970854, 4.971008, 
    4.971807, 4.972627, 4.973881, 4.972935, 4.972168, 4.971625, 4.971332, 
    4.971322, 4.971624, 4.972265, 4.973269, 4.974652, 4.976425, 4.978588, 
    4.981136, 4.984048, 4.987289, 4.990808, 4.994532, 4.998365, 5.002188, 
    5.005852,
  // height(29,31, 0-49)
    4.986139, 4.985011, 4.983933, 4.982914, 4.981956, 4.981061, 4.980238, 
    4.979491, 4.978826, 4.978252, 4.977779, 4.977426, 4.97722, 4.9772, 
    4.977429, 4.977726, 4.970573, 4.971944, 4.973413, 4.974692, 4.97569, 
    4.974526, 4.973392, 4.971966, 4.970906, 4.970163, 4.969861, 4.969983, 
    4.970693, 4.971382, 4.972375, 4.971571, 4.970947, 4.970544, 4.970392, 
    4.970518, 4.970953, 4.971724, 4.972854, 4.974358, 4.976247, 4.978524, 
    4.98118, 4.984198, 4.987542, 4.991161, 4.99498, 4.998902, 5.002809, 
    5.006545,
  // height(29,32, 0-49)
    4.98621, 4.985024, 4.983895, 4.982825, 4.981821, 4.980885, 4.980024, 
    4.979245, 4.978554, 4.977959, 4.97747, 4.977098, 4.97686, 4.97678, 
    4.976899, 4.977179, 4.970335, 4.971414, 4.972563, 4.973532, 4.974247, 
    4.973269, 4.972249, 4.970926, 4.969913, 4.969187, 4.968878, 4.968968, 
    4.969584, 4.97014, 4.970872, 4.970227, 4.969762, 4.969515, 4.969513, 
    4.969784, 4.970358, 4.971261, 4.972516, 4.974138, 4.976139, 4.978522, 
    4.98128, 4.984394, 4.98783, 4.991536, 4.99544, 4.999442, 5.00342, 5.007222,
  // height(29,33, 0-49)
    4.986322, 4.985071, 4.98388, 4.982752, 4.981695, 4.980709, 4.979803, 
    4.978983, 4.978255, 4.977623, 4.977099, 4.976686, 4.976392, 4.976228, 
    4.976206, 4.976455, 4.97019, 4.970946, 4.971748, 4.972381, 4.972796, 
    4.971999, 4.971097, 4.969897, 4.968946, 4.968251, 4.967942, 4.968001, 
    4.96851, 4.968925, 4.969399, 4.968927, 4.968636, 4.968554, 4.968711, 
    4.969135, 4.969853, 4.970891, 4.972271, 4.97401, 4.976117, 4.978599, 
    4.981448, 4.984647, 4.988163, 4.991945, 4.995917, 4.999985, 5.00402, 
    5.007871,
  // height(29,34, 0-49)
    4.986467, 4.98515, 4.983893, 4.982704, 4.981585, 4.980543, 4.979585, 
    4.978714, 4.977937, 4.977258, 4.976682, 4.976209, 4.97584, 4.975573, 
    4.9754, 4.975558, 4.97007, 4.970491, 4.970932, 4.971223, 4.971337, 
    4.970714, 4.969939, 4.968884, 4.968016, 4.967366, 4.967063, 4.967083, 
    4.967473, 4.967741, 4.967969, 4.967685, 4.967576, 4.96767, 4.967996, 
    4.96858, 4.969448, 4.970625, 4.972131, 4.973985, 4.976196, 4.978769, 
    4.981701, 4.984973, 4.988553, 4.992392, 4.996415, 5.000526, 5.0046, 
    5.008479,
  // height(29,35, 0-49)
    4.986632, 4.985251, 4.98393, 4.982677, 4.981496, 4.980392, 4.979373, 
    4.978443, 4.977607, 4.976867, 4.976226, 4.97568, 4.975222, 4.97484, 
    4.974514, 4.974512, 4.969934, 4.970024, 4.970108, 4.97006, 4.969883, 
    4.969428, 4.968791, 4.967904, 4.967138, 4.966548, 4.966253, 4.966227, 
    4.96648, 4.966601, 4.966601, 4.96651, 4.966591, 4.96687, 4.967371, 
    4.968122, 4.969146, 4.970466, 4.972102, 4.974071, 4.976381, 4.979041, 
    4.982045, 4.985377, 4.989005, 4.99288, 4.996932, 5.001062, 5.005144, 
    5.009022,
  // height(29,36, 0-49)
    4.986797, 4.985363, 4.983984, 4.98267, 4.981424, 4.980255, 4.97917, 
    4.978174, 4.977268, 4.976458, 4.97574, 4.97511, 4.974553, 4.974052, 
    4.973577, 4.973351, 4.969756, 4.969531, 4.96927, 4.968902, 4.968448, 
    4.968158, 4.967667, 4.966969, 4.966328, 4.965811, 4.965522, 4.965443, 
    4.965545, 4.965516, 4.965311, 4.965418, 4.965693, 4.96616, 4.966842, 
    4.967765, 4.968948, 4.970416, 4.972183, 4.974266, 4.976675, 4.979414, 
    4.98248, 4.985857, 4.989515, 4.993406, 4.99746, 5.001577, 5.005634, 
    5.009474,
  // height(29,37, 0-49)
    4.986938, 4.985464, 4.984036, 4.982665, 4.981359, 4.980126, 4.978973, 
    4.977904, 4.976924, 4.976033, 4.97523, 4.974505, 4.973844, 4.973222, 
    4.972605, 4.972109, 4.969525, 4.969004, 4.968421, 4.967756, 4.967048, 
    4.966916, 4.966578, 4.966092, 4.965594, 4.965162, 4.964882, 4.964739, 
    4.964676, 4.9645, 4.964114, 4.96442, 4.964892, 4.965548, 4.966413, 
    4.96751, 4.968857, 4.970472, 4.972372, 4.974567, 4.97707, 4.979882, 
    4.983001, 4.986409, 4.990077, 4.993959, 4.997983, 5.002053, 5.006046, 
    5.009804,
  // height(29,38, 0-49)
    4.987028, 4.985529, 4.984065, 4.982647, 4.981288, 4.979993, 4.978771, 
    4.977629, 4.976569, 4.975593, 4.974696, 4.973871, 4.973101, 4.972361, 
    4.971611, 4.970821, 4.969233, 4.968444, 4.967564, 4.96663, 4.965697, 
    4.965714, 4.965539, 4.96528, 4.964942, 4.964607, 4.964337, 4.964119, 
    4.963884, 4.963566, 4.96303, 4.963531, 4.964195, 4.965038, 4.966087, 
    4.967357, 4.968866, 4.970628, 4.972659, 4.974966, 4.977559, 4.980438, 
    4.983595, 4.98702, 4.990678, 4.994521, 4.998483, 5.002466, 5.006349, 
    5.009973,
  // height(29,39, 0-49)
    4.98703, 4.985528, 4.984045, 4.982595, 4.981189, 4.97984, 4.978554, 
    4.977337, 4.976196, 4.975132, 4.974139, 4.97321, 4.972332, 4.971474, 
    4.970599, 4.969515, 4.96888, 4.967854, 4.966705, 4.965531, 4.964404, 
    4.964564, 4.964558, 4.964538, 4.964377, 4.964149, 4.963889, 4.963593, 
    4.96318, 4.96273, 4.962073, 4.962762, 4.963613, 4.964639, 4.965863, 
    4.967302, 4.96897, 4.970879, 4.973037, 4.975451, 4.978129, 4.981064, 
    4.984251, 4.987672, 4.991296, 4.995074, 4.998935, 5.002787, 5.006506, 
    5.009941,
  // height(29,40, 0-49)
    4.986917, 4.985433, 4.98395, 4.982483, 4.981046, 4.979649, 4.978304, 
    4.977018, 4.975799, 4.974646, 4.973557, 4.972527, 4.971539, 4.970568, 
    4.969579, 4.968217, 4.968469, 4.967233, 4.965849, 4.964469, 4.963177, 
    4.963475, 4.963636, 4.963868, 4.963894, 4.963784, 4.963535, 4.963162, 
    4.962571, 4.962003, 4.961255, 4.962122, 4.963151, 4.964351, 4.965744, 
    4.967346, 4.969165, 4.971212, 4.973492, 4.976008, 4.978761, 4.981743, 
    4.984945, 4.988344, 4.991908, 4.995585, 4.999307, 5.002978, 5.006479, 
    5.00966,
  // height(29,41, 0-49)
    4.986656, 4.985214, 4.983752, 4.982286, 4.980833, 4.979402, 4.978008, 
    4.976662, 4.975368, 4.97413, 4.97295, 4.971819, 4.970726, 4.969647, 
    4.968551, 4.96694, 4.968, 4.966581, 4.964995, 4.963443, 4.96202, 
    4.962448, 4.962779, 4.963267, 4.963491, 4.963505, 4.963273, 4.962823, 
    4.962065, 4.961395, 4.960584, 4.96162, 4.962814, 4.964176, 4.965727, 
    4.967481, 4.969442, 4.971618, 4.974011, 4.976619, 4.979436, 4.98245, 
    4.98565, 4.989006, 4.992481, 4.996022, 4.99956, 5.002998, 5.00622, 5.00908,
  // height(29,42, 0-49)
    4.986219, 4.984845, 4.983426, 4.981982, 4.980528, 4.979081, 4.977652, 
    4.976253, 4.974894, 4.973581, 4.972313, 4.971088, 4.969896, 4.968716, 
    4.96752, 4.965698, 4.967477, 4.965904, 4.964147, 4.962456, 4.960933, 
    4.961483, 4.961984, 4.962727, 4.963152, 4.963299, 4.96309, 4.962575, 
    4.961663, 4.96091, 4.960064, 4.961257, 4.962603, 4.964114, 4.96581, 
    4.967701, 4.969793, 4.972085, 4.974578, 4.977262, 4.980129, 4.98316, 
    4.986334, 4.989621, 4.992977, 4.996344, 4.99965, 5.0028, 5.00568, 5.00815,
  // height(29,43, 0-49)
    4.985586, 4.984303, 4.982952, 4.981551, 4.980116, 4.978669, 4.977219, 
    4.975782, 4.97437, 4.97299, 4.971644, 4.970334, 4.969049, 4.967778, 
    4.966492, 4.964496, 4.966899, 4.965197, 4.963301, 4.961505, 4.959913, 
    4.960582, 4.961247, 4.96224, 4.962868, 4.963152, 4.962977, 4.962408, 
    4.961366, 4.960551, 4.959695, 4.961031, 4.962516, 4.964162, 4.965988, 
    4.968001, 4.970206, 4.972599, 4.975173, 4.977917, 4.980814, 4.983839, 
    4.986966, 4.990153, 4.993352, 4.996504, 4.999529, 5.002333, 5.004804, 
    5.006812,
  // height(29,44, 0-49)
    4.984741, 4.983572, 4.98231, 4.980974, 4.979583, 4.978152, 4.9767, 
    4.975242, 4.973791, 4.972355, 4.970943, 4.969557, 4.968193, 4.966837, 
    4.96547, 4.96334, 4.966269, 4.964459, 4.962457, 4.960586, 4.958953, 
    4.959734, 4.960559, 4.961791, 4.962621, 4.963047, 4.962915, 4.962311, 
    4.961167, 4.960318, 4.959472, 4.96094, 4.96255, 4.964314, 4.966252, 
    4.968369, 4.970668, 4.973141, 4.975777, 4.978558, 4.981461, 4.984454, 
    4.987502, 4.990557, 4.993561, 4.996449, 4.999139, 5.001537, 5.003535, 
    5.00501,
  // height(29,45, 0-49)
    4.983676, 4.982643, 4.981495, 4.980247, 4.978919, 4.977528, 4.976092, 
    4.974628, 4.973153, 4.971678, 4.970212, 4.968764, 4.967327, 4.965899, 
    4.964459, 4.962228, 4.965582, 4.963693, 4.96161, 4.959693, 4.958048, 
    4.958934, 4.95991, 4.961367, 4.962389, 4.962958, 4.962886, 4.962271, 
    4.961058, 4.960199, 4.959386, 4.960973, 4.962695, 4.964563, 4.966595, 
    4.968796, 4.971167, 4.973697, 4.976369, 4.979159, 4.982038, 4.984967, 
    4.987901, 4.990783, 4.99355, 4.996124, 4.998423, 5.000354, 5.001812, 
    5.002688,
  // height(29,46, 0-49)
    4.982392, 4.981516, 4.980502, 4.979363, 4.978121, 4.976789, 4.97539, 
    4.973942, 4.972459, 4.970959, 4.969454, 4.967954, 4.96646, 4.964968, 
    4.963467, 4.961162, 4.96484, 4.962892, 4.96076, 4.958823, 4.957186, 
    4.958171, 4.959288, 4.960949, 4.962153, 4.962865, 4.962866, 4.962266, 
    4.961024, 4.960183, 4.959423, 4.961119, 4.962938, 4.964893, 4.967002, 
    4.969267, 4.971686, 4.974245, 4.976924, 4.979692, 4.982513, 4.985339, 
    4.988117, 4.990781, 4.993258, 4.995465, 4.997318, 4.998721, 4.999578, 
    4.999793,
  // height(29,47, 0-49)
    4.980901, 4.9802, 4.979339, 4.97833, 4.977193, 4.975943, 4.9746, 
    4.973184, 4.971713, 4.970206, 4.968677, 4.967138, 4.965598, 4.964054, 
    4.962501, 4.960147, 4.964045, 4.96206, 4.959902, 4.957967, 4.956358, 
    4.957434, 4.958677, 4.960518, 4.961888, 4.96274, 4.962831, 4.962277, 
    4.961047, 4.960255, 4.959564, 4.961359, 4.963265, 4.965293, 4.967459, 
    4.969764, 4.972204, 4.974763, 4.977415, 4.980123, 4.982846, 4.985526, 
    4.988099, 4.990493, 4.992628, 4.994412, 4.995758, 4.996574, 4.996771, 
    4.996272,
  // height(29,48, 0-49)
    4.979223, 4.978709, 4.978018, 4.977159, 4.976146, 4.974998, 4.973732, 
    4.972368, 4.970926, 4.969428, 4.967888, 4.966326, 4.96475, 4.963166, 
    4.961571, 4.959184, 4.963201, 4.961198, 4.959035, 4.957121, 4.955557, 
    4.956709, 4.958065, 4.960053, 4.961572, 4.96256, 4.962756, 4.96228, 
    4.961107, 4.960392, 4.959789, 4.961674, 4.963654, 4.965738, 4.967942, 
    4.970265, 4.972701, 4.975228, 4.977816, 4.980423, 4.983, 4.985481, 
    4.987796, 4.989864, 4.991597, 4.992898, 4.993679, 4.993851, 4.993337, 
    4.992082,
  // height(29,49, 0-49)
    4.977364, 4.976999, 4.976442, 4.975697, 4.974771, 4.973678, 4.972433, 
    4.97105, 4.96955, 4.967954, 4.966277, 4.964537, 4.96275, 4.960918, 
    4.959042, 4.955583, 4.965085, 4.962095, 4.958641, 4.955575, 4.95313, 
    4.956073, 4.959288, 4.963607, 4.966753, 4.968592, 4.96859, 4.966987, 
    4.963706, 4.96112, 4.958558, 4.960826, 4.963123, 4.965455, 4.967843, 
    4.970289, 4.972789, 4.975318, 4.977843, 4.980316, 4.982681, 4.984867, 
    4.986794, 4.988374, 4.989514, 4.990113, 4.990091, 4.989372, 4.987904, 
    4.98567 ;

 totalHeight =
  // totalHeight(0,0, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // totalHeight(0,1, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // totalHeight(0,2, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // totalHeight(0,3, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // totalHeight(0,4, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // totalHeight(0,5, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // totalHeight(0,6, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // totalHeight(0,7, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // totalHeight(0,8, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // totalHeight(0,9, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // totalHeight(0,10, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // totalHeight(0,11, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // totalHeight(0,12, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // totalHeight(0,13, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // totalHeight(0,14, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // totalHeight(0,15, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // totalHeight(0,16, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // totalHeight(0,17, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // totalHeight(0,18, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // totalHeight(0,19, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // totalHeight(0,20, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 30, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // totalHeight(0,21, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 30, 5, 5, 5, 5, 5, 5, 5, 10, 
    10, 10, 10, 10, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5,
  // totalHeight(0,22, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 30, 5, 5, 5, 5, 5, 5, 10, 
    10, 10, 10, 10, 10, 10, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5,
  // totalHeight(0,23, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 30, 5, 5, 5, 5, 5, 10, 10, 
    10, 10, 10, 10, 10, 10, 10, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5,
  // totalHeight(0,24, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 30, 5, 5, 5, 5, 5, 10, 10, 
    10, 10, 10, 10, 10, 10, 10, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5,
  // totalHeight(0,25, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 30, 5, 5, 5, 5, 5, 10, 10, 
    10, 10, 10, 10, 10, 10, 10, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5,
  // totalHeight(0,26, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 30, 5, 5, 5, 5, 5, 10, 10, 
    10, 10, 10, 10, 10, 10, 10, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5,
  // totalHeight(0,27, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 30, 5, 5, 5, 5, 5, 10, 10, 
    10, 10, 10, 10, 10, 10, 10, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5,
  // totalHeight(0,28, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 30, 5, 5, 5, 5, 5, 5, 10, 
    10, 10, 10, 10, 10, 10, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5,
  // totalHeight(0,29, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 30, 5, 5, 5, 5, 5, 5, 5, 10, 
    10, 10, 10, 10, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5,
  // totalHeight(0,30, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // totalHeight(0,31, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // totalHeight(0,32, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // totalHeight(0,33, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // totalHeight(0,34, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // totalHeight(0,35, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // totalHeight(0,36, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // totalHeight(0,37, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // totalHeight(0,38, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // totalHeight(0,39, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // totalHeight(0,40, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // totalHeight(0,41, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // totalHeight(0,42, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // totalHeight(0,43, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // totalHeight(0,44, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // totalHeight(0,45, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // totalHeight(0,46, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // totalHeight(0,47, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // totalHeight(0,48, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // totalHeight(0,49, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // totalHeight(1,0, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // totalHeight(1,1, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // totalHeight(1,2, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // totalHeight(1,3, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // totalHeight(1,4, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // totalHeight(1,5, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // totalHeight(1,6, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // totalHeight(1,7, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // totalHeight(1,8, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // totalHeight(1,9, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5.000001, 5.000003, 5.000003, 5.000003, 5.000003, 5.000003, 5.000001, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // totalHeight(1,10, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 
    5.00001, 5.000023, 5.000029, 5.00003, 5.000029, 5.000023, 5.00001, 
    5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // totalHeight(1,11, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000005, 
    5.000022, 5.000071, 5.000165, 5.000208, 5.000218, 5.000208, 5.000165, 
    5.000071, 5.000022, 5.000005, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5,
  // totalHeight(1,12, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000009, 
    5.000041, 5.000161, 5.000472, 5.00103, 5.001293, 5.001361, 5.001293, 
    5.00103, 5.000472, 5.000161, 5.000041, 5.000009, 5.000001, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // totalHeight(1,13, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000013, 
    5.000065, 5.00028, 5.000989, 5.002667, 5.005479, 5.00688, 5.007271, 
    5.00688, 5.005479, 5.002667, 5.000989, 5.00028, 5.000065, 5.000013, 
    5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // totalHeight(1,14, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000016, 
    5.000087, 5.000412, 5.001609, 5.005196, 5.012874, 5.024823, 5.031068, 
    5.032917, 5.031068, 5.024823, 5.012874, 5.005196, 5.001609, 5.000412, 
    5.000087, 5.000016, 5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // totalHeight(1,15, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000018, 
    5.000104, 5.000527, 5.002232, 5.007843, 5.023126, 5.05233, 5.093832, 
    5.116333, 5.123362, 5.116333, 5.093832, 5.05233, 5.023126, 5.007843, 
    5.002232, 5.000527, 5.000104, 5.000018, 5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5,
  // totalHeight(1,16, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000016, 5.000111, 
    5.000595, 5.002696, 5.010195, 5.032046, 5.08562, 5.174296, 5.284347, 
    5.345138, 5.365025, 5.345138, 5.284347, 5.174296, 5.08562, 5.032046, 
    5.010195, 5.002696, 5.000595, 5.00011, 5.000018, 5.000002, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5,
  // totalHeight(1,17, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000013, 5.000091, 
    5.000609, 5.00287, 5.011568, 5.038834, 5.107607, 5.255316, 5.45458, 
    5.654781, 5.766831, 5.805127, 5.766831, 5.654781, 5.45458, 5.255316, 
    5.107607, 5.038834, 5.011568, 5.002866, 5.000595, 5.000104, 5.000016, 
    5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // totalHeight(1,18, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000008, 5.00006, 5.000425, 
    5.002811, 5.011596, 5.041329, 5.121252, 5.288161, 5.587032, 5.889495, 
    6.114048, 6.247925, 6.296353, 6.247925, 6.114048, 5.889495, 5.587032, 
    5.288161, 5.121252, 5.041325, 5.011568, 5.002696, 5.000527, 5.000087, 
    5.000013, 5.000001, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // totalHeight(1,19, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000003, 5.000028, 5.000218, 
    5.001533, 5.011003, 5.039038, 5.121291, 5.303221, 5.596775, 6.011393, 
    6.30257, 6.444544, 6.550306, 6.591668, 6.550305, 6.444544, 6.30257, 
    6.011393, 5.596775, 5.303215, 5.121252, 5.038834, 5.010195, 5.002232, 
    5.000412, 5.000065, 5.000009, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // totalHeight(1,20, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000014, 30, 5.039814, 
    5.109214, 5.288445, 5.596817, 5.95014, 6.326973, 6.498679, 6.541141, 
    6.600243, 6.624728, 6.600243, 6.541141, 6.498679, 6.326972, 5.950134, 
    5.596775, 5.288161, 5.107607, 5.032046, 5.007843, 5.001609, 5.00028, 
    5.000041, 5.000005, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // totalHeight(1,21, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 30, 5.108829, 
    5.260567, 5.588036, 6.011554, 6.326994, 6.546953, 6.566364, 6.535832, 
    6.558554, 6.576564, 6.558554, 6.535832, 6.566363, 6.546951, 6.326972, 
    6.011393, 5.587032, 5.255316, 5.08562, 5.023126, 5.005196, 5.000989, 
    5.000161, 5.000022, 5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // totalHeight(1,22, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 30, 5.226802, 5.467532, 
    5.892158, 6.303021, 6.498741, 6.56637, 6.621973, 6.765517, 6.920608, 
    6.987292, 6.920608, 6.765517, 6.621973, 6.566362, 6.498679, 6.30257, 
    5.889495, 5.45458, 5.174296, 5.05233, 5.012874, 5.002667, 5.000472, 
    5.000071, 5.00001, 5.000001, 5, 5, 5, 5, 5, 5, 5, 5,
  // totalHeight(1,23, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 30, 5.378377, 5.679589, 
    6.119381, 6.445471, 6.541272, 6.535846, 6.765518, 7.138705, 7.442398, 
    7.559381, 7.442398, 7.138703, 6.765517, 6.535831, 6.541141, 6.444544, 
    6.114048, 5.654781, 5.284347, 5.093832, 5.024823, 5.005479, 5.00103, 
    5.000165, 5.000023, 5.000003, 5, 5, 5, 5, 5, 5, 5, 5,
  // totalHeight(1,24, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 30, 5.461733, 5.797845, 
    6.254579, 6.551452, 6.600401, 6.558572, 6.920609, 7.442399, 7.841739, 
    7.990802, 7.841739, 7.442398, 6.920608, 6.558555, 6.600243, 6.550306, 
    6.247925, 5.766831, 5.345138, 5.116333, 5.031068, 5.00688, 5.001293, 
    5.000208, 5.000029, 5.000003, 5, 5, 5, 5, 5, 5, 5, 5,
  // totalHeight(1,25, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 30, 5.488677, 5.83798, 
    6.303374, 6.592873, 6.624895, 6.576583, 6.987293, 7.559382, 7.990802, 
    8.150589, 7.990803, 7.559381, 6.987291, 6.576564, 6.624729, 6.591668, 
    6.296353, 5.805127, 5.365025, 5.123362, 5.032917, 5.007271, 5.001361, 
    5.000218, 5.00003, 5.000003, 5, 5, 5, 5, 5, 5, 5, 5,
  // totalHeight(1,26, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 30, 5.461732, 5.797844, 
    6.254579, 6.551452, 6.600401, 6.558572, 6.920609, 7.442398, 7.841739, 
    7.990802, 7.841739, 7.442398, 6.920608, 6.558555, 6.600243, 6.550306, 
    6.247925, 5.766831, 5.345138, 5.116333, 5.031068, 5.00688, 5.001293, 
    5.000208, 5.000029, 5.000003, 5, 5, 5, 5, 5, 5, 5, 5,
  // totalHeight(1,27, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 30, 5.378368, 
    5.679588, 6.119381, 6.445471, 6.541272, 6.535846, 6.765518, 7.138705, 
    7.442398, 7.55938, 7.442398, 7.138704, 6.765517, 6.535832, 6.541142, 
    6.444544, 6.114048, 5.654781, 5.284347, 5.093832, 5.024823, 5.005479, 
    5.00103, 5.000165, 5.000023, 5.000003, 5, 5, 5, 5, 5, 5, 5, 5,
  // totalHeight(1,28, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000009, 30, 5.226734, 
    5.467518, 5.892155, 6.303021, 6.498741, 6.56637, 6.621974, 6.765516, 
    6.920608, 6.987291, 6.920608, 6.765516, 6.621973, 6.566363, 6.498679, 
    6.30257, 5.889495, 5.45458, 5.174296, 5.05233, 5.012874, 5.002667, 
    5.000472, 5.000071, 5.00001, 5.000001, 5, 5, 5, 5, 5, 5, 5, 5,
  // totalHeight(1,29, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000013, 5.00007, 30, 
    5.108382, 5.260472, 5.588021, 6.011552, 6.326994, 6.546954, 6.566364, 
    6.535832, 6.558555, 6.576563, 6.558555, 6.535832, 6.566363, 6.546951, 
    6.326972, 6.011393, 5.587032, 5.255316, 5.08562, 5.023126, 5.005196, 
    5.000989, 5.000161, 5.000022, 5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // totalHeight(1,30, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000017, 5.000138, 5.000946, 
    5.005786, 5.03459, 5.108321, 5.288314, 5.5968, 5.950139, 6.326973, 
    6.49868, 6.541142, 6.600243, 6.624728, 6.600243, 6.541142, 6.498679, 
    6.326972, 5.950134, 5.596775, 5.288161, 5.107607, 5.032046, 5.007843, 
    5.001609, 5.00028, 5.000041, 5.000005, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // totalHeight(1,31, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000005, 5.000042, 5.000306, 
    5.001886, 5.010614, 5.038951, 5.121276, 5.303219, 5.596775, 6.011393, 
    6.30257, 6.444544, 6.550306, 6.591668, 6.550306, 6.444544, 6.30257, 
    6.011393, 5.596775, 5.303215, 5.121252, 5.038834, 5.010195, 5.002232, 
    5.000412, 5.000065, 5.000009, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // totalHeight(1,32, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000009, 5.000072, 5.000477, 
    5.002755, 5.011584, 5.041328, 5.121252, 5.288161, 5.587032, 5.889495, 
    6.114048, 6.247925, 6.296353, 6.247925, 6.114048, 5.889495, 5.587032, 
    5.288161, 5.121252, 5.041325, 5.011568, 5.002696, 5.000527, 5.000087, 
    5.000013, 5.000001, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // totalHeight(1,33, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000014, 5.000097, 
    5.000602, 5.002868, 5.011568, 5.038834, 5.107607, 5.255316, 5.45458, 
    5.654781, 5.766831, 5.805127, 5.766831, 5.654781, 5.45458, 5.255316, 
    5.107607, 5.038834, 5.011568, 5.002866, 5.000595, 5.000104, 5.000016, 
    5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // totalHeight(1,34, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000017, 5.00011, 
    5.000595, 5.002696, 5.010195, 5.032046, 5.08562, 5.174296, 5.284347, 
    5.345138, 5.365025, 5.345138, 5.284347, 5.174296, 5.08562, 5.032046, 
    5.010195, 5.002696, 5.000595, 5.00011, 5.000018, 5.000002, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5,
  // totalHeight(1,35, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000018, 
    5.000104, 5.000527, 5.002232, 5.007843, 5.023126, 5.05233, 5.093832, 
    5.116333, 5.123362, 5.116333, 5.093832, 5.05233, 5.023126, 5.007843, 
    5.002232, 5.000527, 5.000104, 5.000018, 5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5,
  // totalHeight(1,36, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000016, 
    5.000087, 5.000412, 5.001609, 5.005196, 5.012874, 5.024823, 5.031068, 
    5.032917, 5.031068, 5.024823, 5.012874, 5.005196, 5.001609, 5.000412, 
    5.000087, 5.000016, 5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // totalHeight(1,37, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000013, 
    5.000065, 5.00028, 5.000989, 5.002667, 5.005479, 5.00688, 5.007271, 
    5.00688, 5.005479, 5.002667, 5.000989, 5.00028, 5.000065, 5.000013, 
    5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // totalHeight(1,38, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000009, 
    5.000041, 5.000161, 5.000472, 5.00103, 5.001293, 5.001361, 5.001293, 
    5.00103, 5.000472, 5.000161, 5.000041, 5.000009, 5.000001, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // totalHeight(1,39, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000005, 
    5.000022, 5.000071, 5.000165, 5.000208, 5.000218, 5.000208, 5.000165, 
    5.000071, 5.000022, 5.000005, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5,
  // totalHeight(1,40, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 
    5.00001, 5.000023, 5.000029, 5.00003, 5.000029, 5.000023, 5.00001, 
    5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // totalHeight(1,41, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5.000001, 5.000003, 5.000003, 5.000003, 5.000003, 5.000003, 5.000001, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // totalHeight(1,42, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // totalHeight(1,43, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // totalHeight(1,44, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // totalHeight(1,45, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // totalHeight(1,46, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // totalHeight(1,47, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // totalHeight(1,48, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // totalHeight(1,49, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // totalHeight(2,0, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // totalHeight(2,1, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // totalHeight(2,2, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // totalHeight(2,3, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5.000001, 5.000001, 5.000001, 5.000001, 5.000001, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // totalHeight(2,4, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 
    5.000003, 5.000006, 5.000008, 5.000009, 5.000008, 5.000006, 5.000003, 
    5.000001, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // totalHeight(2,5, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 
    5.000003, 5.000009, 5.000018, 5.00003, 5.000037, 5.000041, 5.000037, 
    5.00003, 5.000018, 5.000009, 5.000003, 5.000001, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // totalHeight(2,6, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000008, 
    5.00002, 5.000044, 5.000084, 5.000135, 5.000167, 5.000179, 5.000167, 
    5.000135, 5.000084, 5.000044, 5.00002, 5.000008, 5.000002, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // totalHeight(2,7, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000004, 5.000013, 
    5.000036, 5.000087, 5.000192, 5.000359, 5.000562, 5.000698, 5.000745, 
    5.000698, 5.000562, 5.000359, 5.000192, 5.000087, 5.000036, 5.000013, 
    5.000004, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // totalHeight(2,8, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000005, 
    5.000019, 5.000055, 5.000149, 5.000361, 5.000768, 5.001396, 5.002146, 
    5.002654, 5.002829, 5.002654, 5.002146, 5.001396, 5.000768, 5.000361, 
    5.000149, 5.000055, 5.000019, 5.000005, 5.000001, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5,
  // totalHeight(2,9, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000007, 5.000025, 
    5.00008, 5.00023, 5.000596, 5.001375, 5.002819, 5.004971, 5.00749, 
    5.009201, 5.009799, 5.009201, 5.00749, 5.004971, 5.002819, 5.001375, 
    5.000596, 5.00023, 5.00008, 5.000025, 5.000007, 5.000001, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5,
  // totalHeight(2,10, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000008, 5.000031, 
    5.000104, 5.000319, 5.000876, 5.002162, 5.004771, 5.009418, 5.016093, 
    5.023739, 5.028931, 5.030761, 5.028931, 5.023739, 5.016093, 5.009418, 
    5.004771, 5.002162, 5.000876, 5.000319, 5.000104, 5.000031, 5.000008, 
    5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // totalHeight(2,11, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.00001, 5.000034, 
    5.000126, 5.000408, 5.001172, 5.003046, 5.007127, 5.014987, 5.028435, 
    5.046975, 5.067611, 5.08152, 5.086449, 5.08152, 5.067611, 5.046975, 
    5.028435, 5.014987, 5.007127, 5.003045, 5.001171, 5.000405, 5.000127, 
    5.000036, 5.00001, 5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // totalHeight(2,12, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000009, 5.000036, 5.000136, 
    5.000466, 5.001442, 5.003905, 5.00958, 5.021203, 5.042273, 5.076715, 
    5.121716, 5.169673, 5.201324, 5.212531, 5.201324, 5.169673, 5.121716, 
    5.076715, 5.042273, 5.021201, 5.009576, 5.003897, 5.00143, 5.000474, 
    5.000143, 5.000039, 5.00001, 5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // totalHeight(2,13, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000008, 5.000033, 5.000133, 
    5.000481, 5.00157, 5.004634, 5.011772, 5.027131, 5.05641, 5.105655, 
    5.181499, 5.273223, 5.364344, 5.422204, 5.4425, 5.422204, 5.364344, 
    5.273223, 5.181498, 5.105653, 5.056403, 5.02711, 5.011728, 5.004572, 
    5.001609, 5.000513, 5.000149, 5.000039, 5.00001, 5.000002, 5, 5, 5, 5, 5, 
    5, 5, 5, 5,
  // totalHeight(2,14, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000007, 5.000029, 5.000118, 5.000446, 
    5.001536, 5.004781, 5.013485, 5.031936, 5.068588, 5.132482, 5.229629, 
    5.367397, 5.516597, 5.650199, 5.73082, 5.75868, 5.73082, 5.650199, 
    5.516597, 5.367393, 5.229616, 5.132443, 5.068489, 5.031737, 5.013205, 
    5.004946, 5.001672, 5.000513, 5.000143, 5.000036, 5.000008, 5.000001, 5, 
    5, 5, 5, 5, 5, 5, 5,
  // totalHeight(2,15, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000004, 5.000021, 5.000093, 5.000368, 
    5.001338, 5.004398, 5.013077, 5.035445, 5.07743, 5.152986, 5.270136, 
    5.425341, 5.623005, 5.808567, 5.954159, 6.038265, 6.066943, 6.038265, 
    5.954158, 5.808562, 5.622989, 5.425284, 5.269968, 5.152572, 5.076609, 
    5.034278, 5.01373, 5.004946, 5.001609, 5.000474, 5.000127, 5.000031, 
    5.000007, 5.000001, 5, 5, 5, 5, 5, 5, 5,
  // totalHeight(2,16, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000014, 5.000063, 5.000268, 5.001024, 
    5.003561, 5.011195, 5.031907, 5.083897, 5.166404, 5.297246, 5.471339, 
    5.663941, 5.881144, 6.054009, 6.170801, 6.238191, 6.261086, 6.23819, 
    6.170798, 6.053992, 5.881079, 5.663725, 5.470706, 5.295689, 5.163324, 
    5.079466, 5.034278, 5.013205, 5.004572, 5.00143, 5.000405, 5.000104, 
    5.000025, 5.000005, 5, 5, 5, 5, 5, 5, 5,
  // totalHeight(2,17, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000008, 5.000038, 5.000165, 5.00067, 
    5.002472, 5.008275, 5.024992, 5.068762, 5.178341, 5.314689, 5.498798, 
    5.701071, 5.878989, 6.057094, 6.174425, 6.241654, 6.28508, 6.300066, 
    6.285078, 6.24164, 6.174369, 6.056881, 5.878283, 5.699006, 5.493689, 
    5.304491, 5.163324, 5.076609, 5.031737, 5.011728, 5.003897, 5.001171, 
    5.000319, 5.00008, 5.000019, 5.000004, 5, 5, 5, 5, 5, 5,
  // totalHeight(2,18, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5.000003, 5.000017, 5.000082, 5.000356, 5.001401, 
    5.005028, 5.016359, 5.047846, 5.129076, 5.339933, 5.523062, 5.725195, 
    5.900149, 6.010222, 6.107472, 6.153584, 6.174073, 6.196599, 6.204854, 
    6.196589, 6.174033, 6.153419, 6.106858, 6.008182, 5.894237, 5.710595, 
    5.493689, 5.295689, 5.152572, 5.068489, 5.02711, 5.009576, 5.003045, 
    5.000876, 5.00023, 5.000055, 5.000013, 5.000002, 5, 5, 5, 5, 5,
  // totalHeight(2,19, 0-49)
    5, 5, 5, 5, 5, 5, 5.000001, 5.000007, 5.000029, 5.000135, 5.000575, 
    5.002245, 5.008015, 5.025926, 5.074886, 5.206708, 5.580922, 5.772137, 
    5.930871, 6.024444, 6.039964, 6.04226, 6.020387, 6.004436, 6.009708, 
    6.012484, 6.009684, 6.004327, 6.019951, 6.040654, 6.034697, 6.009424, 
    5.894236, 5.699005, 5.470706, 5.269968, 5.132443, 5.056403, 5.021201, 
    5.007127, 5.002162, 5.000596, 5.000149, 5.000036, 5.000008, 5.000001, 5, 
    5, 5, 5,
  // totalHeight(2,20, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5.000001, 5.00001, 5.000042, 5.000171, 5.000613, 
    5.001966, 5.005518, 5.013143, 30, 6.070654, 6.10031, 6.109229, 6.073961, 
    5.989838, 5.897338, 5.812802, 5.764136, 5.750331, 5.746961, 5.750273, 
    5.763871, 5.811723, 5.893331, 5.976495, 6.034697, 6.008182, 5.878282, 
    5.663725, 5.425284, 5.229616, 5.105653, 5.042273, 5.014987, 5.004771, 
    5.001375, 5.000361, 5.000087, 5.00002, 5.000003, 5, 5, 5, 5,
  // totalHeight(2,21, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5.000003, 5.000014, 5.000054, 5.000195, 5.00063, 
    5.001772, 5.004181, 30, 6.513035, 6.426273, 6.282675, 6.110457, 5.917133, 
    5.702082, 5.514227, 5.387189, 5.318944, 5.296926, 5.318848, 5.386738, 
    5.51234, 5.694969, 5.893331, 6.040654, 6.106857, 6.056882, 5.88108, 
    5.622988, 5.367393, 5.181498, 5.076715, 5.028435, 5.009418, 5.002819, 
    5.000768, 5.000192, 5.000044, 5.000009, 5.000001, 5, 5, 5,
  // totalHeight(2,22, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000004, 5.000016, 5.000055, 5.000182, 
    5.000515, 5.001205, 30, 6.890601, 6.696692, 6.413081, 6.125101, 5.847679, 
    5.523096, 5.231614, 5.02129, 4.898302, 4.858558, 4.898164, 5.020628, 
    5.228783, 5.512339, 5.811723, 6.019951, 6.153419, 6.174369, 6.053992, 
    5.808561, 5.516597, 5.273223, 5.121716, 5.046975, 5.016093, 5.004971, 
    5.001396, 5.000359, 5.000084, 5.000018, 5.000003, 5, 5, 5,
  // totalHeight(2,23, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000004, 5.000016, 5.000049, 5.000141, 
    5.000327, 30, 7.175317, 6.901651, 6.513165, 6.143483, 5.81144, 5.400992, 
    5.024344, 4.753988, 4.602839, 4.55656, 4.602668, 4.753143, 5.020628, 
    5.386737, 5.76387, 6.004326, 6.174033, 6.241639, 6.170797, 5.954158, 
    5.650199, 5.364344, 5.169673, 5.067611, 5.023739, 5.00749, 5.002146, 
    5.000562, 5.000135, 5.00003, 5.000006, 5.000001, 5, 5,
  // totalHeight(2,24, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000006, 5.00002, 5.000057, 5.000128, 
    30, 7.33971, 7.028852, 6.586917, 6.171556, 5.805634, 5.335411, 4.902411, 
    4.603594, 4.448595, 4.40392, 4.448415, 4.602663, 4.89816, 5.318843, 
    5.750269, 6.009683, 6.196589, 6.285078, 6.23819, 6.038265, 5.73082, 
    5.422204, 5.201324, 5.08152, 5.028931, 5.009201, 5.002654, 5.000698, 
    5.000167, 5.000037, 5.000008, 5.000001, 5, 5,
  // totalHeight(2,25, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000003, 5.000013, 5.000041, 5.000108, 
    5.000237, 30, 7.394997, 7.072412, 6.612961, 6.182293, 5.805012, 5.31426, 
    4.862948, 4.55748, 4.40407, 4.360934, 4.403889, 4.556526, 4.858529, 
    5.296904, 5.746947, 6.012478, 6.204852, 6.300065, 6.261086, 6.066943, 
    5.75868, 5.4425, 5.212531, 5.086449, 5.030761, 5.009799, 5.002829, 
    5.000745, 5.000179, 5.000041, 5.000009, 5.000001, 5, 5,
  // totalHeight(2,26, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000003, 5.000014, 5.000048, 5.000146, 
    5.00039, 5.000851, 30, 7.33743, 7.027562, 6.586339, 6.171353, 5.805575, 
    5.335398, 4.902407, 4.603593, 4.448595, 4.403919, 4.448415, 4.602663, 
    4.898159, 5.318843, 5.750269, 6.009683, 6.196589, 6.285078, 6.23819, 
    6.038265, 5.73082, 5.422204, 5.201324, 5.08152, 5.028931, 5.009201, 
    5.002654, 5.000698, 5.000167, 5.000037, 5.000008, 5.000001, 5, 5,
  // totalHeight(2,27, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5.000003, 5.000013, 5.000049, 5.000171, 5.000519, 
    5.001362, 5.002976, 30, 7.16783, 6.897426, 6.511255, 6.142797, 5.811236, 
    5.40094, 5.024333, 4.753986, 4.602839, 4.55656, 4.602669, 4.753144, 
    5.020627, 5.386737, 5.76387, 6.004327, 6.174033, 6.24164, 6.170797, 
    5.954158, 5.650199, 5.364344, 5.169673, 5.067611, 5.023739, 5.00749, 
    5.002146, 5.000562, 5.000135, 5.00003, 5.000006, 5.000001, 5, 5,
  // totalHeight(2,28, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5.000002, 5.00001, 5.000044, 5.000165, 5.000557, 
    5.001666, 5.004333, 5.009483, 30, 6.869401, 6.684888, 6.407736, 6.123141, 
    5.847076, 5.522937, 5.231577, 5.021283, 4.898301, 4.858558, 4.898164, 
    5.020629, 5.228784, 5.51234, 5.811723, 6.019951, 6.153419, 6.174369, 
    6.053992, 5.808561, 5.516597, 5.273223, 5.121716, 5.046975, 5.016093, 
    5.004971, 5.001396, 5.000359, 5.000084, 5.000018, 5.000003, 5, 5, 5,
  // totalHeight(2,29, 0-49)
    5, 5, 5, 5, 5, 5, 5.000001, 5.000007, 5.000031, 5.00013, 5.000485, 
    5.001624, 5.004813, 5.012438, 5.027185, 30, 6.458423, 6.39655, 6.269349, 
    6.105521, 5.915573, 5.701647, 5.514119, 5.387164, 5.318938, 5.296925, 
    5.318848, 5.386738, 5.51234, 5.694969, 5.893331, 6.040654, 6.106858, 
    6.056882, 5.88108, 5.622988, 5.367393, 5.181498, 5.076715, 5.028435, 
    5.009418, 5.002819, 5.000768, 5.000192, 5.000044, 5.000009, 5.000001, 5, 
    5, 5,
  // totalHeight(2,30, 0-49)
    5, 5, 5, 5, 5, 5, 5.000004, 5.000019, 5.000091, 5.000392, 5.001544, 
    5.005568, 5.018255, 5.053765, 5.13902, 5.339774, 5.824156, 5.992731, 
    6.068674, 6.060568, 5.985876, 5.89627, 5.812539, 5.764076, 5.750317, 
    5.746958, 5.750272, 5.763871, 5.811723, 5.893331, 5.976495, 6.034697, 
    6.008182, 5.878283, 5.663725, 5.425284, 5.229616, 5.105653, 5.042273, 
    5.014987, 5.004771, 5.001375, 5.000361, 5.000087, 5.00002, 5.000003, 5, 
    5, 5, 5,
  // totalHeight(2,31, 0-49)
    5, 5, 5, 5, 5, 5, 5.000002, 5.000012, 5.000059, 5.000257, 5.001028, 
    5.003737, 5.01235, 5.036781, 5.097425, 5.235366, 5.544514, 5.750298, 
    5.92068, 6.020491, 6.03864, 6.041875, 6.020286, 6.00441, 6.009703, 
    6.012483, 6.009684, 6.004327, 6.019951, 6.040655, 6.034697, 6.009424, 
    5.894237, 5.699006, 5.470706, 5.269968, 5.132443, 5.056403, 5.021201, 
    5.007127, 5.002162, 5.000596, 5.000149, 5.000036, 5.000008, 5.000001, 5, 
    5, 5, 5,
  // totalHeight(2,32, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5.000005, 5.000028, 5.000126, 5.000518, 5.00194, 
    5.006609, 5.020349, 5.056161, 5.140028, 5.324083, 5.513662, 5.720868, 
    5.898491, 6.009674, 6.107315, 6.153543, 6.174064, 6.196596, 6.204853, 
    6.196589, 6.174033, 6.153419, 6.106858, 6.008182, 5.894237, 5.710595, 
    5.493689, 5.295689, 5.152572, 5.068489, 5.02711, 5.009576, 5.003045, 
    5.000876, 5.00023, 5.000055, 5.000013, 5.000002, 5, 5, 5, 5, 5,
  // totalHeight(2,33, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000011, 5.000051, 5.000216, 5.000844, 
    5.002991, 5.009605, 5.02779, 5.072512, 5.172647, 5.311225, 5.497193, 
    5.700458, 5.878788, 6.057036, 6.17441, 6.241651, 6.28508, 6.300066, 
    6.285078, 6.241639, 6.174369, 6.056882, 5.878283, 5.699006, 5.493689, 
    5.304491, 5.163324, 5.076609, 5.031737, 5.011728, 5.003897, 5.001171, 
    5.000319, 5.00008, 5.000019, 5.000004, 5, 5, 5, 5, 5, 5,
  // totalHeight(2,34, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5.000003, 5.000018, 5.000078, 5.000318, 5.001177, 
    5.003963, 5.012051, 5.033063, 5.082146, 5.165304, 5.29673, 5.471141, 
    5.663877, 5.881125, 6.054005, 6.170801, 6.238191, 6.261086, 6.238191, 
    6.170798, 6.053992, 5.88108, 5.663725, 5.470706, 5.295689, 5.163324, 
    5.079466, 5.034278, 5.013205, 5.004572, 5.00143, 5.000405, 5.000104, 
    5.000025, 5.000005, 5, 5, 5, 5, 5, 5, 5,
  // totalHeight(2,35, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000006, 5.000025, 5.000106, 5.000411, 
    5.001449, 5.004638, 5.0134, 5.034968, 5.077124, 5.152843, 5.270081, 
    5.425323, 5.623, 5.808566, 5.954159, 6.038265, 6.066944, 6.038265, 
    5.954159, 5.808562, 5.622989, 5.425284, 5.269968, 5.152572, 5.076609, 
    5.034278, 5.01373, 5.004946, 5.001609, 5.000474, 5.000127, 5.000031, 
    5.000007, 5.000001, 5, 5, 5, 5, 5, 5, 5,
  // totalHeight(2,36, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000007, 5.000031, 5.000127, 
    5.000473, 5.001596, 5.004863, 5.013367, 5.031859, 5.068552, 5.132469, 
    5.229624, 5.367395, 5.516597, 5.650199, 5.73082, 5.75868, 5.73082, 
    5.650199, 5.516597, 5.367393, 5.229616, 5.132443, 5.068489, 5.031737, 
    5.013205, 5.004946, 5.001672, 5.000513, 5.000143, 5.000036, 5.000008, 
    5.000001, 5, 5, 5, 5, 5, 5, 5, 5,
  // totalHeight(2,37, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000009, 5.000036, 5.000139, 
    5.000494, 5.001589, 5.004607, 5.011755, 5.027123, 5.056408, 5.105654, 
    5.181498, 5.273223, 5.364344, 5.422204, 5.4425, 5.422204, 5.364344, 
    5.273223, 5.181498, 5.105653, 5.056403, 5.02711, 5.011728, 5.004572, 
    5.001609, 5.000513, 5.000149, 5.000039, 5.00001, 5.000002, 5, 5, 5, 5, 5, 
    5, 5, 5, 5,
  // totalHeight(2,38, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.00001, 5.000037, 5.000138, 
    5.00047, 5.001437, 5.003901, 5.009578, 5.021202, 5.042273, 5.076715, 
    5.121716, 5.169673, 5.201324, 5.212531, 5.201324, 5.169673, 5.121716, 
    5.076715, 5.042273, 5.021201, 5.009576, 5.003897, 5.00143, 5.000474, 
    5.000143, 5.000039, 5.00001, 5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // totalHeight(2,39, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.00001, 5.000034, 
    5.000126, 5.000407, 5.001172, 5.003045, 5.007127, 5.014987, 5.028435, 
    5.046975, 5.067611, 5.08152, 5.086449, 5.08152, 5.067611, 5.046975, 
    5.028435, 5.014987, 5.007127, 5.003045, 5.001171, 5.000405, 5.000127, 
    5.000036, 5.00001, 5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // totalHeight(2,40, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000008, 5.000031, 
    5.000104, 5.000319, 5.000876, 5.002162, 5.004771, 5.009418, 5.016093, 
    5.023739, 5.028931, 5.030761, 5.028931, 5.023739, 5.016093, 5.009418, 
    5.004771, 5.002162, 5.000876, 5.000319, 5.000104, 5.000031, 5.000008, 
    5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // totalHeight(2,41, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000007, 5.000025, 
    5.00008, 5.00023, 5.000596, 5.001375, 5.002819, 5.004971, 5.00749, 
    5.009201, 5.009799, 5.009201, 5.00749, 5.004971, 5.002819, 5.001375, 
    5.000596, 5.00023, 5.00008, 5.000025, 5.000007, 5.000001, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5,
  // totalHeight(2,42, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000005, 
    5.000019, 5.000055, 5.000149, 5.000361, 5.000768, 5.001396, 5.002146, 
    5.002654, 5.002829, 5.002654, 5.002146, 5.001396, 5.000768, 5.000361, 
    5.000149, 5.000055, 5.000019, 5.000005, 5.000001, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5,
  // totalHeight(2,43, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000004, 5.000013, 
    5.000036, 5.000087, 5.000192, 5.000359, 5.000562, 5.000698, 5.000745, 
    5.000698, 5.000562, 5.000359, 5.000192, 5.000087, 5.000036, 5.000013, 
    5.000004, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // totalHeight(2,44, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000008, 
    5.00002, 5.000044, 5.000084, 5.000135, 5.000167, 5.000179, 5.000167, 
    5.000135, 5.000084, 5.000044, 5.00002, 5.000008, 5.000002, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // totalHeight(2,45, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 
    5.000003, 5.000009, 5.000018, 5.00003, 5.000037, 5.000041, 5.000037, 
    5.00003, 5.000018, 5.000009, 5.000003, 5.000001, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // totalHeight(2,46, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 
    5.000003, 5.000006, 5.000008, 5.000009, 5.000008, 5.000006, 5.000003, 
    5.000001, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // totalHeight(2,47, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5.000001, 5.000001, 5.000001, 5.000001, 5.000001, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // totalHeight(2,48, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // totalHeight(2,49, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // totalHeight(3,0, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 
    5.000003, 5.000006, 5.00001, 5.000014, 5.000018, 5.000019, 5.000018, 
    5.000014, 5.00001, 5.000006, 5.000003, 5.000001, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // totalHeight(3,1, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000007, 
    5.000014, 5.000024, 5.000038, 5.000054, 5.000065, 5.000069, 5.000065, 
    5.000054, 5.000038, 5.000024, 5.000014, 5.000007, 5.000002, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // totalHeight(3,2, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000005, 
    5.000013, 5.000025, 5.000051, 5.000089, 5.000139, 5.000192, 5.00023, 
    5.000245, 5.00023, 5.000192, 5.000139, 5.000089, 5.000051, 5.000025, 
    5.000013, 5.000005, 5.000001, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // totalHeight(3,3, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000003, 5.000008, 5.00002, 
    5.000045, 5.000092, 5.000175, 5.000303, 5.000471, 5.000645, 5.000771, 
    5.000815, 5.000771, 5.000645, 5.000471, 5.000303, 5.000175, 5.000092, 
    5.000045, 5.00002, 5.000008, 5.000003, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5,
  // totalHeight(3,4, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000004, 5.000012, 5.00003, 
    5.00007, 5.000153, 5.000309, 5.000576, 5.000975, 5.001488, 5.002019, 
    5.0024, 5.002537, 5.0024, 5.002019, 5.001488, 5.000975, 5.000576, 
    5.000309, 5.000153, 5.00007, 5.00003, 5.000012, 5.000004, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5,
  // totalHeight(3,5, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000005, 5.000016, 
    5.000041, 5.000101, 5.000232, 5.000495, 5.000975, 5.001767, 5.002935, 
    5.004404, 5.005916, 5.006993, 5.007383, 5.006993, 5.005916, 5.004404, 
    5.002935, 5.001767, 5.000974, 5.000495, 5.000232, 5.000101, 5.000041, 
    5.000016, 5.000005, 5.000001, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // totalHeight(3,6, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000007, 5.00002, 5.000052, 
    5.000135, 5.000328, 5.000727, 5.001502, 5.002871, 5.005065, 5.008235, 
    5.012152, 5.016148, 5.018981, 5.020005, 5.018981, 5.016148, 5.012152, 
    5.008235, 5.005065, 5.00287, 5.001501, 5.000726, 5.000327, 5.000136, 
    5.000052, 5.00002, 5.000007, 5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // totalHeight(3,7, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000008, 5.000022, 5.000062, 
    5.000168, 5.000426, 5.000994, 5.002136, 5.004256, 5.007876, 5.013505, 
    5.021459, 5.0311, 5.040833, 5.047673, 5.050141, 5.047673, 5.040833, 
    5.0311, 5.021459, 5.013503, 5.007874, 5.004254, 5.00213, 5.000989, 
    5.000427, 5.000171, 5.000064, 5.000023, 5.000008, 5.000002, 5, 5, 5, 5, 
    5, 5, 5, 5, 5,
  // totalHeight(3,8, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000008, 5.000023, 5.000071, 
    5.000197, 5.000516, 5.001256, 5.002826, 5.005837, 5.011214, 5.020035, 
    5.033278, 5.051542, 5.073155, 5.094623, 5.109491, 5.114835, 5.109491, 
    5.094623, 5.073154, 5.05154, 5.033274, 5.020027, 5.011199, 5.005819, 
    5.002808, 5.001259, 5.000525, 5.000204, 5.000074, 5.000025, 5.000008, 
    5.000002, 5, 5, 5, 5, 5, 5, 5, 5,
  // totalHeight(3,9, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000008, 5.000024, 5.000072, 5.000215, 
    5.000583, 5.001472, 5.003447, 5.007477, 5.01482, 5.027332, 5.046957, 
    5.07516, 5.112832, 5.155911, 5.197577, 5.225729, 5.235758, 5.225728, 
    5.197576, 5.155908, 5.112823, 5.075142, 5.046923, 5.027278, 5.014745, 
    5.00741, 5.003462, 5.001504, 5.000608, 5.000228, 5.00008, 5.000026, 
    5.000009, 5.000002, 5, 5, 5, 5, 5, 5, 5,
  // totalHeight(3,10, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000007, 5.000022, 5.000071, 5.000216, 
    5.00061, 5.001602, 5.003899, 5.008797, 5.018371, 5.034782, 5.061243, 
    5.100461, 5.15364, 5.221577, 5.295402, 5.36382, 5.408352, 5.423996, 
    5.408351, 5.363815, 5.29539, 5.221547, 5.153577, 5.100338, 5.061041, 
    5.034512, 5.018124, 5.008841, 5.004006, 5.001688, 5.000662, 5.000242, 
    5.000082, 5.000026, 5.000008, 5.000002, 5, 5, 5, 5, 5, 5,
  // totalHeight(3,11, 0-49)
    5, 5, 5, 5, 5, 5, 5.000001, 5.000006, 5.000021, 5.000064, 5.000203, 
    5.000594, 5.001617, 5.004089, 5.009582, 5.020787, 5.04175, 5.075024, 
    5.125049, 5.193873, 5.280046, 5.383638, 5.488432, 5.579867, 5.636599, 
    5.656176, 5.636593, 5.57985, 5.488389, 5.383534, 5.279824, 5.193449, 
    5.124352, 5.074101, 5.040899, 5.020916, 5.009921, 5.004369, 5.001788, 
    5.000681, 5.000242, 5.00008, 5.000025, 5.000008, 5.000002, 5, 5, 5, 5, 5,
  // totalHeight(3,12, 0-49)
    5, 5, 5, 5, 5, 5, 5.000005, 5.000017, 5.000055, 5.000177, 5.000535, 
    5.001513, 5.003968, 5.009657, 5.021753, 5.045288, 5.087358, 5.14761, 
    5.230261, 5.333305, 5.449304, 5.57871, 5.698251, 5.795069, 5.852182, 
    5.871558, 5.852166, 5.795019, 5.698119, 5.578391, 5.448622, 5.331985, 
    5.228084, 5.144711, 5.084641, 5.045663, 5.022761, 5.010503, 5.004496, 
    5.001788, 5.000662, 5.000228, 5.000074, 5.000023, 5.000007, 5.000001, 5, 
    5, 5, 5,
  // totalHeight(3,13, 0-49)
    5, 5, 5, 5, 5, 5.000002, 5.000013, 5.000043, 5.000142, 5.000446, 
    5.001304, 5.003549, 5.008974, 5.021013, 5.045398, 5.090425, 5.167326, 
    5.262846, 5.378967, 5.506453, 5.631666, 5.760675, 5.867614, 5.947062, 
    5.992007, 6.007091, 5.991964, 5.946927, 5.867256, 5.75981, 5.629799, 
    5.502812, 5.372893, 5.25464, 5.159427, 5.091476, 5.048205, 5.023404, 
    5.010503, 5.004369, 5.001688, 5.000608, 5.000204, 5.000064, 5.00002, 
    5.000005, 5, 5, 5, 5,
  // totalHeight(3,14, 0-49)
    5, 5, 5, 5, 5.000001, 5.000009, 5.000031, 5.000105, 5.00034, 5.001029, 
    5.002908, 5.007648, 5.018635, 5.041913, 5.086556, 5.164249, 5.291772, 
    5.421392, 5.55587, 5.681244, 5.783919, 5.882294, 5.952684, 5.99908, 
    6.024866, 6.03354, 6.024758, 5.998743, 5.951796, 5.880162, 5.77933, 
    5.672307, 5.540854, 5.400769, 5.271254, 5.167127, 5.093842, 5.048205, 
    5.022761, 5.009921, 5.004006, 5.001504, 5.000525, 5.000171, 5.000052, 
    5.000016, 5.000004, 5, 5, 5,
  // totalHeight(3,15, 0-49)
    5, 5, 5, 5, 5.000005, 5.00002, 5.000069, 5.000233, 5.000735, 5.002163, 
    5.005921, 5.015044, 5.035314, 5.076136, 5.14962, 5.26931, 5.461556, 
    5.608839, 5.731626, 5.821412, 5.873544, 5.920516, 5.942305, 5.950413, 
    5.955587, 5.957473, 5.955333, 5.949632, 5.940266, 5.915689, 5.863268, 
    5.801664, 5.698636, 5.56323, 5.414839, 5.276899, 5.167127, 5.091476, 
    5.045663, 5.020916, 5.00884, 5.003462, 5.001259, 5.000427, 5.000136, 
    5.000041, 5.000012, 5.000003, 5, 5,
  // totalHeight(3,16, 0-49)
    5, 5, 5, 5.000002, 5.000011, 5.000041, 5.000143, 5.000468, 5.001436, 
    5.004103, 5.010897, 5.026792, 5.060598, 5.124972, 5.232549, 5.396155, 
    5.662586, 5.799902, 5.878317, 5.906157, 5.892824, 5.879972, 5.850737, 
    5.821409, 5.806584, 5.801819, 5.806024, 5.819709, 5.846377, 5.869823, 
    5.871604, 5.866385, 5.813318, 5.711125, 5.5706, 5.414839, 5.271254, 
    5.159427, 5.084641, 5.040899, 5.018124, 5.00741, 5.002808, 5.000989, 
    5.000327, 5.000101, 5.00003, 5.000008, 5.000001, 5,
  // totalHeight(3,17, 0-49)
    5, 5, 5.000001, 5.000005, 5.000021, 5.000075, 5.000259, 5.000828, 
    5.002479, 5.006911, 5.017881, 5.042683, 5.093165, 5.18362, 5.322259, 
    5.521502, 5.866402, 5.969814, 5.983183, 5.936786, 5.854723, 5.780489, 
    5.701207, 5.636169, 5.601222, 5.58957, 5.600065, 5.632699, 5.692458, 
    5.76054, 5.814003, 5.863031, 5.867137, 5.816883, 5.711125, 5.56323, 
    5.400769, 5.25464, 5.144711, 5.0741, 5.034512, 5.014745, 5.005819, 
    5.00213, 5.000726, 5.000232, 5.00007, 5.00002, 5.000005, 5,
  // totalHeight(3,18, 0-49)
    5, 5, 5.000002, 5.000009, 5.000031, 5.000117, 5.000395, 5.001246, 
    5.003667, 5.010052, 5.025521, 5.059556, 5.126149, 5.238306, 5.394081, 
    5.615667, 6.035935, 6.101533, 6.04922, 5.929343, 5.78085, 5.644381, 
    5.515065, 5.414158, 5.357251, 5.337825, 5.354997, 5.407474, 5.498516, 
    5.607554, 5.707836, 5.802571, 5.86004, 5.867137, 5.813318, 5.698636, 
    5.540854, 5.372893, 5.228083, 5.124352, 5.061041, 5.027278, 5.011199, 
    5.004254, 5.001501, 5.000495, 5.000153, 5.000045, 5.000013, 5.000002,
  // totalHeight(3,19, 0-49)
    5, 5, 5.000002, 5.000011, 5.000038, 5.00014, 5.000471, 5.001475, 
    5.004326, 5.011827, 5.029943, 5.069492, 5.145236, 5.266404, 5.417098, 
    5.657688, 6.133231, 6.183744, 6.085767, 5.90326, 5.691944, 5.490312, 
    5.308599, 5.169163, 5.086947, 5.058302, 5.082806, 5.156998, 5.279012, 
    5.426208, 5.569045, 5.70021, 5.80257, 5.863031, 5.866385, 5.801664, 
    5.672307, 5.502812, 5.331985, 5.193449, 5.100338, 5.046923, 5.020027, 
    5.007874, 5.00287, 5.000974, 5.000309, 5.000092, 5.000025, 5.000007,
  // totalHeight(3,20, 0-49)
    5, 5, 5.000001, 5.000006, 5.000022, 5.000076, 5.000246, 5.000745, 
    5.002099, 5.005454, 5.012992, 5.028082, 5.054316, 5.092286, 5.134862, 30, 
    6.537839, 6.444597, 6.224334, 5.931908, 5.627497, 5.341224, 5.09673, 
    4.91181, 4.799217, 4.759322, 4.791854, 4.890079, 5.043821, 5.226887, 
    5.408791, 5.569041, 5.707834, 5.814003, 5.871604, 5.863268, 5.779329, 
    5.629799, 5.448622, 5.279824, 5.153577, 5.075142, 5.033274, 5.013503, 
    5.005065, 5.001767, 5.000576, 5.000175, 5.000051, 5.000014,
  // totalHeight(3,21, 0-49)
    5, 5, 5, 5.000002, 5.000011, 5.000037, 5.000119, 5.000364, 5.001029, 
    5.002694, 5.006472, 5.01416, 5.027897, 5.048741, 5.073972, 30, 6.715348, 
    6.582877, 6.306049, 5.934135, 5.539999, 5.157746, 4.834559, 4.587932, 
    4.433352, 4.378251, 4.422956, 4.55676, 4.757838, 4.992012, 5.226871, 
    5.426194, 5.607547, 5.760535, 5.869822, 5.915688, 5.880161, 5.75981, 
    5.578391, 5.383534, 5.221547, 5.112823, 5.05154, 5.021459, 5.008235, 
    5.002935, 5.000975, 5.000303, 5.000089, 5.000024,
  // totalHeight(3,22, 0-49)
    5, 5, 5, 5, 5.000004, 5.000016, 5.000052, 5.00016, 5.000462, 5.001224, 
    5.002986, 5.006641, 5.013321, 5.023751, 5.036767, 30, 6.819324, 6.665093, 
    6.350619, 5.917248, 5.445622, 4.973551, 4.571023, 4.255342, 4.050066, 
    3.976002, 4.036703, 4.214768, 4.470624, 4.757758, 5.043741, 5.278961, 
    5.498487, 5.692443, 5.846371, 5.940264, 5.951795, 5.867255, 5.69812, 
    5.488389, 5.29539, 5.155908, 5.073154, 5.0311, 5.012152, 5.004404, 
    5.001488, 5.000471, 5.000139, 5.000038,
  // totalHeight(3,23, 0-49)
    5, 5, 5, 5, 5.000001, 5.000007, 5.000022, 5.00007, 5.000204, 5.000552, 
    5.001373, 5.003109, 5.006342, 5.011469, 5.017878, 30, 6.881858, 6.715767, 
    6.377157, 5.89924, 5.365091, 4.814788, 4.335211, 3.944315, 3.680533, 
    3.584269, 3.664799, 3.895799, 4.214448, 4.556406, 4.88979, 5.156824, 
    5.407378, 5.63265, 5.819686, 5.949622, 5.99874, 5.946925, 5.795018, 
    5.57985, 5.363815, 5.197576, 5.094623, 5.040833, 5.016148, 5.005916, 
    5.002019, 5.000645, 5.000192, 5.000054,
  // totalHeight(3,24, 0-49)
    5, 5, 5, 5, 5, 5.000004, 5.000014, 5.000044, 5.000131, 5.000354, 
    5.000885, 5.002009, 5.004103, 5.00741, 5.011444, 30, 6.913795, 6.743283, 
    6.393038, 5.88919, 5.313772, 4.708361, 4.169513, 3.717096, 3.405324, 
    3.291309, 3.388295, 3.663615, 4.035308, 4.421719, 4.790909, 5.082253, 
    5.354696, 5.599913, 5.805953, 5.955301, 6.024744, 5.991959, 5.852164, 
    5.636593, 5.40835, 5.225728, 5.109491, 5.047673, 5.018981, 5.006993, 
    5.0024, 5.000771, 5.00023, 5.000065,
  // totalHeight(3,25, 0-49)
    5, 5, 5, 5, 5.000001, 5.000007, 5.000023, 5.000068, 5.000196, 5.000519, 
    5.001256, 5.00277, 5.005505, 5.009689, 5.014659, 30, 6.917509, 6.746934, 
    6.394336, 5.883124, 5.294426, 4.670211, 4.109842, 3.634244, 3.304592, 
    3.184185, 3.287201, 3.579186, 3.97121, 4.374317, 4.756428, 5.056643, 
    5.336924, 5.589113, 5.801601, 5.957374, 6.033497, 6.007074, 5.871552, 
    5.656174, 5.423996, 5.235758, 5.114835, 5.050141, 5.020005, 5.007383, 
    5.002537, 5.000815, 5.000245, 5.000069,
  // totalHeight(3,26, 0-49)
    5, 5, 5, 5, 5.000005, 5.000018, 5.000054, 5.000162, 5.000451, 5.001157, 
    5.00272, 5.005827, 5.011258, 5.019319, 5.028754, 30, 6.889607, 6.723534, 
    6.378369, 5.879577, 5.308405, 4.705863, 4.168527, 3.716762, 3.405225, 
    3.291283, 3.388287, 3.663613, 4.035307, 4.421719, 4.790908, 5.082252, 
    5.354695, 5.599913, 5.805953, 5.955301, 6.024744, 5.991959, 5.852164, 
    5.636593, 5.40835, 5.225728, 5.109491, 5.047673, 5.018981, 5.006993, 
    5.0024, 5.000771, 5.00023, 5.000065,
  // totalHeight(3,27, 0-49)
    5, 5, 5, 5.000003, 5.000013, 5.000042, 5.000131, 5.000385, 5.001048, 
    5.002628, 5.006048, 5.012661, 5.02387, 5.039977, 5.058367, 30, 6.826754, 
    6.670672, 6.343395, 5.876875, 5.352436, 4.808751, 4.332749, 3.943442, 
    3.680258, 3.58419, 3.664778, 3.895793, 4.214446, 4.556406, 4.889789, 
    5.156823, 5.407378, 5.63265, 5.819686, 5.949621, 5.99874, 5.946925, 
    5.795018, 5.57985, 5.363815, 5.197576, 5.094623, 5.040833, 5.016148, 
    5.005916, 5.002019, 5.000645, 5.000192, 5.000054,
  // totalHeight(3,28, 0-49)
    5, 5, 5.000001, 5.000009, 5.000028, 5.000093, 5.000291, 5.000842, 
    5.002254, 5.005562, 5.012565, 5.025754, 5.047345, 5.076943, 5.108829, 30, 
    6.720564, 6.584433, 6.289873, 5.876649, 5.422355, 4.96215, 4.566208, 
    4.253551, 4.049467, 3.975818, 4.036649, 4.214753, 4.470621, 4.757757, 
    5.04374, 5.27896, 5.498487, 5.692443, 5.846371, 5.940264, 5.951794, 
    5.867256, 5.69812, 5.488389, 5.29539, 5.155908, 5.073154, 5.0311, 
    5.012152, 5.004404, 5.001488, 5.000471, 5.000139, 5.000038,
  // totalHeight(3,29, 0-49)
    5, 5, 5.000004, 5.000016, 5.000057, 5.000186, 5.000579, 5.001659, 
    5.004405, 5.010764, 5.024003, 5.048273, 5.086257, 5.134563, 5.180684, 30, 
    6.556565, 6.454806, 6.209808, 5.869759, 5.502885, 5.139183, 4.826483, 
    4.584808, 4.432256, 4.377896, 4.422847, 4.556728, 4.757828, 4.99201, 
    5.226871, 5.426193, 5.607547, 5.760535, 5.869822, 5.915688, 5.880161, 
    5.75981, 5.578391, 5.383534, 5.221547, 5.112823, 5.05154, 5.021459, 
    5.008235, 5.002935, 5.000975, 5.000303, 5.000089, 5.000024,
  // totalHeight(3,30, 0-49)
    5, 5.000002, 5.000008, 5.000027, 5.0001, 5.000338, 5.001072, 5.003178, 
    5.008781, 5.022519, 5.053143, 5.113769, 5.216212, 5.355342, 5.494076, 
    5.709598, 6.125762, 6.156536, 6.034242, 5.81732, 5.566053, 5.311934, 
    5.084235, 4.906974, 4.7975, 4.758753, 4.791675, 4.890025, 5.043805, 
    5.226883, 5.40879, 5.569041, 5.707834, 5.814003, 5.871604, 5.863268, 
    5.779329, 5.629799, 5.448622, 5.279824, 5.153577, 5.075142, 5.033274, 
    5.013503, 5.005065, 5.001767, 5.000576, 5.000175, 5.000051, 5.000014,
  // totalHeight(3,31, 0-49)
    5, 5.000001, 5.000006, 5.000023, 5.000086, 5.000294, 5.000936, 5.002785, 
    5.007725, 5.019886, 5.047167, 5.101953, 5.197631, 5.337241, 5.499212, 
    5.707389, 6.101362, 6.130861, 6.032712, 5.862597, 5.666519, 5.477023, 
    5.3025, 5.166655, 5.086007, 5.057975, 5.082697, 5.156963, 5.279002, 
    5.426205, 5.569045, 5.70021, 5.80257, 5.863031, 5.866385, 5.801664, 
    5.672307, 5.502812, 5.331985, 5.193449, 5.100338, 5.046923, 5.020027, 
    5.007874, 5.00287, 5.000974, 5.000309, 5.000092, 5.000025, 5.000007,
  // totalHeight(3,32, 0-49)
    5, 5, 5.000003, 5.000016, 5.000057, 5.000198, 5.000641, 5.001941, 
    5.005484, 5.014384, 5.034873, 5.077482, 5.155878, 5.27987, 5.442998, 
    5.649105, 5.993998, 6.054826, 6.009722, 5.902009, 5.764829, 5.636314, 
    5.511456, 5.412694, 5.356704, 5.337633, 5.354934, 5.407454, 5.49851, 
    5.607553, 5.707836, 5.802571, 5.86004, 5.867137, 5.813318, 5.698636, 
    5.540854, 5.372893, 5.228083, 5.124352, 5.061041, 5.027278, 5.011199, 
    5.004254, 5.001501, 5.000495, 5.000153, 5.000045, 5.000013, 5.000002,
  // totalHeight(3,33, 0-49)
    5, 5, 5.000001, 5.000009, 5.000031, 5.000113, 5.000374, 5.00116, 
    5.003356, 5.009038, 5.022561, 5.051877, 5.108922, 5.206487, 5.349631, 
    5.540675, 5.829793, 5.934906, 5.95664, 5.919773, 5.845279, 5.775891, 
    5.699202, 5.635369, 5.600927, 5.589468, 5.600031, 5.632689, 5.692454, 
    5.760539, 5.814003, 5.863031, 5.867137, 5.816883, 5.711125, 5.563231, 
    5.400769, 5.25464, 5.144711, 5.0741, 5.034512, 5.014745, 5.005819, 
    5.00213, 5.000726, 5.000232, 5.00007, 5.00002, 5.000005, 5,
  // totalHeight(3,34, 0-49)
    5, 5, 5, 5.000003, 5.000016, 5.000058, 5.000192, 5.000611, 5.001822, 
    5.00506, 5.013054, 5.031149, 5.068315, 5.13659, 5.246739, 5.405913, 
    5.637955, 5.777564, 5.862308, 5.896429, 5.887648, 5.877523, 5.849693, 
    5.821001, 5.806437, 5.801769, 5.806009, 5.819705, 5.846376, 5.869823, 
    5.871605, 5.866385, 5.813318, 5.711125, 5.5706, 5.414839, 5.271254, 
    5.159427, 5.084641, 5.040899, 5.018124, 5.00741, 5.002808, 5.000989, 
    5.000327, 5.000101, 5.00003, 5.000008, 5.000001, 5,
  // totalHeight(3,35, 0-49)
    5, 5, 5, 5.000001, 5.000007, 5.000026, 5.000089, 5.00029, 5.000893, 
    5.002561, 5.006839, 5.016948, 5.038792, 5.081545, 5.156356, 5.273779, 
    5.448004, 5.596495, 5.722991, 5.816328, 5.870923, 5.919303, 5.941797, 
    5.950219, 5.955517, 5.957448, 5.955325, 5.949628, 5.940266, 5.915689, 
    5.863268, 5.801664, 5.698636, 5.56323, 5.414839, 5.276899, 5.167127, 
    5.091476, 5.045663, 5.020916, 5.00884, 5.003462, 5.001259, 5.000427, 
    5.000136, 5.000041, 5.000012, 5.000003, 5, 5,
  // totalHeight(3,36, 0-49)
    5, 5, 5, 5, 5.000002, 5.000011, 5.000038, 5.000125, 5.000399, 5.001182, 
    5.00327, 5.008418, 5.020082, 5.044224, 5.089479, 5.166116, 5.285483, 
    5.41548, 5.55173, 5.678836, 5.782701, 5.881738, 5.952456, 5.998994, 
    6.024836, 6.033529, 6.024755, 5.998743, 5.951795, 5.880162, 5.77933, 
    5.672307, 5.540854, 5.400769, 5.271254, 5.167127, 5.093842, 5.048205, 
    5.022761, 5.009921, 5.004006, 5.001504, 5.000525, 5.000171, 5.000052, 
    5.000016, 5.000004, 5, 5, 5,
  // totalHeight(3,37, 0-49)
    5, 5, 5, 5, 5, 5.000004, 5.000015, 5.000051, 5.000163, 5.000501, 
    5.001435, 5.003837, 5.00953, 5.021924, 5.046564, 5.091146, 5.164802, 
    5.260377, 5.377213, 5.50543, 5.631152, 5.760442, 5.867519, 5.947026, 
    5.991995, 6.007086, 5.991962, 5.946927, 5.867255, 5.75981, 5.629799, 
    5.502812, 5.372893, 5.25464, 5.159427, 5.091476, 5.048205, 5.023404, 
    5.010503, 5.004369, 5.001688, 5.000608, 5.000204, 5.000064, 5.00002, 
    5.000005, 5, 5, 5, 5,
  // totalHeight(3,38, 0-49)
    5, 5, 5, 5, 5, 5, 5.000005, 5.00002, 5.000062, 5.000195, 5.00058, 
    5.001613, 5.004166, 5.009988, 5.022183, 5.045549, 5.086459, 5.146701, 
    5.229607, 5.33292, 5.449109, 5.578621, 5.698215, 5.795055, 5.852177, 
    5.871556, 5.852166, 5.79502, 5.69812, 5.578392, 5.448622, 5.331985, 
    5.228083, 5.144711, 5.084641, 5.045663, 5.022761, 5.010503, 5.004496, 
    5.001788, 5.000662, 5.000228, 5.000074, 5.000023, 5.000007, 5.000001, 5, 
    5, 5, 5,
  // totalHeight(3,39, 0-49)
    5, 5, 5, 5, 5, 5, 5.000001, 5.000007, 5.000022, 5.000071, 5.000218, 
    5.000627, 5.001684, 5.004201, 5.00973, 5.020876, 5.04146, 5.074723, 
    5.124831, 5.193744, 5.27998, 5.383608, 5.48842, 5.579863, 5.636596, 
    5.656175, 5.636593, 5.57985, 5.488389, 5.383535, 5.279824, 5.193449, 
    5.124352, 5.0741, 5.040899, 5.020916, 5.009921, 5.004369, 5.001788, 
    5.000681, 5.000242, 5.00008, 5.000025, 5.000008, 5.000002, 5, 5, 5, 5, 5,
  // totalHeight(3,40, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000008, 5.000024, 5.000075, 5.000226, 
    5.00063, 5.001637, 5.003948, 5.008826, 5.018284, 5.034691, 5.061178, 
    5.100423, 5.153621, 5.221567, 5.295398, 5.363819, 5.408352, 5.423996, 
    5.408351, 5.363815, 5.29539, 5.221547, 5.153577, 5.100338, 5.061041, 
    5.034512, 5.018124, 5.00884, 5.004006, 5.001688, 5.000662, 5.000242, 
    5.000082, 5.000026, 5.000008, 5.000002, 5, 5, 5, 5, 5, 5,
  // totalHeight(3,41, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000008, 5.000024, 5.000076, 5.00022, 
    5.000594, 5.001486, 5.003456, 5.007452, 5.014793, 5.027314, 5.046945, 
    5.075154, 5.112829, 5.15591, 5.197577, 5.225729, 5.235758, 5.225728, 
    5.197576, 5.155908, 5.112823, 5.075142, 5.046923, 5.027278, 5.014745, 
    5.00741, 5.003462, 5.001504, 5.000608, 5.000228, 5.00008, 5.000026, 
    5.000009, 5.000002, 5, 5, 5, 5, 5, 5, 5,
  // totalHeight(3,42, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000008, 5.000024, 5.000072, 
    5.0002, 5.000521, 5.001258, 5.002819, 5.00583, 5.011209, 5.020034, 
    5.033277, 5.051541, 5.073155, 5.094623, 5.109491, 5.114835, 5.109491, 
    5.094623, 5.073154, 5.05154, 5.033274, 5.020027, 5.011199, 5.005819, 
    5.002808, 5.001259, 5.000525, 5.000204, 5.000074, 5.000025, 5.000008, 
    5.000002, 5, 5, 5, 5, 5, 5, 5, 5,
  // totalHeight(3,43, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000008, 5.000023, 5.000063, 
    5.00017, 5.000428, 5.000993, 5.002134, 5.004256, 5.007876, 5.013503, 
    5.021459, 5.0311, 5.040833, 5.047673, 5.050141, 5.047673, 5.040833, 
    5.0311, 5.021459, 5.013503, 5.007874, 5.004254, 5.00213, 5.000989, 
    5.000427, 5.000171, 5.000064, 5.000023, 5.000008, 5.000002, 5, 5, 5, 5, 
    5, 5, 5, 5, 5,
  // totalHeight(3,44, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000007, 5.00002, 5.000052, 
    5.000136, 5.000328, 5.000727, 5.001502, 5.002871, 5.005065, 5.008235, 
    5.012152, 5.016148, 5.018981, 5.020005, 5.018981, 5.016148, 5.012152, 
    5.008235, 5.005065, 5.00287, 5.001501, 5.000726, 5.000327, 5.000136, 
    5.000052, 5.00002, 5.000007, 5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // totalHeight(3,45, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000005, 5.000016, 
    5.000041, 5.000101, 5.000232, 5.000495, 5.000975, 5.001767, 5.002935, 
    5.004404, 5.005916, 5.006993, 5.007383, 5.006993, 5.005916, 5.004404, 
    5.002935, 5.001767, 5.000974, 5.000495, 5.000232, 5.000101, 5.000041, 
    5.000016, 5.000005, 5.000001, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // totalHeight(3,46, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000004, 5.000012, 5.00003, 
    5.00007, 5.000153, 5.000309, 5.000576, 5.000975, 5.001488, 5.002019, 
    5.0024, 5.002537, 5.0024, 5.002019, 5.001488, 5.000975, 5.000576, 
    5.000309, 5.000153, 5.00007, 5.00003, 5.000012, 5.000004, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5,
  // totalHeight(3,47, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000003, 5.000008, 5.00002, 
    5.000045, 5.000092, 5.000175, 5.000303, 5.000471, 5.000645, 5.000771, 
    5.000815, 5.000771, 5.000645, 5.000471, 5.000303, 5.000175, 5.000092, 
    5.000045, 5.00002, 5.000008, 5.000003, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5,
  // totalHeight(3,48, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000005, 
    5.000013, 5.000025, 5.000051, 5.000089, 5.000139, 5.000192, 5.000231, 
    5.000245, 5.000231, 5.000192, 5.000139, 5.000089, 5.000051, 5.000025, 
    5.000013, 5.000005, 5.000001, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // totalHeight(3,49, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000006, 
    5.000012, 5.000023, 5.000038, 5.000055, 5.000067, 5.000071, 5.000067, 
    5.000055, 5.000038, 5.000023, 5.000012, 5.000006, 5.000002, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // totalHeight(4,0, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000006, 5.000013, 
    5.000028, 5.000057, 5.000112, 5.000206, 5.000354, 5.000569, 5.00085, 
    5.001171, 5.001479, 5.001697, 5.001776, 5.001697, 5.001479, 5.001171, 
    5.00085, 5.000569, 5.000354, 5.000206, 5.000112, 5.000057, 5.000028, 
    5.000013, 5.000006, 5.000001, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // totalHeight(4,1, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000003, 5.000008, 5.000018, 5.000039, 
    5.000082, 5.000166, 5.000319, 5.000575, 5.000974, 5.001544, 5.002285, 
    5.003127, 5.003933, 5.004504, 5.00471, 5.004504, 5.003933, 5.003127, 
    5.002285, 5.001544, 5.000974, 5.000575, 5.000319, 5.000166, 5.000082, 
    5.000038, 5.000018, 5.000008, 5.000003, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // totalHeight(4,2, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000004, 5.00001, 5.000022, 5.00005, 
    5.000111, 5.000235, 5.000467, 5.000876, 5.001545, 5.002564, 5.003994, 
    5.005826, 5.00789, 5.009855, 5.011244, 5.011746, 5.011244, 5.009855, 
    5.00789, 5.005825, 5.003993, 5.002563, 5.001543, 5.000874, 5.000466, 
    5.000235, 5.000111, 5.00005, 5.000022, 5.00001, 5.000004, 5, 5, 5, 5, 5, 
    5, 5, 5, 5,
  // totalHeight(4,3, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000005, 5.000011, 5.000026, 5.000062, 
    5.000142, 5.000312, 5.000645, 5.001252, 5.002286, 5.003933, 5.006382, 
    5.00975, 5.014007, 5.018755, 5.023253, 5.026416, 5.027557, 5.026416, 
    5.023252, 5.018755, 5.014006, 5.009748, 5.006378, 5.003928, 5.002279, 
    5.001247, 5.000645, 5.000314, 5.000144, 5.000063, 5.000027, 5.000011, 
    5.000005, 5.000001, 5, 5, 5, 5, 5, 5, 5,
  // totalHeight(4,4, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000005, 5.000012, 5.00003, 5.000073, 
    5.000174, 5.000391, 5.000835, 5.001678, 5.003172, 5.005635, 5.009448, 
    5.014966, 5.022386, 5.031617, 5.041789, 5.051358, 5.058033, 5.060435, 
    5.058033, 5.051356, 5.041786, 5.031611, 5.022377, 5.014951, 5.009429, 
    5.005613, 5.003155, 5.001675, 5.00084, 5.000397, 5.000178, 5.000076, 
    5.000031, 5.000013, 5.000005, 5.000001, 5, 5, 5, 5, 5, 5,
  // totalHeight(4,5, 0-49)
    5, 5, 5, 5, 5, 5, 5.000002, 5.000006, 5.000013, 5.000031, 5.000082, 
    5.0002, 5.000464, 5.00102, 5.002115, 5.004128, 5.00759, 5.013093, 
    5.021336, 5.032907, 5.048047, 5.066521, 5.086531, 5.105149, 5.117974, 
    5.122565, 5.117973, 5.105145, 5.086521, 5.066501, 5.048014, 5.032856, 
    5.021269, 5.01302, 5.007533, 5.004119, 5.002128, 5.001039, 5.00048, 
    5.00021, 5.000087, 5.000034, 5.000014, 5.000006, 5.000002, 5, 5, 5, 5, 5,
  // totalHeight(4,6, 0-49)
    5, 5, 5, 5, 5, 5.000001, 5.000006, 5.000013, 5.000033, 5.000086, 
    5.000218, 5.00052, 5.001176, 5.002513, 5.005054, 5.009583, 5.017104, 
    5.028571, 5.04509, 5.06742, 5.095617, 5.129127, 5.164507, 5.196824, 
    5.218638, 5.226384, 5.218632, 5.196807, 5.164472, 5.12906, 5.095507, 
    5.067253, 5.04487, 5.028332, 5.016919, 5.009551, 5.005095, 5.002568, 
    5.001224, 5.00055, 5.000236, 5.000094, 5.000036, 5.000015, 5.000007, 
    5.000002, 5, 5, 5, 5,
  // totalHeight(4,7, 0-49)
    5, 5, 5, 5, 5, 5.000005, 5.000013, 5.000032, 5.000086, 5.000224, 
    5.000552, 5.001284, 5.002817, 5.005834, 5.011383, 5.020915, 5.036179, 
    5.058282, 5.0886, 5.12762, 5.174555, 5.228317, 5.28298, 5.331494, 
    5.363276, 5.374424, 5.363256, 5.331442, 5.282871, 5.228115, 5.174216, 
    5.12711, 5.08793, 5.057558, 5.035612, 5.020813, 5.011489, 5.00599, 
    5.002948, 5.001372, 5.000603, 5.00025, 5.000099, 5.000037, 5.000015, 
    5.000006, 5.000001, 5, 5, 5,
  // totalHeight(4,8, 0-49)
    5, 5, 5, 5, 5.000004, 5.000011, 5.00003, 5.000083, 5.000219, 5.000553, 
    5.001321, 5.002983, 5.00635, 5.012745, 5.024074, 5.042771, 5.071508, 
    5.110453, 5.160557, 5.220954, 5.288945, 5.363122, 5.434719, 5.495795, 
    5.534249, 5.547521, 5.534192, 5.49565, 5.434417, 5.36256, 5.288007, 
    5.219527, 5.158675, 5.108407, 5.069887, 5.04248, 5.024346, 5.013159, 
    5.006711, 5.003231, 5.001469, 5.000631, 5.000257, 5.000099, 5.000036, 
    5.000014, 5.000005, 5.000001, 5, 5,
  // totalHeight(4,9, 0-49)
    5, 5, 5, 5.000003, 5.00001, 5.000027, 5.000073, 5.000201, 5.000522, 
    5.001283, 5.002978, 5.006522, 5.013456, 5.026117, 5.047627, 5.081541, 
    5.131313, 5.193063, 5.26604, 5.346703, 5.429886, 5.515448, 5.592755, 
    5.65555, 5.693194, 5.705945, 5.693052, 5.655185, 5.592003, 5.51405, 
    5.427536, 5.343099, 5.261235, 5.187773, 5.12704, 5.0808, 5.048308, 
    5.027168, 5.014386, 5.00718, 5.00338, 5.001504, 5.000631, 5.00025, 
    5.000094, 5.000034, 5.000013, 5.000005, 5, 5,
  // totalHeight(4,10, 0-49)
    5, 5, 5.000001, 5.000008, 5.000023, 5.000062, 5.000174, 5.000464, 
    5.001174, 5.002803, 5.006311, 5.01339, 5.026711, 5.050013, 5.087704, 
    5.143996, 5.222599, 5.309128, 5.400571, 5.490787, 5.573659, 5.653591, 
    5.720015, 5.770827, 5.799431, 5.808886, 5.799106, 5.770001, 5.718316, 
    5.65044, 5.568353, 5.482604, 5.389545, 5.296785, 5.212377, 5.142366, 
    5.089346, 5.052536, 5.028989, 5.015037, 5.007341, 5.00338, 5.001469, 
    5.000603, 5.000236, 5.000087, 5.000031, 5.000011, 5.000004, 5,
  // totalHeight(4,11, 0-49)
    5, 5.000001, 5.000006, 5.000018, 5.000051, 5.000142, 5.000389, 5.00101, 
    5.002481, 5.005745, 5.012537, 5.025723, 5.049498, 5.089058, 5.149407, 
    5.233919, 5.346392, 5.451672, 5.547588, 5.628493, 5.690985, 5.747229, 
    5.788034, 5.816257, 5.830287, 5.834641, 5.829595, 5.814518, 5.784492, 
    5.740716, 5.680092, 5.611754, 5.524933, 5.425946, 5.324495, 5.230956, 
    5.153233, 5.094786, 5.05476, 5.029618, 5.015037, 5.00718, 5.003231, 
    5.001372, 5.00055, 5.00021, 5.000076, 5.000027, 5.00001, 5.000003,
  // totalHeight(4,12, 0-49)
    5, 5.000003, 5.000013, 5.000038, 5.000109, 5.000305, 5.000814, 5.002055, 
    5.004901, 5.011015, 5.023273, 5.046094, 5.08526, 5.146695, 5.233996, 
    5.347453, 5.493467, 5.603019, 5.683767, 5.735504, 5.761001, 5.781113, 
    5.78789, 5.788424, 5.785759, 5.784305, 5.784378, 5.784986, 5.780982, 
    5.768596, 5.740397, 5.704315, 5.641876, 5.555245, 5.451858, 5.343374, 
    5.242486, 5.158862, 5.096653, 5.05476, 5.028989, 5.014386, 5.006711, 
    5.002948, 5.001224, 5.00048, 5.000178, 5.000063, 5.000022, 5.000008,
  // totalHeight(4,13, 0-49)
    5.000001, 5.000009, 5.000026, 5.000077, 5.000224, 5.000611, 5.001587, 
    5.003901, 5.009038, 5.019696, 5.040237, 5.07673, 5.135884, 5.222372, 
    5.33526, 5.470407, 5.644621, 5.740721, 5.789155, 5.798397, 5.778439, 
    5.757261, 5.727443, 5.699325, 5.679906, 5.672492, 5.677281, 5.692876, 
    5.71471, 5.734662, 5.742108, 5.744841, 5.718772, 5.661288, 5.574646, 
    5.467301, 5.352917, 5.246391, 5.158862, 5.094786, 5.052536, 5.027167, 
    5.013159, 5.00599, 5.002568, 5.001039, 5.000397, 5.000144, 5.00005, 
    5.000018,
  // totalHeight(4,14, 0-49)
    5.000004, 5.000016, 5.000051, 5.00015, 5.000423, 5.001134, 5.002876, 
    5.006879, 5.015491, 5.032723, 5.064547, 5.118182, 5.199555, 5.309104, 
    5.438466, 5.581018, 5.776528, 5.845946, 5.853991, 5.817026, 5.75099, 
    5.688416, 5.622475, 5.56643, 5.530651, 5.517122, 5.525881, 5.554883, 
    5.600159, 5.649828, 5.690797, 5.731436, 5.745387, 5.726641, 5.672071, 
    5.58408, 5.472425, 5.352917, 5.242486, 5.153233, 5.089346, 5.048308, 
    5.024346, 5.011489, 5.005095, 5.002128, 5.00084, 5.000314, 5.000111, 
    5.000039,
  // totalHeight(4,15, 0-49)
    5.000009, 5.00003, 5.000093, 5.000268, 5.000741, 5.001943, 5.004808, 
    5.011213, 5.02456, 5.050291, 5.095673, 5.167803, 5.269303, 5.393564, 
    5.523967, 5.657652, 5.868953, 5.907986, 5.878179, 5.799743, 5.692262, 
    5.590435, 5.489555, 5.406311, 5.354075, 5.333925, 5.345757, 5.386508, 
    5.452232, 5.527853, 5.598085, 5.67159, 5.722934, 5.744675, 5.730055, 
    5.67552, 5.58408, 5.467301, 5.343374, 5.230956, 5.142365, 5.080799, 
    5.04248, 5.020813, 5.009551, 5.004119, 5.001675, 5.000645, 5.000236, 
    5.000084,
  // totalHeight(4,16, 0-49)
    5.000016, 5.000051, 5.000154, 5.000436, 5.001185, 5.003041, 5.007361, 
    5.016769, 5.035784, 5.071095, 5.130445, 5.218989, 5.333667, 5.459665, 
    5.573878, 5.686548, 5.908281, 5.92311, 5.866307, 5.756901, 5.615705, 
    5.477578, 5.342819, 5.232497, 5.162915, 5.135132, 5.148944, 5.199866, 
    5.28306, 5.380913, 5.476108, 5.57633, 5.659531, 5.718256, 5.744269, 
    5.730054, 5.672071, 5.574646, 5.451857, 5.324495, 5.212377, 5.12704, 
    5.069887, 5.035612, 5.016918, 5.007533, 5.003155, 5.001247, 5.000467, 
    5.000169,
  // totalHeight(4,17, 0-49)
    5.000024, 5.000076, 5.000226, 5.000637, 5.0017, 5.004287, 5.01019, 
    5.022752, 5.047452, 5.091729, 5.162721, 5.26203, 5.379788, 5.493896, 
    5.577772, 5.66574, 5.886785, 5.890759, 5.822771, 5.696401, 5.531397, 
    5.360797, 5.193435, 5.055688, 4.967145, 4.93014, 4.944488, 5.003893, 
    5.101617, 5.218238, 5.334838, 5.456188, 5.56532, 5.655404, 5.718253, 
    5.744672, 5.726639, 5.661288, 5.555245, 5.425946, 5.296785, 5.187774, 
    5.108407, 5.057558, 5.028332, 5.01302, 5.005613, 5.00228, 5.000876, 
    5.000325,
  // totalHeight(4,18, 0-49)
    5.000031, 5.000098, 5.00029, 5.000809, 5.002132, 5.005311, 5.012467, 
    5.027443, 5.05629, 5.106589, 5.184099, 5.286392, 5.397364, 5.489583, 
    5.535452, 5.605662, 5.800894, 5.810308, 5.749249, 5.622153, 5.445377, 
    5.247847, 5.050285, 4.884759, 4.775092, 4.726635, 4.739514, 4.805339, 
    4.914531, 5.046517, 5.181646, 5.319603, 5.449533, 5.565309, 5.659521, 
    5.722928, 5.745382, 5.718771, 5.641876, 5.524933, 5.389545, 5.261234, 
    5.158674, 5.08793, 5.04487, 5.021269, 5.009429, 5.003929, 5.001545, 
    5.000584,
  // totalHeight(4,19, 0-49)
    5.000033, 5.000104, 5.000303, 5.000842, 5.002212, 5.00549, 5.012845, 
    5.02818, 5.057574, 5.108389, 5.185361, 5.283393, 5.381967, 5.449668, 
    5.45941, 5.528225, 5.651516, 5.679839, 5.644249, 5.534561, 5.360603, 
    5.14432, 4.920958, 4.727758, 4.594412, 4.531527, 4.540184, 4.609795, 
    4.727152, 4.870959, 5.022038, 5.172999, 5.319552, 5.45614, 5.576295, 
    5.67157, 5.731426, 5.744835, 5.704313, 5.611754, 5.482604, 5.343098, 
    5.219526, 5.12711, 5.067253, 5.032856, 5.014951, 5.00638, 5.002567, 
    5.000986,
  // totalHeight(4,20, 0-49)
    5.000022, 5.000071, 5.000206, 5.000566, 5.001461, 5.003547, 5.008075, 
    5.017149, 5.033758, 5.061057, 5.100434, 5.148736, 5.196876, 5.232886, 
    5.249486, 30, 5.72522, 5.722096, 5.663104, 5.536474, 5.342846, 5.092929, 
    4.832631, 4.601823, 4.436234, 4.352537, 4.352442, 4.422397, 4.544476, 
    4.696456, 4.860911, 5.021814, 5.181428, 5.334681, 5.476007, 5.598027, 
    5.690766, 5.742093, 5.74039, 5.680089, 5.568351, 5.427535, 5.288007, 
    5.174216, 5.095507, 5.048014, 5.022378, 5.00975, 5.003997, 5.001556,
  // totalHeight(4,21, 0-49)
    5.000014, 5.000044, 5.000126, 5.000348, 5.000903, 5.002204, 5.005051, 
    5.010816, 5.021541, 5.039646, 5.06693, 5.102845, 5.142964, 5.179457, 
    5.204838, 30, 5.693264, 5.683771, 5.624491, 5.49779, 5.296422, 5.020554, 
    4.725423, 4.45422, 4.252345, 4.146114, 4.139155, 4.214416, 4.347202, 
    4.512626, 4.695527, 4.870046, 5.045835, 5.217789, 5.380641, 5.527698, 
    5.649745, 5.734621, 5.768576, 5.740706, 5.650436, 5.514049, 5.36256, 
    5.228116, 5.12906, 5.066501, 5.031611, 5.014006, 5.005826, 5.002292,
  // totalHeight(4,22, 0-49)
    5.000008, 5.000024, 5.000072, 5.000199, 5.000521, 5.00129, 5.002997, 
    5.006517, 5.013214, 5.024857, 5.043125, 5.068581, 5.099402, 5.130821, 
    5.156437, 30, 5.645344, 5.631002, 5.571152, 5.445369, 5.241158, 4.948497, 
    4.63036, 4.328893, 4.096667, 3.969621, 3.954431, 4.03174, 4.170502, 
    4.343932, 4.540859, 4.72441, 4.91267, 5.100444, 5.282361, 5.451836, 
    5.599946, 5.7146, 5.780928, 5.784469, 5.718306, 5.591999, 5.434416, 
    5.28287, 5.164471, 5.086521, 5.041785, 5.018754, 5.007888, 5.003124,
  // totalHeight(4,23, 0-49)
    5.000003, 5.000014, 5.000041, 5.000118, 5.000312, 5.000783, 5.001848, 
    5.004087, 5.008446, 5.016229, 5.028857, 5.047226, 5.070715, 5.096325, 
    5.118713, 30, 5.596464, 5.578844, 5.518146, 5.392861, 5.187092, 4.88203, 
    4.546795, 4.220427, 3.96124, 3.815448, 3.794108, 3.875613, 4.021391, 
    4.202407, 4.412063, 4.602664, 4.800696, 5.001018, 5.198163, 5.385542, 
    5.554357, 5.692601, 5.784849, 5.814455, 5.769972, 5.655174, 5.495645, 
    5.33144, 5.196806, 5.105144, 5.051356, 5.023251, 5.009851, 5.003916,
  // totalHeight(4,24, 0-49)
    5.000002, 5.000011, 5.000033, 5.000093, 5.000248, 5.000626, 5.001483, 
    5.003294, 5.006839, 5.01322, 5.023686, 5.039129, 5.059257, 5.081702, 
    5.101663, 30, 5.556334, 5.537187, 5.476232, 5.351586, 5.145324, 4.83245, 
    4.485684, 4.140932, 3.860631, 3.700632, 3.676901, 3.765053, 3.9187, 
    4.106887, 4.327, 4.52336, 4.728728, 4.937836, 5.14499, 5.343493, 
    5.524635, 5.676622, 5.784046, 5.829436, 5.799034, 5.693022, 5.534179, 
    5.363252, 5.21863, 5.117971, 5.058032, 5.026413, 5.011236, 5.004478,
  // totalHeight(4,25, 0-49)
    5.000005, 5.000016, 5.000045, 5.000125, 5.000327, 5.000806, 5.00187, 
    5.004066, 5.00826, 5.015623, 5.027387, 5.044277, 5.06568, 5.088906, 
    5.109101, 30, 5.530094, 5.511153, 5.450953, 5.327627, 5.122614, 4.808633, 
    4.459426, 4.109352, 3.822037, 3.657288, 3.633398, 3.724782, 3.881723, 
    4.07268, 4.296721, 4.495244, 4.70334, 4.915673, 5.126443, 5.328887, 
    5.514308, 5.670983, 5.783531, 5.834264, 5.808712, 5.705871, 5.54749, 
    5.374413, 5.226382, 5.122564, 5.060434, 5.027554, 5.011736, 5.004682,
  // totalHeight(4,26, 0-49)
    5.00001, 5.00003, 5.000083, 5.000225, 5.000573, 5.001377, 5.003111, 
    5.006579, 5.012978, 5.023774, 5.040254, 5.062696, 5.089457, 5.116624, 
    5.138906, 30, 5.520136, 5.503262, 5.445169, 5.324215, 5.122498, 4.814704, 
    4.473166, 4.133136, 3.856438, 3.698707, 3.676142, 3.764788, 3.918613, 
    4.10686, 4.326991, 4.523357, 4.728727, 4.937836, 5.144989, 5.343493, 
    5.524634, 5.676622, 5.784046, 5.829436, 5.799034, 5.693022, 5.534179, 
    5.363252, 5.21863, 5.117971, 5.058032, 5.026413, 5.011236, 5.004478,
  // totalHeight(4,27, 0-49)
    5.000019, 5.000056, 5.000157, 5.000415, 5.001042, 5.002456, 5.005435, 
    5.011232, 5.021597, 5.038417, 5.062864, 5.094123, 5.128512, 5.160077, 
    5.183197, 30, 5.526995, 5.513671, 5.458173, 5.339542, 5.142099, 4.846486, 
    4.52138, 4.204391, 3.952483, 3.811342, 3.79244, 3.875007, 4.021184, 
    4.202338, 4.412041, 4.602656, 4.800694, 5.001017, 5.198163, 5.385541, 
    5.554357, 5.692601, 5.784849, 5.814455, 5.769972, 5.655174, 5.495645, 
    5.33144, 5.196806, 5.105144, 5.051356, 5.023251, 5.009851, 5.003916,
  // totalHeight(4,28, 0-49)
    5.000035, 5.0001, 5.000277, 5.000724, 5.001793, 5.004173, 5.009095, 
    5.018476, 5.034788, 5.060286, 5.095444, 5.137174, 5.178433, 5.210751, 
    5.229156, 30, 5.549765, 5.540964, 5.487337, 5.369511, 5.17579, 4.895623, 
    4.591888, 4.304254, 4.082989, 3.963053, 3.951664, 4.030686, 4.170128, 
    4.343802, 4.540814, 4.724395, 4.912664, 5.100442, 5.28236, 5.451836, 
    5.599946, 5.7146, 5.780928, 5.784469, 5.718305, 5.591999, 5.434416, 
    5.28287, 5.164471, 5.086521, 5.041785, 5.018754, 5.007888, 5.003124,
  // totalHeight(4,29, 0-49)
    5.000054, 5.000159, 5.000442, 5.001153, 5.00284, 5.006568, 5.014205, 
    5.028555, 5.05294, 5.08968, 5.137436, 5.189026, 5.232651, 5.257787, 
    5.262488, 30, 5.584862, 5.579939, 5.525392, 5.405305, 5.214372, 4.952533, 
    4.675216, 4.421723, 4.234072, 4.137152, 4.135252, 4.212865, 4.346626, 
    4.51242, 4.695455, 4.870021, 5.045825, 5.217786, 5.380639, 5.527698, 
    5.649745, 5.734621, 5.768576, 5.740706, 5.650436, 5.514049, 5.36256, 
    5.228116, 5.12906, 5.066501, 5.031611, 5.014006, 5.005826, 5.002292,
  // totalHeight(4,30, 0-49)
    5.000076, 5.000227, 5.000637, 5.001688, 5.004233, 5.010009, 5.022226, 
    5.046075, 5.08837, 5.154881, 5.244466, 5.342824, 5.423133, 5.457164, 
    5.429102, 5.460217, 5.513269, 5.527208, 5.492916, 5.390181, 5.221525, 
    4.998848, 4.766492, 4.560466, 4.413423, 4.341393, 4.347546, 4.42042, 
    4.543725, 4.696185, 4.860814, 5.02178, 5.181416, 5.334677, 5.476006, 
    5.598026, 5.690766, 5.742093, 5.74039, 5.680089, 5.568351, 5.427535, 
    5.288007, 5.174216, 5.095507, 5.048014, 5.022378, 5.00975, 5.003997, 
    5.001556,
  // totalHeight(4,31, 0-49)
    5.000073, 5.000221, 5.000621, 5.001653, 5.00416, 5.009876, 5.02202, 
    5.045835, 5.088351, 5.155962, 5.249051, 5.356033, 5.453192, 5.513427, 
    5.51753, 5.549628, 5.688647, 5.683352, 5.618227, 5.4899, 5.309708, 
    5.098572, 4.885837, 4.704521, 4.580997, 4.524658, 4.537004, 4.608436, 
    4.726605, 4.870749, 5.021959, 5.17297, 5.319542, 5.456137, 5.576294, 
    5.671569, 5.731426, 5.744835, 5.704313, 5.611754, 5.482604, 5.343098, 
    5.219526, 5.12711, 5.067253, 5.032856, 5.014951, 5.00638, 5.002567, 
    5.000986,
  // totalHeight(4,32, 0-49)
    5.000058, 5.000175, 5.000499, 5.001343, 5.003422, 5.008226, 5.018595, 
    5.039321, 5.077241, 5.13961, 5.229686, 5.340741, 5.453701, 5.542929, 
    5.586711, 5.634364, 5.810377, 5.794869, 5.715106, 5.578702, 5.402011, 
    5.211908, 5.024439, 4.868459, 4.765963, 4.722025, 4.737376, 4.804413, 
    4.91415, 5.046367, 5.181589, 5.319583, 5.449525, 5.565306, 5.65952, 
    5.722928, 5.745382, 5.718771, 5.641876, 5.524932, 5.389545, 5.261234, 
    5.158674, 5.08793, 5.04487, 5.021269, 5.009429, 5.003929, 5.001545, 
    5.000584,
  // totalHeight(4,33, 0-49)
    5.00004, 5.000121, 5.000348, 5.000955, 5.002475, 5.006059, 5.013967, 
    5.030193, 5.060858, 5.113483, 5.193935, 5.30105, 5.422253, 5.535433, 
    5.617548, 5.69124, 5.875936, 5.864213, 5.786301, 5.657351, 5.496267, 
    5.333714, 5.17509, 5.044634, 4.961142, 4.927159, 4.943112, 5.003295, 
    5.101369, 5.218139, 5.334802, 5.456174, 5.565315, 5.655402, 5.718253, 
    5.744672, 5.726639, 5.661288, 5.555245, 5.425946, 5.296785, 5.187774, 
    5.108407, 5.057558, 5.028332, 5.01302, 5.005613, 5.00228, 5.000876, 
    5.000325,
  // totalHeight(4,34, 0-49)
    5.000024, 5.000075, 5.000218, 5.000609, 5.001614, 5.004035, 5.009521, 
    5.021117, 5.043819, 5.084566, 5.150602, 5.245469, 5.363938, 5.490148, 
    5.602442, 5.704795, 5.886364, 5.892461, 5.832005, 5.724312, 5.588806, 
    5.458125, 5.330325, 5.225271, 5.159105, 5.133275, 5.148096, 5.1995, 
    5.282907, 5.380851, 5.476084, 5.576321, 5.659528, 5.718254, 5.744268, 
    5.730054, 5.672071, 5.574646, 5.451857, 5.324495, 5.212377, 5.12704, 
    5.069887, 5.035612, 5.016918, 5.007533, 5.003155, 5.001247, 5.000467, 
    5.000169,
  // totalHeight(4,35, 0-49)
    5.000014, 5.000041, 5.000124, 5.000355, 5.000961, 5.002462, 5.00596, 
    5.013583, 5.029061, 5.058093, 5.107836, 5.184575, 5.289448, 5.414499, 
    5.54309, 5.668658, 5.844255, 5.878744, 5.849082, 5.774486, 5.672875, 
    5.577171, 5.48142, 5.401774, 5.351748, 5.332812, 5.345255, 5.386293, 
    5.452143, 5.527818, 5.598071, 5.671585, 5.722932, 5.744674, 5.730054, 
    5.67552, 5.58408, 5.467301, 5.343374, 5.230956, 5.142365, 5.080799, 
    5.04248, 5.020813, 5.009551, 5.004119, 5.001675, 5.000645, 5.000236, 
    5.000084,
  // totalHeight(4,36, 0-49)
    5.000007, 5.000022, 5.000065, 5.00019, 5.000528, 5.001387, 5.003449, 
    5.008088, 5.01785, 5.036942, 5.071377, 5.128031, 5.211954, 5.322424, 
    5.450345, 5.586574, 5.754741, 5.821698, 5.831575, 5.79887, 5.73787, 
    5.679853, 5.617424, 5.563701, 5.529284, 5.51648, 5.525597, 5.554762, 
    5.600111, 5.649807, 5.69079, 5.731433, 5.745385, 5.72664, 5.672071, 
    5.58408, 5.472425, 5.352917, 5.242486, 5.153233, 5.089346, 5.048308, 
    5.024346, 5.011489, 5.005095, 5.002128, 5.00084, 5.000314, 5.000111, 
    5.000039,
  // totalHeight(4,37, 0-49)
    5.000002, 5.000011, 5.000032, 5.000094, 5.00027, 5.000727, 5.001855, 
    5.004479, 5.010196, 5.021828, 5.043808, 5.082083, 5.142909, 5.230166, 
    5.342067, 5.472644, 5.628459, 5.722989, 5.773468, 5.786318, 5.77012, 
    5.752038, 5.724462, 5.697757, 5.679138, 5.672138, 5.677126, 5.692811, 
    5.714684, 5.734652, 5.742105, 5.744839, 5.718772, 5.661288, 5.574646, 
    5.467301, 5.352917, 5.246391, 5.158862, 5.094786, 5.052536, 5.027167, 
    5.013159, 5.00599, 5.002568, 5.001039, 5.000397, 5.000144, 5.00005, 
    5.000018,
  // totalHeight(4,38, 0-49)
    5, 5.000005, 5.000015, 5.000044, 5.000129, 5.000355, 5.000931, 5.002315, 
    5.005435, 5.012023, 5.025013, 5.048794, 5.088931, 5.150884, 5.237588, 
    5.348084, 5.483159, 5.591568, 5.673834, 5.728097, 5.756079, 5.778114, 
    5.786222, 5.787565, 5.785347, 5.784119, 5.784297, 5.784952, 5.780969, 
    5.768591, 5.740396, 5.704315, 5.641877, 5.555245, 5.451857, 5.343374, 
    5.242486, 5.158862, 5.096653, 5.05476, 5.028989, 5.014386, 5.006711, 
    5.002948, 5.001224, 5.00048, 5.000178, 5.000063, 5.000022, 5.000008,
  // totalHeight(4,39, 0-49)
    5, 5.000001, 5.000007, 5.00002, 5.000057, 5.000163, 5.000438, 5.00112, 
    5.002711, 5.006193, 5.013331, 5.026992, 5.051274, 5.091135, 5.151162, 
    5.233976, 5.340683, 5.445152, 5.541938, 5.624341, 5.688284, 5.745618, 
    5.787155, 5.815814, 5.830077, 5.834549, 5.829556, 5.814503, 5.784487, 
    5.740712, 5.680091, 5.611754, 5.524933, 5.425946, 5.324495, 5.230956, 
    5.153233, 5.094786, 5.05476, 5.029618, 5.015037, 5.00718, 5.003231, 
    5.001372, 5.00055, 5.00021, 5.000076, 5.000027, 5.00001, 5.000003,
  // totalHeight(4,40, 0-49)
    5, 5, 5.000002, 5.000009, 5.000025, 5.00007, 5.000193, 5.000509, 
    5.001269, 5.002991, 5.006652, 5.013947, 5.027512, 5.050968, 5.088504, 
    5.143935, 5.219826, 5.305856, 5.397701, 5.488678, 5.572298, 5.652788, 
    5.719582, 5.770612, 5.799332, 5.808841, 5.799087, 5.769994, 5.718313, 
    5.650439, 5.568352, 5.482605, 5.389545, 5.296785, 5.212377, 5.142365, 
    5.089346, 5.052536, 5.028989, 5.015037, 5.007341, 5.00338, 5.001469, 
    5.000603, 5.000236, 5.000087, 5.000031, 5.000011, 5.000004, 5,
  // totalHeight(4,41, 0-49)
    5, 5, 5, 5.000003, 5.000011, 5.000029, 5.000081, 5.000217, 5.000558, 
    5.001357, 5.003117, 5.006752, 5.013795, 5.026531, 5.047973, 5.081492, 
    5.130116, 5.191607, 5.264742, 5.345742, 5.429265, 5.515083, 5.592558, 
    5.655453, 5.693151, 5.705927, 5.693044, 5.655183, 5.592001, 5.51405, 
    5.427535, 5.343099, 5.261235, 5.187774, 5.12704, 5.080799, 5.048308, 
    5.027167, 5.014386, 5.00718, 5.00338, 5.001504, 5.000631, 5.00025, 
    5.000094, 5.000034, 5.000013, 5.000005, 5, 5,
  // totalHeight(4,42, 0-49)
    5, 5, 5, 5, 5.000005, 5.000012, 5.000032, 5.000088, 5.000232, 5.00058, 
    5.001373, 5.003073, 5.006487, 5.012912, 5.024214, 5.042749, 5.071041, 
    5.10987, 5.16003, 5.220561, 5.28869, 5.362971, 5.434639, 5.495757, 
    5.534231, 5.547513, 5.534188, 5.495649, 5.434417, 5.36256, 5.288007, 
    5.219526, 5.158674, 5.108407, 5.069887, 5.04248, 5.024346, 5.013159, 
    5.006711, 5.003231, 5.001469, 5.000631, 5.000257, 5.000099, 5.000036, 
    5.000014, 5.000005, 5.000001, 5, 5,
  // totalHeight(4,43, 0-49)
    5, 5, 5, 5, 5.000001, 5.000005, 5.000013, 5.000034, 5.000092, 5.000234, 
    5.000571, 5.001317, 5.002868, 5.005898, 5.011437, 5.020907, 5.036011, 
    5.058069, 5.088407, 5.127475, 5.17446, 5.228262, 5.28295, 5.331479, 
    5.36327, 5.374421, 5.363255, 5.331441, 5.28287, 5.228115, 5.174216, 
    5.12711, 5.08793, 5.057558, 5.035612, 5.020813, 5.011489, 5.00599, 
    5.002948, 5.001372, 5.000603, 5.00025, 5.000099, 5.000037, 5.000015, 
    5.000006, 5.000001, 5, 5, 5,
  // totalHeight(4,44, 0-49)
    5, 5, 5, 5, 5, 5.000001, 5.000006, 5.000014, 5.000034, 5.00009, 5.000225, 
    5.000533, 5.001195, 5.002535, 5.005076, 5.009581, 5.017048, 5.028498, 
    5.045024, 5.067372, 5.095585, 5.129107, 5.164498, 5.196819, 5.218636, 
    5.226383, 5.218631, 5.196807, 5.164472, 5.12906, 5.095506, 5.067253, 
    5.044869, 5.028332, 5.016918, 5.009551, 5.005095, 5.002568, 5.001224, 
    5.00055, 5.000236, 5.000094, 5.000036, 5.000015, 5.000007, 5.000002, 5, 
    5, 5, 5,
  // totalHeight(4,45, 0-49)
    5, 5, 5, 5, 5, 5, 5.000002, 5.000006, 5.000013, 5.000032, 5.000083, 
    5.000204, 5.000471, 5.001028, 5.002122, 5.004128, 5.007573, 5.013069, 
    5.021315, 5.032892, 5.048037, 5.066514, 5.086528, 5.105148, 5.117975, 
    5.122566, 5.117973, 5.105145, 5.086521, 5.0665, 5.048013, 5.032856, 
    5.021268, 5.013019, 5.007533, 5.004119, 5.002128, 5.001039, 5.00048, 
    5.00021, 5.000087, 5.000034, 5.000014, 5.000006, 5.000002, 5, 5, 5, 5, 5,
  // totalHeight(4,46, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000005, 5.000012, 5.00003, 5.000074, 
    5.000175, 5.000395, 5.000838, 5.001678, 5.003167, 5.005628, 5.009441, 
    5.01496, 5.022381, 5.031613, 5.041788, 5.051359, 5.058036, 5.060439, 
    5.058036, 5.051358, 5.041786, 5.03161, 5.022376, 5.014949, 5.009427, 
    5.005613, 5.003155, 5.001675, 5.00084, 5.000397, 5.000178, 5.000076, 
    5.000031, 5.000013, 5.000005, 5.000001, 5, 5, 5, 5, 5, 5,
  // totalHeight(4,47, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000005, 5.000011, 5.000026, 5.000062, 
    5.000143, 5.000313, 5.000644, 5.001248, 5.002281, 5.003928, 5.006376, 
    5.009744, 5.014003, 5.018755, 5.023259, 5.026426, 5.027568, 5.026426, 
    5.023259, 5.018755, 5.014002, 5.009743, 5.006373, 5.003924, 5.002277, 
    5.001245, 5.000643, 5.000314, 5.000143, 5.000063, 5.000027, 5.000011, 
    5.000005, 5.000001, 5, 5, 5, 5, 5, 5, 5,
  // totalHeight(4,48, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000004, 5.00001, 5.000022, 5.000049, 
    5.000109, 5.000232, 5.000462, 5.000867, 5.001534, 5.002549, 5.003979, 
    5.005815, 5.007891, 5.009873, 5.011274, 5.01178, 5.011274, 5.009873, 
    5.007891, 5.005815, 5.003978, 5.002548, 5.001532, 5.000866, 5.000462, 
    5.000232, 5.000109, 5.000049, 5.000022, 5.00001, 5.000004, 5, 5, 5, 5, 5, 
    5, 5, 5, 5,
  // totalHeight(4,49, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000005, 5.000012, 5.00003, 
    5.000065, 5.000139, 5.000275, 5.000512, 5.000896, 5.001465, 5.002233, 
    5.00314, 5.004033, 5.004668, 5.004897, 5.004668, 5.004033, 5.00314, 
    5.002233, 5.001465, 5.000896, 5.000512, 5.000275, 5.000139, 5.000065, 
    5.00003, 5.000012, 5.000005, 5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // totalHeight(5,0, 0-49)
    5, 5, 5, 5, 5, 5, 5.000002, 5.000006, 5.000013, 5.000028, 5.000061, 
    5.00013, 5.000265, 5.000516, 5.00096, 5.001699, 5.002862, 5.004584, 
    5.006996, 5.010178, 5.014109, 5.018611, 5.023259, 5.027408, 5.030265, 
    5.031285, 5.030264, 5.027405, 5.023253, 5.018603, 5.014096, 5.010162, 
    5.006977, 5.004565, 5.002849, 5.001694, 5.000961, 5.00052, 5.000268, 
    5.000132, 5.000062, 5.000028, 5.000013, 5.000006, 5.000002, 5, 5, 5, 5, 5,
  // totalHeight(5,1, 0-49)
    5, 5, 5, 5, 5, 5.000004, 5.000008, 5.000015, 5.000031, 5.000068, 
    5.000149, 5.000312, 5.000626, 5.0012, 5.002189, 5.003802, 5.006291, 
    5.0099, 5.01486, 5.021302, 5.029162, 5.038113, 5.047316, 5.055529, 
    5.06116, 5.063167, 5.061155, 5.05552, 5.047298, 5.038086, 5.029122, 
    5.021251, 5.0148, 5.00984, 5.006246, 5.003785, 5.002189, 5.001209, 
    5.000637, 5.00032, 5.000154, 5.000071, 5.000032, 5.000015, 5.000008, 
    5.000004, 5, 5, 5, 5,
  // totalHeight(5,2, 0-49)
    5, 5, 5, 5, 5.000005, 5.000009, 5.000016, 5.000033, 5.000074, 5.000168, 
    5.000363, 5.000746, 5.001466, 5.00274, 5.004883, 5.00829, 5.013408, 
    5.020618, 5.030261, 5.042474, 5.057049, 5.073393, 5.08998, 5.104668, 
    5.114639, 5.118178, 5.114626, 5.10464, 5.089929, 5.07331, 5.056931, 
    5.042319, 5.030082, 5.020443, 5.013276, 5.008237, 5.00488, 5.002761, 
    5.001492, 5.000769, 5.000379, 5.000178, 5.000082, 5.000035, 5.000017, 
    5.000009, 5.000005, 5.000001, 5, 5,
  // totalHeight(5,3, 0-49)
    5, 5, 5, 5.000004, 5.000009, 5.000016, 5.000034, 5.000081, 5.000184, 
    5.000405, 5.000853, 5.001713, 5.00328, 5.005985, 5.010404, 5.017234, 
    5.027194, 5.040734, 5.058229, 5.079662, 5.104465, 5.131642, 5.158663, 
    5.182254, 5.198014, 5.203566, 5.197978, 5.182171, 5.158515, 5.131409, 
    5.104133, 5.079228, 5.057729, 5.040246, 5.026826, 5.017087, 5.010396, 
    5.006039, 5.00335, 5.001772, 5.000896, 5.000432, 5.000201, 5.000089, 
    5.000038, 5.000018, 5.00001, 5.000006, 5.000001, 5,
  // totalHeight(5,4, 0-49)
    5, 5, 5.000002, 5.000008, 5.000016, 5.000034, 5.000082, 5.000193, 
    5.000432, 5.000931, 5.001913, 5.003746, 5.006992, 5.012434, 5.021055, 
    5.033954, 5.052146, 5.075799, 5.105033, 5.139303, 5.177319, 5.217662, 
    5.25659, 5.289864, 5.311574, 5.319134, 5.311477, 5.289647, 5.256206, 
    5.217056, 5.176451, 5.13817, 5.103726, 5.074522, 5.051179, 5.033571, 
    5.021023, 5.012565, 5.007167, 5.003901, 5.002026, 5.001004, 5.000476, 
    5.000216, 5.000093, 5.00004, 5.000018, 5.00001, 5.000005, 5,
  // totalHeight(5,5, 0-49)
    5, 5.000001, 5.000006, 5.000015, 5.000033, 5.000081, 5.000193, 5.000442, 
    5.000971, 5.002039, 5.004083, 5.00779, 5.014157, 5.024488, 5.040304, 
    5.063102, 5.094024, 5.131987, 5.176251, 5.225178, 5.276432, 5.328592, 
    5.376917, 5.417064, 5.442416, 5.451099, 5.442188, 5.416547, 5.376002, 
    5.32715, 5.274362, 5.222458, 5.173093, 5.128881, 5.09165, 5.062176, 
    5.040218, 5.024799, 5.014578, 5.008171, 5.004367, 5.002228, 5.001084, 
    5.000504, 5.000224, 5.000095, 5.00004, 5.000018, 5.000009, 5.000004,
  // totalHeight(5,6, 0-49)
    5.000001, 5.000005, 5.000013, 5.000031, 5.000074, 5.000183, 5.00043, 
    5.000967, 5.002075, 5.004246, 5.008282, 5.015374, 5.02715, 5.045572, 
    5.072659, 5.110019, 5.15846, 5.213607, 5.273174, 5.334088, 5.393208, 
    5.450352, 5.500582, 5.540859, 5.565177, 5.573293, 5.564681, 5.539737, 
    5.498604, 5.447233, 5.388718, 5.328151, 5.266213, 5.206674, 5.153087, 
    5.107989, 5.072482, 5.046282, 5.028121, 5.016266, 5.008961, 5.004705, 
    5.002356, 5.001125, 5.000514, 5.000224, 5.000093, 5.000038, 5.000018, 
    5.000008,
  // totalHeight(5,7, 0-49)
    5.000004, 5.00001, 5.000028, 5.000067, 5.000166, 5.0004, 5.000918, 
    5.002015, 5.004214, 5.008401, 5.015932, 5.02872, 5.04916, 5.079797, 
    5.122718, 5.178854, 5.248075, 5.319426, 5.389174, 5.453479, 5.509659, 
    5.560696, 5.602446, 5.634424, 5.65239, 5.658066, 5.651396, 5.632189, 
    5.598525, 5.554535, 5.500804, 5.441733, 5.375283, 5.305392, 5.237004, 
    5.174875, 5.122472, 5.081369, 5.051301, 5.030718, 5.017484, 5.009469, 
    5.004883, 5.002399, 5.001125, 5.000504, 5.000216, 5.000089, 5.000036, 
    5.000016,
  // totalHeight(5,8, 0-49)
    5.000009, 5.000022, 5.000058, 5.000145, 5.000354, 5.000831, 5.001863, 
    5.003988, 5.008126, 5.015749, 5.028997, 5.050632, 5.083705, 5.130813, 
    5.193053, 5.269456, 5.35902, 5.440007, 5.509358, 5.56441, 5.604834, 
    5.638444, 5.662354, 5.67907, 5.686673, 5.688493, 5.684813, 5.674917, 
    5.655134, 5.627209, 5.588828, 5.543271, 5.484299, 5.414421, 5.338465, 
    5.262632, 5.193025, 5.134175, 5.088205, 5.054886, 5.03237, 5.018123, 
    5.009644, 5.004883, 5.002356, 5.001084, 5.000476, 5.000201, 5.000082, 
    5.000034,
  // totalHeight(5,9, 0-49)
    5.000019, 5.000048, 5.00012, 5.000298, 5.000716, 5.001643, 5.003593, 
    5.007489, 5.014842, 5.027926, 5.049793, 5.083932, 5.133445, 5.199761, 
    5.281408, 5.374544, 5.47942, 5.558947, 5.615193, 5.648915, 5.663444, 
    5.671911, 5.672351, 5.669973, 5.665254, 5.662431, 5.661954, 5.662679, 
    5.659845, 5.652761, 5.636622, 5.613993, 5.574114, 5.516903, 5.445178, 
    5.364569, 5.282547, 5.20661, 5.142382, 5.092508, 5.056751, 5.032938, 
    5.018123, 5.009469, 5.004705, 5.002228, 5.001004, 5.000433, 5.00018, 
    5.000075,
  // totalHeight(5,10, 0-49)
    5.000036, 5.000093, 5.000239, 5.000585, 5.001373, 5.003076, 5.006561, 
    5.013308, 5.02562, 5.046711, 5.08042, 5.130344, 5.198357, 5.283011, 
    5.378876, 5.479668, 5.591911, 5.658225, 5.691349, 5.696425, 5.68037, 
    5.66087, 5.636159, 5.613672, 5.596256, 5.58842, 5.590661, 5.601462, 
    5.615591, 5.630049, 5.638243, 5.642887, 5.629557, 5.59555, 5.540604, 
    5.467718, 5.383308, 5.296116, 5.215004, 5.146606, 5.093976, 5.056751, 
    5.03237, 5.017484, 5.008961, 5.004367, 5.002027, 5.000896, 5.000381, 
    5.000162,
  // totalHeight(5,11, 0-49)
    5.000071, 5.000181, 5.000453, 5.001088, 5.002494, 5.005449, 5.011323, 
    5.022336, 5.041712, 5.073508, 5.121789, 5.189017, 5.274099, 5.371275, 
    5.471056, 5.567159, 5.679311, 5.724144, 5.729917, 5.705225, 5.659316, 
    5.612999, 5.564149, 5.522204, 5.492456, 5.479336, 5.483345, 5.502607, 
    5.531834, 5.56584, 5.596796, 5.628322, 5.64375, 5.638568, 5.609673, 
    5.556548, 5.482425, 5.39456, 5.302978, 5.217842, 5.146606, 5.092508, 
    5.054886, 5.030718, 5.016266, 5.008171, 5.003901, 5.001774, 5.000774, 
    5.000335,
  // totalHeight(5,12, 0-49)
    5.000131, 5.00033, 5.000812, 5.001908, 5.004274, 5.00911, 5.018438, 
    5.035336, 5.0639, 5.108568, 5.172517, 5.255433, 5.351807, 5.45142, 
    5.54234, 5.622025, 5.729712, 5.750149, 5.730207, 5.67971, 5.608513, 
    5.538956, 5.468381, 5.40834, 5.366759, 5.347938, 5.352461, 5.37809, 
    5.419709, 5.470071, 5.520361, 5.575464, 5.617815, 5.642097, 5.643387, 
    5.618141, 5.565696, 5.48967, 5.398307, 5.302978, 5.215004, 5.142382, 
    5.088205, 5.051301, 5.028121, 5.014579, 5.007169, 5.003353, 5.001502, 
    5.000663,
  // totalHeight(5,13, 0-49)
    5.000229, 5.000569, 5.001369, 5.00315, 5.006894, 5.014339, 5.02826, 
    5.052577, 5.091915, 5.1502, 5.228284, 5.321659, 5.420121, 5.510469, 
    5.580884, 5.636158, 5.738116, 5.735927, 5.695858, 5.626519, 5.536742, 
    5.448798, 5.359662, 5.283228, 5.230228, 5.205044, 5.208557, 5.238231, 
    5.289241, 5.352497, 5.418259, 5.492509, 5.55786, 5.608896, 5.639956, 
    5.645646, 5.622089, 5.568675, 5.48967, 5.39456, 5.296116, 5.20661, 
    5.134175, 5.081369, 5.046282, 5.0248, 5.012568, 5.006046, 5.00278, 
    5.001256,
  // totalHeight(5,14, 0-49)
    5.000374, 5.000917, 5.002163, 5.004873, 5.010436, 5.021191, 5.040668, 
    5.073408, 5.123923, 5.194474, 5.282308, 5.378265, 5.468612, 5.539557, 
    5.581494, 5.609149, 5.704862, 5.684734, 5.631863, 5.551764, 5.45104, 
    5.350298, 5.246478, 5.15581, 5.091814, 5.059381, 5.060057, 5.091223, 
    5.148467, 5.22124, 5.298869, 5.387869, 5.471773, 5.545377, 5.60301, 
    5.638582, 5.646293, 5.622088, 5.565695, 5.482424, 5.383307, 5.282547, 
    5.193025, 5.122472, 5.072483, 5.040219, 5.021027, 5.010407, 5.004912, 
    5.002266,
  // totalHeight(5,15, 0-49)
    5.000567, 5.001374, 5.003187, 5.00704, 5.014763, 5.029299, 5.054786, 
    5.09597, 5.156433, 5.235746, 5.326997, 5.417121, 5.49086, 5.535902, 
    5.545708, 5.546775, 5.632914, 5.60088, 5.542744, 5.459904, 5.356049, 
    5.248635, 5.134977, 5.033073, 4.95883, 4.918158, 4.913803, 4.943549, 
    5.003622, 5.082602, 5.168946, 5.268797, 5.367137, 5.458964, 5.538911, 
    5.600954, 5.638575, 5.645641, 5.618137, 5.556546, 5.467716, 5.364568, 
    5.262632, 5.174875, 5.10799, 5.062179, 5.033578, 5.017106, 5.008286, 
    5.003901,
  // totalHeight(5,16, 0-49)
    5.000793, 5.001904, 5.004345, 5.009432, 5.01941, 5.037717, 5.06884, 
    5.117216, 5.184804, 5.268004, 5.356136, 5.433732, 5.48586, 5.502688, 
    5.480472, 5.459173, 5.525829, 5.488203, 5.431913, 5.353796, 5.254422, 
    5.146871, 5.029435, 4.92056, 4.837578, 4.787774, 4.775797, 4.80067, 
    4.859735, 4.941498, 5.033751, 5.14112, 5.250391, 5.356567, 5.454606, 
    5.538887, 5.602984, 5.639937, 5.643376, 5.609665, 5.5406, 5.445177, 
    5.338465, 5.237003, 5.153089, 5.091654, 5.05119, 5.026856, 5.013346, 
    5.006411,
  // totalHeight(5,17, 0-49)
    5.001009, 5.002405, 5.005424, 5.01161, 5.023516, 5.044888, 5.080247, 
    5.133332, 5.204224, 5.28643, 5.36658, 5.428285, 5.457914, 5.448078, 
    5.397178, 5.359798, 5.38727, 5.349489, 5.301646, 5.235264, 5.147697, 
    5.046798, 4.932895, 4.822896, 4.733915, 4.674499, 4.651908, 4.667727, 
    4.721311, 4.802092, 4.897588, 5.009571, 5.126815, 5.244068, 5.35647, 
    5.458864, 5.5453, 5.608845, 5.642067, 5.638551, 5.595541, 5.5169, 
    5.414419, 5.305392, 5.206675, 5.128885, 5.074537, 5.040285, 5.020535, 
    5.010053,
  // totalHeight(5,18, 0-49)
    5.001149, 5.002726, 5.006095, 5.012916, 5.025878, 5.048788, 5.085967, 
    5.140407, 5.210714, 5.288495, 5.358942, 5.405567, 5.415976, 5.384698, 
    5.312162, 5.264491, 5.221843, 5.186554, 5.153127, 5.1055, 5.037116, 
    4.949855, 4.847899, 4.744311, 4.653742, 4.585035, 4.548517, 4.550172, 
    4.592954, 4.668444, 4.76445, 4.87837, 5.000965, 5.126472, 5.250022, 
    5.366846, 5.471569, 5.55773, 5.617738, 5.643708, 5.629535, 5.574101, 
    5.484294, 5.375281, 5.266214, 5.1731, 5.103745, 5.057774, 5.03019, 
    5.015046,
  // totalHeight(5,19, 0-49)
    5.001132, 5.00268, 5.005971, 5.012604, 5.025155, 5.04725, 5.082956, 
    5.134978, 5.201641, 5.274235, 5.337543, 5.374701, 5.373543, 5.330182, 
    5.248117, 5.187968, 5.03577, 5.00039, 4.986063, 4.964749, 4.923753, 
    4.857672, 4.777114, 4.68915, 4.603427, 4.527005, 4.473067, 4.454343, 
    4.479911, 4.545097, 4.638662, 4.751842, 4.87722, 5.008308, 5.14009, 
    5.268059, 5.38738, 5.492204, 5.575282, 5.62822, 5.642832, 5.613966, 
    5.543258, 5.441728, 5.32815, 5.222465, 5.138189, 5.079276, 5.042429, 
    5.021496,
  // totalHeight(5,20, 0-49)
    5.000885, 5.002056, 5.004517, 5.009397, 5.018436, 5.033949, 5.05833, 
    5.092862, 5.13604, 5.182454, 5.22361, 5.251111, 5.26051, 5.253445, 
    5.236856, 30, 4.882641, 4.890296, 4.897371, 4.893323, 4.87047, 4.819962, 
    4.758723, 4.686413, 4.605082, 4.517176, 4.437809, 4.388928, 4.388727, 
    4.437592, 4.525457, 4.634996, 4.760348, 4.894176, 5.031245, 5.167237, 
    5.297763, 5.417573, 5.519956, 5.596563, 5.638118, 5.636558, 5.588799, 
    5.500793, 5.388714, 5.274365, 5.176466, 5.104169, 5.057017, 5.029309,
  // totalHeight(5,21, 0-49)
    5.000641, 5.001482, 5.003266, 5.006831, 5.013499, 5.025104, 5.043731, 
    5.070997, 5.106867, 5.148563, 5.190476, 5.225755, 5.249031, 5.258772, 
    5.257997, 30, 4.74108, 4.76133, 4.784954, 4.801523, 4.801844, 4.771854, 
    4.732392, 4.676557, 4.600542, 4.503641, 4.402691, 4.328095, 4.306149, 
    4.341571, 4.42612, 4.532413, 4.657756, 4.794104, 4.93592, 5.078889, 
    5.218863, 5.351027, 5.469194, 5.565336, 5.629769, 5.652613, 5.627135, 
    5.554501, 5.447219, 5.327146, 5.217059, 5.131421, 5.073335, 5.038131,
  // totalHeight(5,22, 0-49)
    5.000444, 5.00103, 5.002293, 5.004852, 5.009718, 5.018359, 5.0326, 
    5.054197, 5.084013, 5.121048, 5.161894, 5.201262, 5.233709, 5.255754, 
    5.267343, 30, 4.627163, 4.653697, 4.689208, 4.723159, 4.745467, 4.737381, 
    4.725026, 4.694858, 4.635277, 4.538174, 4.417841, 4.312981, 4.261384, 
    4.275565, 4.351222, 4.44836, 4.569024, 4.704297, 4.848145, 4.995989, 
    5.143591, 5.286217, 5.41789, 5.530775, 5.614996, 5.659525, 5.65497, 
    5.598444, 5.498568, 5.375984, 5.256189, 5.158487, 5.089858, 5.047126,
  // totalHeight(5,23, 0-49)
    5.000326, 5.000756, 5.0017, 5.003643, 5.007394, 5.014186, 5.025643, 
    5.043532, 5.069174, 5.102598, 5.141809, 5.182737, 5.220225, 5.249777, 
    5.26927, 30, 4.542715, 4.572813, 4.616893, 4.664588, 4.705509, 4.716725, 
    4.729808, 4.725214, 4.68426, 4.591591, 4.457345, 4.326142, 4.246144, 
    4.238336, 4.303779, 4.389193, 4.502711, 4.634574, 4.778222, 4.928749, 
    5.081713, 5.232281, 5.374473, 5.500473, 5.600245, 5.662012, 5.674566, 
    5.632014, 5.539653, 5.416502, 5.289604, 5.182093, 5.104459, 5.055098,
  // totalHeight(5,24, 0-49)
    5.000295, 5.00068, 5.00153, 5.00328, 5.006674, 5.012842, 5.023315, 
    5.039814, 5.063758, 5.095514, 5.133634, 5.174624, 5.213623, 5.245886, 
    5.268474, 30, 4.488168, 4.520331, 4.569875, 4.626774, 4.680708, 4.705749, 
    4.737486, 4.751808, 4.725004, 4.637198, 4.495549, 4.347715, 4.248083, 
    4.223984, 4.28151, 4.357102, 4.464386, 4.592849, 4.73542, 4.886861, 
    5.042512, 5.19742, 5.345583, 5.479222, 5.588269, 5.660618, 5.684098, 
    5.651032, 5.564503, 5.442098, 5.311407, 5.19786, 5.114362, 5.060548,
  // totalHeight(5,25, 0-49)
    5.000359, 5.000815, 5.001808, 5.003817, 5.007643, 5.014476, 5.025854, 
    5.043424, 5.068394, 5.100799, 5.138853, 5.178908, 5.216267, 5.246636, 
    5.267615, 30, 4.464517, 4.497284, 4.548565, 4.608568, 4.667108, 4.6971, 
    4.73595, 4.757792, 4.737058, 4.652288, 4.509429, 4.356791, 4.250607, 
    4.22062, 4.27515, 4.34684, 4.451613, 4.57867, 4.72073, 4.872409, 
    5.028946, 5.185324, 5.335518, 5.471749, 5.583937, 5.659878, 5.6871, 
    5.657343, 5.572935, 5.450924, 5.319024, 5.203423, 5.117879, 5.062491,
  // totalHeight(5,26, 0-49)
    5.000526, 5.001181, 5.002566, 5.005302, 5.010374, 5.01916, 5.033297, 
    5.054275, 5.082738, 5.117734, 5.156352, 5.194211, 5.226768, 5.250868, 
    5.265858, 30, 4.47485, 4.506453, 4.555189, 4.611245, 4.664432, 4.688535, 
    4.720223, 4.735377, 4.710451, 4.625587, 4.487513, 4.343034, 4.245784, 
    4.222999, 4.281123, 4.356955, 4.46433, 4.592826, 4.735413, 4.886859, 
    5.042512, 5.19742, 5.345583, 5.479222, 5.588269, 5.660618, 5.684098, 
    5.651031, 5.564503, 5.442098, 5.311407, 5.19786, 5.114362, 5.060548,
  // totalHeight(5,27, 0-49)
    5.000805, 5.001794, 5.003833, 5.007775, 5.014898, 5.026875, 5.045452, 
    5.071789, 5.105519, 5.144054, 5.182762, 5.21631, 5.240609, 5.254356, 
    5.259472, 30, 4.523546, 4.551486, 4.592946, 4.637959, 4.676403, 4.684864, 
    4.697034, 4.693454, 4.655822, 4.568797, 4.441556, 4.316923, 4.241585, 
    4.236356, 4.302987, 4.388885, 4.502593, 4.634529, 4.778204, 4.928742, 
    5.081711, 5.232281, 5.374472, 5.500473, 5.600244, 5.662012, 5.674566, 
    5.632014, 5.539653, 5.416502, 5.289604, 5.182093, 5.104459, 5.055098,
  // totalHeight(5,28, 0-49)
    5.001189, 5.002643, 5.005589, 5.011191, 5.021119, 5.037401, 5.061837, 
    5.094956, 5.134828, 5.176611, 5.213614, 5.239749, 5.252041, 5.251792, 
    5.243953, 30, 4.61626, 4.63638, 4.665257, 4.692745, 4.709127, 4.695071, 
    4.679724, 4.649843, 4.594497, 4.505446, 4.395233, 4.299756, 4.254767, 
    4.27263, 4.350018, 4.447882, 4.568835, 4.704223, 4.848115, 4.995977, 
    5.143586, 5.286216, 5.417889, 5.530774, 5.614996, 5.659525, 5.65497, 
    5.598445, 5.498568, 5.375984, 5.256189, 5.158487, 5.089858, 5.047126,
  // totalHeight(5,29, 0-49)
    5.001638, 5.003657, 5.007708, 5.01534, 5.02871, 5.05025, 5.081713, 
    5.122604, 5.168763, 5.212454, 5.244812, 5.259601, 5.255975, 5.238696, 
    5.215979, 30, 4.757369, 4.761571, 4.770969, 4.774717, 4.763777, 4.723468, 
    4.678093, 4.621346, 4.550265, 4.463518, 4.37518, 4.311992, 4.297986, 
    4.337866, 4.424553, 4.531772, 4.657499, 4.794, 4.935878, 5.078872, 
    5.218856, 5.351024, 5.469192, 5.565335, 5.629769, 5.652613, 5.627135, 
    5.554501, 5.447219, 5.327146, 5.217059, 5.131421, 5.073335, 5.038131,
  // totalHeight(5,30, 0-49)
    5.002085, 5.004748, 5.010147, 5.020489, 5.03899, 5.069524, 5.115261, 
    5.176115, 5.24598, 5.31214, 5.358694, 5.372374, 5.346906, 5.283526, 
    5.188242, 5.105539, 4.913468, 4.864236, 4.846265, 4.829531, 4.79874, 
    4.743309, 4.680916, 4.612876, 4.541994, 4.469274, 4.40619, 4.370837, 
    4.379624, 4.433442, 4.523681, 4.634262, 4.760047, 4.894053, 5.031196, 
    5.167217, 5.297757, 5.417571, 5.519956, 5.596563, 5.638118, 5.636558, 
    5.588799, 5.500793, 5.388714, 5.274365, 5.176466, 5.104169, 5.057017, 
    5.029309,
  // totalHeight(5,31, 0-49)
    5.002143, 5.004889, 5.010488, 5.021266, 5.040632, 5.072723, 5.12099, 
    5.185519, 5.260214, 5.332315, 5.385979, 5.407974, 5.391459, 5.335916, 
    5.244624, 5.177097, 5.096328, 5.048657, 5.011378, 4.966193, 4.904812, 
    4.824902, 4.735695, 4.645541, 4.563855, 4.495916, 4.451912, 4.441776, 
    4.473276, 4.541901, 4.637214, 4.751214, 4.876952, 5.008195, 5.140043, 
    5.268041, 5.387373, 5.492201, 5.575282, 5.62822, 5.642832, 5.613966, 
    5.543258, 5.441728, 5.328151, 5.222465, 5.138189, 5.079276, 5.042429, 
    5.021496,
  // totalHeight(5,32, 0-49)
    5.001922, 5.004405, 5.009535, 5.019537, 5.037773, 5.068523, 5.115789, 
    5.180799, 5.258986, 5.338832, 5.40467, 5.442245, 5.443079, 5.405014, 
    5.329818, 5.271312, 5.264867, 5.214771, 5.161846, 5.095674, 5.012313, 
    4.915738, 4.80939, 4.706865, 4.621886, 4.561248, 4.53286, 4.540988, 
    4.588072, 4.666042, 4.76333, 4.877868, 5.000745, 5.126377, 5.249983, 
    5.366829, 5.471562, 5.557727, 5.617737, 5.643708, 5.629536, 5.574101, 
    5.484294, 5.375281, 5.266214, 5.1731, 5.103745, 5.057774, 5.03019, 
    5.015046,
  // totalHeight(5,33, 0-49)
    5.00155, 5.003578, 5.007845, 5.01632, 5.032094, 5.059364, 5.102615, 
    5.16453, 5.242973, 5.328912, 5.40777, 5.464293, 5.487687, 5.473557, 
    5.422353, 5.376557, 5.412996, 5.361646, 5.298301, 5.217968, 5.119894, 
    5.013451, 4.898541, 4.791826, 4.709034, 4.656785, 4.640617, 4.661203, 
    4.717844, 4.800365, 4.89677, 5.009197, 5.126649, 5.243997, 5.35644, 
    5.458851, 5.545294, 5.608843, 5.642066, 5.638551, 5.595541, 5.5169, 
    5.414419, 5.305392, 5.206675, 5.128885, 5.074537, 5.040285, 5.020535, 
    5.010053,
  // totalHeight(5,34, 0-49)
    5.001143, 5.002663, 5.005934, 5.012573, 5.025232, 5.04776, 5.084791, 
    5.14025, 5.21467, 5.302464, 5.391526, 5.466604, 5.514605, 5.528172, 
    5.505728, 5.478414, 5.53635, 5.487955, 5.419987, 5.331903, 5.225847, 
    5.115927, 5, 4.895658, 4.818719, 4.774924, 4.767848, 4.796153, 4.857343, 
    4.940302, 5.033179, 5.140856, 5.250273, 5.356515, 5.454584, 5.538877, 
    5.60298, 5.639935, 5.643376, 5.609665, 5.5406, 5.445177, 5.338465, 
    5.237003, 5.153089, 5.091654, 5.05119, 5.026856, 5.013346, 5.006411,
  // totalHeight(5,35, 0-49)
    5.000779, 5.001836, 5.004165, 5.009008, 5.018488, 5.035882, 5.065555, 
    5.112102, 5.1783, 5.262308, 5.355819, 5.445318, 5.51646, 5.558745, 
    5.567586, 5.563785, 5.631766, 5.591699, 5.525231, 5.435889, 5.328604, 
    5.221323, 5.110783, 5.013813, 4.944966, 4.909076, 4.90834, 4.940494, 
    5.002017, 5.0818, 5.168562, 5.26862, 5.367057, 5.45893, 5.538898, 
    5.600948, 5.638573, 5.645639, 5.618137, 5.556546, 5.467717, 5.364568, 
    5.262632, 5.174875, 5.10799, 5.062179, 5.033578, 5.017106, 5.008286, 
    5.003901,
  // totalHeight(5,36, 0-49)
    5.000493, 5.00118, 5.002732, 5.006036, 5.012685, 5.025267, 5.047535, 
    5.084073, 5.139023, 5.213765, 5.304395, 5.400975, 5.489923, 5.558537, 
    5.598734, 5.621789, 5.695973, 5.669862, 5.611474, 5.527821, 5.42626, 
    5.327377, 5.227425, 5.141449, 5.081936, 5.053137, 5.056394, 5.089209, 
    5.147419, 5.22072, 5.298621, 5.387753, 5.471721, 5.545353, 5.603, 
    5.638578, 5.646291, 5.622087, 5.565695, 5.482424, 5.383308, 5.282547, 
    5.193025, 5.122472, 5.072483, 5.040219, 5.021027, 5.010407, 5.004912, 
    5.002266,
  // totalHeight(5,37, 0-49)
    5.000292, 5.00071, 5.00168, 5.003798, 5.008177, 5.016725, 5.032395, 
    5.059221, 5.101714, 5.163327, 5.244109, 5.338745, 5.436703, 5.525202, 
    5.5934, 5.644053, 5.725108, 5.718331, 5.675017, 5.604451, 5.51567, 
    5.430519, 5.345299, 5.272915, 5.223416, 5.200871, 5.206166, 5.236938, 
    5.288577, 5.352169, 5.418102, 5.492436, 5.557827, 5.608882, 5.639949, 
    5.645644, 5.622088, 5.568674, 5.489669, 5.39456, 5.296116, 5.20661, 
    5.134175, 5.081369, 5.046282, 5.0248, 5.012568, 5.006046, 5.00278, 
    5.001256,
  // totalHeight(5,38, 0-49)
    5.000163, 5.000402, 5.000972, 5.002252, 5.004967, 5.01043, 5.02079, 
    5.039236, 5.069869, 5.116913, 5.18307, 5.267374, 5.363808, 5.462077, 
    5.550688, 5.62586, 5.715589, 5.73241, 5.710911, 5.660795, 5.591628, 
    5.525109, 5.458025, 5.401213, 5.362216, 5.345235, 5.350946, 5.377285, 
    5.419301, 5.469871, 5.520268, 5.57542, 5.617796, 5.642089, 5.643384, 
    5.61814, 5.565695, 5.489669, 5.398307, 5.302978, 5.215004, 5.142382, 
    5.088205, 5.051301, 5.028121, 5.014579, 5.007169, 5.003353, 5.001502, 
    5.000663,
  // totalHeight(5,39, 0-49)
    5.000086, 5.000216, 5.000532, 5.00126, 5.002849, 5.006141, 5.012588, 
    5.024494, 5.045127, 5.078468, 5.128332, 5.196746, 5.282134, 5.37842, 
    5.476128, 5.568144, 5.666311, 5.708275, 5.713571, 5.690119, 5.646567, 
    5.603043, 5.557014, 5.517471, 5.489532, 5.477641, 5.482416, 5.502121, 
    5.53159, 5.565724, 5.596741, 5.628298, 5.64374, 5.638564, 5.60967, 
    5.556547, 5.482424, 5.39456, 5.302978, 5.217841, 5.146606, 5.092508, 
    5.054886, 5.030718, 5.016266, 5.008171, 5.003901, 5.001774, 5.000774, 
    5.000335,
  // totalHeight(5,40, 0-49)
    5.000043, 5.00011, 5.000275, 5.000667, 5.001546, 5.00342, 5.007205, 
    5.014437, 5.02746, 5.049472, 5.084197, 5.134979, 5.203325, 5.287435, 
    5.381662, 5.479102, 5.581413, 5.64549, 5.67866, 5.685199, 5.671315, 
    5.65408, 5.631466, 5.610655, 5.594442, 5.587394, 5.59011, 5.601179, 
    5.615451, 5.629982, 5.638213, 5.642873, 5.629552, 5.595548, 5.540603, 
    5.467717, 5.383308, 5.296116, 5.215004, 5.146606, 5.093976, 5.056751, 
    5.03237, 5.017484, 5.008961, 5.004367, 5.002027, 5.000896, 5.000381, 
    5.000162,
  // totalHeight(5,41, 0-49)
    5.000021, 5.000053, 5.000136, 5.000334, 5.000796, 5.001806, 5.003906, 
    5.008049, 5.015777, 5.029372, 5.051832, 5.086515, 5.136288, 5.202295, 
    5.282791, 5.373473, 5.471925, 5.54978, 5.606205, 5.641187, 5.657415, 
    5.667536, 5.669413, 5.668134, 5.664176, 5.661833, 5.66164, 5.662522, 
    5.65977, 5.652724, 5.636606, 5.613986, 5.57411, 5.516902, 5.445177, 
    5.364569, 5.282547, 5.20661, 5.142382, 5.092508, 5.056751, 5.032938, 
    5.018123, 5.009469, 5.004705, 5.002228, 5.001004, 5.000433, 5.00018, 
    5.000075,
  // totalHeight(5,42, 0-49)
    5.00001, 5.000026, 5.000064, 5.00016, 5.000389, 5.000905, 5.002008, 
    5.004252, 5.008577, 5.016464, 5.030032, 5.051978, 5.08522, 5.132163, 
    5.193682, 5.268489, 5.354282, 5.43411, 5.503586, 5.559516, 5.601096, 
    5.635793, 5.660614, 5.678005, 5.686062, 5.688162, 5.684644, 5.674834, 
    5.655095, 5.62719, 5.588821, 5.543266, 5.484297, 5.41442, 5.338465, 
    5.262631, 5.193025, 5.134175, 5.088205, 5.054886, 5.03237, 5.018123, 
    5.009644, 5.004883, 5.002356, 5.001084, 5.000476, 5.000201, 5.000082, 
    5.000034,
  // totalHeight(5,43, 0-49)
    5.000005, 5.000013, 5.00003, 5.000073, 5.000181, 5.000431, 5.000981, 
    5.002132, 5.00442, 5.008735, 5.016428, 5.029381, 5.049916, 5.080473, 
    5.122991, 5.178202, 5.245416, 5.316042, 5.385835, 5.450653, 5.507519, 
    5.559199, 5.60148, 5.633844, 5.652066, 5.657897, 5.651314, 5.632151, 
    5.598507, 5.554525, 5.500799, 5.441729, 5.37528, 5.30539, 5.237002, 
    5.174874, 5.122472, 5.081368, 5.051301, 5.030718, 5.017484, 5.009469, 
    5.004883, 5.002399, 5.001125, 5.000504, 5.000216, 5.000089, 5.000036, 
    5.000016,
  // totalHeight(5,44, 0-49)
    5.000001, 5.000006, 5.000015, 5.000033, 5.000081, 5.000196, 5.000456, 
    5.001016, 5.002163, 5.004395, 5.008506, 5.01568, 5.027507, 5.045893, 
    5.072774, 5.109653, 5.157123, 5.211867, 5.271431, 5.332604, 5.392085, 
    5.449572, 5.500086, 5.540573, 5.56503, 5.573226, 5.564657, 5.539729, 
    5.498598, 5.447226, 5.38871, 5.328142, 5.266205, 5.206667, 5.153083, 
    5.107986, 5.07248, 5.046281, 5.028121, 5.016266, 5.008961, 5.004705, 
    5.002356, 5.001125, 5.000514, 5.000224, 5.000093, 5.000038, 5.000018, 
    5.000008,
  // totalHeight(5,45, 0-49)
    5, 5.000002, 5.000007, 5.000016, 5.000035, 5.000085, 5.000203, 5.000461, 
    5.001007, 5.002101, 5.004179, 5.007924, 5.014315, 5.024631, 5.040349, 
    5.062917, 5.093406, 5.131166, 5.175416, 5.224458, 5.275883, 5.328215, 
    5.376691, 5.416956, 5.442389, 5.451115, 5.442218, 5.416569, 5.376009, 
    5.327141, 5.274342, 5.222435, 5.173072, 5.128863, 5.091638, 5.062168, 
    5.040212, 5.024796, 5.014577, 5.00817, 5.004367, 5.002228, 5.001084, 
    5.000504, 5.000224, 5.000095, 5.00004, 5.000018, 5.000009, 5.000004,
  // totalHeight(5,46, 0-49)
    5, 5, 5.000003, 5.000008, 5.000017, 5.000037, 5.000086, 5.0002, 5.000446, 
    5.000955, 5.001951, 5.0038, 5.007055, 5.012488, 5.021063, 5.033856, 
    5.051858, 5.075415, 5.104631, 5.138946, 5.177042, 5.217485, 5.256517, 
    5.289888, 5.311668, 5.319259, 5.311596, 5.289727, 5.256232, 5.217037, 
    5.176403, 5.138111, 5.10367, 5.074477, 5.051146, 5.033548, 5.021009, 
    5.012557, 5.007162, 5.003898, 5.002025, 5.001004, 5.000476, 5.000216, 
    5.000093, 5.00004, 5.000018, 5.00001, 5.000005, 5,
  // totalHeight(5,47, 0-49)
    5, 5, 5, 5.000004, 5.00001, 5.000017, 5.000035, 5.000082, 5.000188, 
    5.000413, 5.000865, 5.001729, 5.003295, 5.005988, 5.010376, 5.017145, 
    5.027009, 5.040486, 5.057955, 5.079401, 5.10426, 5.131539, 5.158699, 
    5.182441, 5.198313, 5.203908, 5.198285, 5.182379, 5.15859, 5.131369, 
    5.104017, 5.079085, 5.057591, 5.040131, 5.026741, 5.017027, 5.010357, 
    5.006016, 5.003337, 5.001766, 5.000893, 5.000431, 5.000199, 5.000088, 
    5.000038, 5.000018, 5.00001, 5.000006, 5.000001, 5,
  // totalHeight(5,48, 0-49)
    5, 5, 5, 5, 5.000005, 5.000009, 5.000016, 5.000033, 5.000074, 5.000168, 
    5.00036, 5.000737, 5.001443, 5.002692, 5.004791, 5.008132, 5.013163, 
    5.020295, 5.029888, 5.0421, 5.056754, 5.073282, 5.09015, 5.105158, 
    5.115366, 5.118993, 5.115357, 5.105136, 5.090113, 5.073223, 5.056668, 
    5.041988, 5.029758, 5.020169, 5.013067, 5.00809, 5.004785, 5.002703, 
    5.001458, 5.00075, 5.000369, 5.000174, 5.000078, 5.000034, 5.000016, 
    5.000009, 5.000005, 5.000001, 5, 5,
  // totalHeight(5,49, 0-49)
    5, 5, 5, 5, 5, 5.000002, 5.000004, 5.00001, 5.000021, 5.000049, 5.00011, 
    5.000237, 5.000488, 5.000957, 5.001791, 5.003193, 5.005428, 5.008776, 
    5.013537, 5.019944, 5.02806, 5.037715, 5.048037, 5.057581, 5.064183, 
    5.06655, 5.064181, 5.057576, 5.048025, 5.037696, 5.028031, 5.019907, 
    5.013492, 5.008731, 5.005393, 5.003181, 5.001791, 5.000962, 5.000493, 
    5.000242, 5.000113, 5.000051, 5.000022, 5.00001, 5.000005, 5.000002, 5, 
    5, 5, 5,
  // totalHeight(6,0, 0-49)
    5.000001, 5.000006, 5.00001, 5.000018, 5.000034, 5.000072, 5.000154, 
    5.000316, 5.000631, 5.001208, 5.002222, 5.003925, 5.006657, 5.010836, 
    5.01693, 5.025394, 5.036568, 5.050474, 5.066961, 5.08557, 5.105506, 
    5.125745, 5.144631, 5.160282, 5.170508, 5.174044, 5.170405, 5.160065, 
    5.144283, 5.12525, 5.104868, 5.084815, 5.066161, 5.049734, 5.036002, 
    5.025083, 5.016811, 5.010836, 5.006715, 5.003999, 5.002289, 5.00126, 
    5.000666, 5.00034, 5.000166, 5.000079, 5.000038, 5.000019, 5.000011, 
    5.000007,
  // totalHeight(6,1, 0-49)
    5.000005, 5.00001, 5.000018, 5.000033, 5.00007, 5.000151, 5.00032, 
    5.000653, 5.001278, 5.002406, 5.004348, 5.007544, 5.012561, 5.020073, 
    5.030783, 5.045307, 5.064008, 5.086517, 5.11232, 5.140503, 5.169809, 
    5.198979, 5.225753, 5.247741, 5.261885, 5.266718, 5.261647, 5.247239, 
    5.224946, 5.197832, 5.168324, 5.13874, 5.110439, 5.084771, 5.062673, 
    5.044592, 5.030516, 5.020079, 5.012699, 5.007718, 5.004508, 5.002532, 
    5.001365, 5.000708, 5.000353, 5.00017, 5.00008, 5.000038, 5.000021, 
    5.000012,
  // totalHeight(6,2, 0-49)
    5.000009, 5.000016, 5.000031, 5.000069, 5.000152, 5.000327, 5.000679, 
    5.001356, 5.002598, 5.004784, 5.008452, 5.014331, 5.023312, 5.036367, 
    5.054408, 5.078065, 5.107471, 5.141197, 5.177971, 5.216177, 5.254053, 
    5.290477, 5.322897, 5.349, 5.365357, 5.37082, 5.364851, 5.347931, 
    5.321181, 5.288037, 5.250886, 5.212396, 5.173913, 5.137403, 5.104555, 
    5.076529, 5.053838, 5.036386, 5.023619, 5.014725, 5.008818, 5.005071, 
    5.002802, 5.001487, 5.000758, 5.000372, 5.000178, 5.000082, 5.000039, 
    5.000021,
  // totalHeight(6,3, 0-49)
    5.000015, 5.000031, 5.000066, 5.000148, 5.000325, 5.000685, 5.001394, 
    5.002722, 5.005103, 5.009176, 5.015826, 5.026171, 5.041471, 5.06295, 
    5.091514, 5.127439, 5.170224, 5.216258, 5.26322, 5.308789, 5.351055, 
    5.389846, 5.422889, 5.44876, 5.464318, 5.469281, 5.463325, 5.446671, 
    5.41954, 5.385091, 5.344875, 5.301375, 5.2552, 5.208684, 5.164347, 
    5.124405, 5.090402, 5.063021, 5.042137, 5.027025, 5.016627, 5.009819, 
    5.005565, 5.003028, 5.001583, 5.000794, 5.000385, 5.00018, 5.000083, 
    5.00004,
  // totalHeight(6,4, 0-49)
    5.000029, 5.000062, 5.00014, 5.00031, 5.000668, 5.001381, 5.002748, 
    5.005244, 5.009598, 5.016839, 5.0283, 5.045533, 5.070081, 5.103135, 
    5.145094, 5.195261, 5.252154, 5.308517, 5.361249, 5.407907, 5.447248, 
    5.481152, 5.508186, 5.528504, 5.5398, 5.542978, 5.537997, 5.524723, 
    5.502158, 5.472632, 5.436204, 5.394633, 5.346801, 5.294731, 5.241333, 
    5.189841, 5.143176, 5.103406, 5.07149, 5.047315, 5.029989, 5.018214, 
    5.010605, 5.005923, 5.003174, 5.001634, 5.000808, 5.000386, 5.00018, 
    5.000086,
  // totalHeight(6,5, 0-49)
    5.000058, 5.000128, 5.000286, 5.000626, 5.001318, 5.002669, 5.005185, 
    5.009661, 5.017243, 5.029462, 5.048134, 5.075124, 5.1119, 5.158987, 
    5.215483, 5.279093, 5.347617, 5.408614, 5.459496, 5.498811, 5.526948, 
    5.548717, 5.563705, 5.573915, 5.578139, 5.578449, 5.57507, 5.567517, 
    5.553593, 5.534558, 5.508757, 5.477044, 5.435779, 5.385819, 5.329535, 
    5.270462, 5.212655, 5.159855, 5.114769, 5.078687, 5.051541, 5.032279, 
    5.019346, 5.011106, 5.006111, 5.003226, 5.001635, 5.000797, 5.000378, 
    5.000181,
  // totalHeight(6,6, 0-49)
    5.000115, 5.000255, 5.000564, 5.001209, 5.002492, 5.00493, 5.009352, 
    5.016989, 5.029522, 5.049008, 5.077607, 5.11707, 5.168053, 5.229499, 
    5.298431, 5.370821, 5.445284, 5.502716, 5.543248, 5.567499, 5.578008, 
    5.582731, 5.581964, 5.579405, 5.574989, 5.571723, 5.570034, 5.569163, 
    5.56598, 5.56068, 5.55012, 5.534544, 5.507586, 5.468422, 5.417926, 
    5.358761, 5.295095, 5.231841, 5.173631, 5.123855, 5.084163, 5.05453, 
    5.033725, 5.019936, 5.011277, 5.006112, 5.003177, 5.001587, 5.000769, 
    5.000376,
  // totalHeight(6,7, 0-49)
    5.000226, 5.000491, 5.001064, 5.002233, 5.004501, 5.008698, 5.016093, 
    5.028466, 5.048059, 5.0773, 5.118228, 5.171681, 5.236503, 5.309232, 
    5.384604, 5.457738, 5.530963, 5.576744, 5.600434, 5.605077, 5.595113, 
    5.581197, 5.563703, 5.547695, 5.534246, 5.527015, 5.526596, 5.532055, 
    5.539679, 5.548707, 5.554925, 5.558561, 5.5509, 5.529508, 5.493343, 
    5.443217, 5.382048, 5.31462, 5.246725, 5.183888, 5.130181, 5.087585, 
    5.056075, 5.034219, 5.019936, 5.011107, 5.005926, 5.003036, 5.001507, 
    5.000752,
  // totalHeight(6,8, 0-49)
    5.000422, 5.000904, 5.001921, 5.003942, 5.007765, 5.014642, 5.026388, 
    5.045363, 5.074217, 5.115291, 5.169679, 5.236262, 5.311226, 5.388562, 
    5.461514, 5.526134, 5.591987, 5.620574, 5.624623, 5.609064, 5.579417, 
    5.548193, 5.515173, 5.486481, 5.46438, 5.452968, 5.453032, 5.463569, 
    5.480635, 5.502585, 5.524538, 5.547294, 5.560452, 5.560471, 5.544627, 
    5.511597, 5.462111, 5.399347, 5.328711, 5.256863, 5.190205, 5.133425, 
    5.088749, 5.056075, 5.033725, 5.019349, 5.010611, 5.00558, 5.002838, 
    5.001445,
  // totalHeight(6,9, 0-49)
    5.000753, 5.001589, 5.003309, 5.006641, 5.012774, 5.023482, 5.041159, 
    5.068617, 5.108491, 5.162234, 5.228955, 5.304729, 5.382974, 5.456024, 
    5.5172, 5.565434, 5.620588, 5.629872, 5.615059, 5.581898, 5.535974, 
    5.490709, 5.444725, 5.404984, 5.375036, 5.359287, 5.358814, 5.372686, 
    5.397056, 5.429439, 5.464555, 5.504181, 5.536883, 5.558599, 5.565522, 
    5.554592, 5.52423, 5.475126, 5.410761, 5.337203, 5.261992, 5.192336, 
    5.133425, 5.087586, 5.054531, 5.032286, 5.018225, 5.009846, 5.005136, 
    5.00267,
  // totalHeight(6,10, 0-49)
    5.001282, 5.002665, 5.005434, 5.010663, 5.020015, 5.035825, 5.060974, 
    5.098361, 5.149876, 5.215099, 5.290311, 5.368649, 5.441668, 5.501667, 
    5.54359, 5.570598, 5.614685, 5.605386, 5.574833, 5.52846, 5.471034, 
    5.416002, 5.360381, 5.31177, 5.275041, 5.254829, 5.25267, 5.267902, 
    5.297109, 5.337039, 5.382149, 5.435371, 5.484737, 5.526087, 5.55515, 
    5.567821, 5.560739, 5.532126, 5.482728, 5.416425, 5.34004, 5.261992, 
    5.190205, 5.130182, 5.084167, 5.051551, 5.03001, 5.016677, 5.008926, 
    5.004739,
  // totalHeight(6,11, 0-49)
    5.002078, 5.004252, 5.008497, 5.016294, 5.029826, 5.051929, 5.085682, 
    5.133456, 5.195515, 5.268737, 5.346379, 5.41946, 5.479264, 5.519618, 
    5.53792, 5.542086, 5.576544, 5.550974, 5.508726, 5.454051, 5.390294, 
    5.330138, 5.268671, 5.213834, 5.171679, 5.146977, 5.141926, 5.156423, 
    5.187869, 5.232409, 5.284306, 5.34762, 5.410196, 5.467977, 5.516637, 
    5.551656, 5.568658, 5.564036, 5.535913, 5.485223, 5.416424, 5.337204, 
    5.256864, 5.183889, 5.12386, 5.078702, 5.04735, 5.027104, 5.014899, 
    5.008082,
  // totalHeight(6,12, 0-49)
    5.003199, 5.006451, 5.012627, 5.023664, 5.042225, 5.071439, 5.11411, 
    5.171338, 5.240982, 5.31694, 5.390095, 5.450813, 5.491652, 5.508848, 
    5.502183, 5.484329, 5.5107, 5.471681, 5.42171, 5.363332, 5.298191, 
    5.237552, 5.174379, 5.116498, 5.070714, 5.04173, 5.032598, 5.044168, 
    5.075143, 5.121388, 5.177038, 5.247113, 5.3195, 5.390254, 5.455167, 
    5.509714, 5.549153, 5.568865, 5.565066, 5.535909, 5.482724, 5.41076, 
    5.328711, 5.246729, 5.17364, 5.114793, 5.071546, 5.042262, 5.023884, 
    5.013244,
  // totalHeight(6,13, 0-49)
    5.004665, 5.00928, 5.017808, 5.032618, 5.056721, 5.093204, 5.144015, 
    5.208309, 5.2812, 5.354035, 5.416568, 5.459991, 5.479059, 5.472442, 
    5.441646, 5.404009, 5.422162, 5.372473, 5.318215, 5.260051, 5.197939, 
    5.141232, 5.080792, 5.023685, 4.976696, 4.944057, 4.92978, 4.936145, 
    4.963764, 5.008761, 5.065294, 5.139062, 5.21817, 5.298661, 5.376439, 
    5.447134, 5.506054, 5.548239, 5.568853, 5.564024, 5.532117, 5.475121, 
    5.399345, 5.314625, 5.231855, 5.159892, 5.10349, 5.063205, 5.036771, 
    5.020852,
  // totalHeight(6,14, 0-49)
    5.006432, 5.012634, 5.023786, 5.042606, 5.072232, 5.115298, 5.172375, 
    5.240322, 5.311727, 5.376356, 5.424157, 5.448103, 5.445302, 5.416306, 
    5.363493, 5.308928, 5.315402, 5.257618, 5.201933, 5.147207, 5.091923, 
    5.043219, 4.99018, 4.938323, 4.893336, 4.858306, 4.838092, 4.836915, 
    4.85803, 4.898629, 4.953203, 5.027792, 5.110849, 5.19822, 5.285783, 
    5.369319, 5.444354, 5.506011, 5.549108, 5.568622, 5.560715, 5.524216, 
    5.462107, 5.382053, 5.295115, 5.212708, 5.143295, 5.09066, 5.054367, 
    5.031552,
  // totalHeight(6,15, 0-49)
    5.008353, 5.01623, 5.03002, 5.052654, 5.087132, 5.135281, 5.196004, 
    5.263953, 5.329874, 5.383046, 5.414553, 5.419429, 5.396732, 5.348141, 
    5.276179, 5.207609, 5.194048, 5.130501, 5.075865, 5.027326, 4.982164, 
    4.945155, 4.904314, 4.862773, 4.823861, 4.788546, 4.762092, 4.751051, 
    4.762189, 4.794866, 4.844478, 4.917047, 5.001487, 5.09321, 5.187871, 
    5.281279, 5.369182, 5.446979, 5.509586, 5.551565, 5.567762, 5.554559, 
    5.511582, 5.443219, 5.358788, 5.270534, 5.190001, 5.124745, 5.077209, 
    5.045891,
  // totalHeight(6,16, 0-49)
    5.010181, 5.019599, 5.035693, 5.061436, 5.099479, 5.150658, 5.212265, 
    5.277219, 5.335279, 5.376088, 5.392232, 5.380555, 5.341426, 5.277007, 
    5.189547, 5.10928, 5.061175, 4.993652, 4.942364, 4.902635, 4.870674, 
    4.848741, 4.82494, 4.799216, 4.771264, 4.738774, 4.706534, 4.683522, 
    4.680879, 4.701571, 4.742841, 4.810379, 4.893664, 4.987398, 5.086774, 
    5.187449, 5.285298, 5.376024, 5.45486, 5.516427, 5.555016, 5.565443, 
    5.544588, 5.493336, 5.417953, 5.329622, 5.241532, 5.164762, 5.10537, 
    5.064186,
  // totalHeight(6,17, 0-49)
    5.011572, 5.022128, 5.039799, 5.067472, 5.107347, 5.159363, 5.219592, 
    5.279918, 5.329862, 5.35982, 5.363729, 5.339694, 5.288814, 5.213394, 
    5.115401, 5.023416, 4.91982, 4.848852, 4.803052, 4.775018, 4.75953, 
    4.755941, 4.754036, 4.749845, 4.738373, 4.712875, 4.676379, 4.639837, 
    4.619423, 4.623429, 4.652407, 4.711521, 4.790933, 4.884343, 4.986193, 
    5.091783, 5.19697, 5.297701, 5.389572, 5.46752, 5.525795, 5.558423, 
    5.560376, 5.529471, 5.46844, 5.385913, 5.294955, 5.209147, 5.138294, 
    5.086379,
  // totalHeight(6,18, 0-49)
    5.012167, 5.023161, 5.04132, 5.069361, 5.109135, 5.160046, 5.217618, 
    5.273468, 5.317338, 5.340284, 5.337028, 5.306277, 5.249497, 5.169226, 
    5.067511, 4.957667, 4.773083, 4.697157, 4.658534, 4.645606, 4.650552, 
    4.668773, 4.693651, 4.71667, 4.727506, 4.714119, 4.676271, 4.625728, 
    4.583766, 4.56583, 4.577911, 4.624625, 4.69708, 4.787639, 4.889681, 
    4.997922, 5.108042, 5.21612, 5.318082, 5.409255, 5.484136, 5.536518, 
    5.560242, 5.550798, 5.507571, 5.435857, 5.34702, 5.255654, 5.174771, 
    5.111942,
  // totalHeight(6,19, 0-49)
    5.011673, 5.022164, 5.039426, 5.06602, 5.103715, 5.152024, 5.206848, 
    5.260324, 5.302584, 5.324714, 5.321186, 5.290559, 5.234613, 5.15659, 
    5.058802, 4.913702, 4.622737, 4.538507, 4.507798, 4.513911, 4.544353, 
    4.588445, 4.64507, 4.700685, 4.73955, 4.744065, 4.709301, 4.645968, 
    4.579593, 4.53436, 4.524497, 4.554203, 4.616135, 4.700994, 4.800754, 
    4.909312, 5.022017, 5.134962, 5.244314, 5.345772, 5.434191, 5.503454, 
    5.546865, 5.558331, 5.534452, 5.477069, 5.394795, 5.301735, 5.213065, 
    5.139863,
  // totalHeight(6,20, 0-49)
    5.009789, 5.018234, 5.032057, 5.053111, 5.08257, 5.119898, 5.161999, 
    5.20331, 5.237241, 5.258398, 5.264359, 5.256173, 5.237612, 5.213781, 
    5.189564, 30, 4.351584, 4.34895, 4.370693, 4.414233, 4.476791, 4.54938, 
    4.639208, 4.728305, 4.795688, 4.818511, 4.786697, 4.708689, 4.613272, 
    4.53438, 4.497091, 4.504663, 4.552106, 4.628093, 4.722847, 4.829231, 
    4.942132, 5.057541, 5.171772, 5.280826, 5.379914, 5.463161, 5.523698, 
    5.554443, 5.54987, 5.508664, 5.436234, 5.345024, 5.251167, 5.168735,
  // totalHeight(6,21, 0-49)
    5.008009, 5.014865, 5.026288, 5.044007, 5.069425, 5.102808, 5.142482, 
    5.184568, 5.223716, 5.254673, 5.273949, 5.280734, 5.276828, 5.265878, 
    5.252289, 30, 4.170659, 4.190443, 4.237646, 4.309671, 4.403232, 4.505134, 
    4.625941, 4.743216, 4.833209, 4.872109, 4.84777, 4.765993, 4.654385, 
    4.551601, 4.492404, 4.478347, 4.510312, 4.576025, 4.664337, 4.767112, 
    4.878688, 4.994842, 5.111915, 5.226116, 5.33296, 5.426864, 5.501005, 
    5.547768, 5.560138, 5.534248, 5.47243, 5.384887, 5.287694, 5.197131,
  // totalHeight(6,22, 0-49)
    5.006531, 5.012131, 5.021671, 5.036806, 5.059116, 5.089477, 5.127281, 
    5.16994, 5.2131, 5.25171, 5.281518, 5.300305, 5.308352, 5.308174, 
    5.303796, 30, 4.030805, 4.065196, 4.131796, 4.227709, 4.348972, 4.477757, 
    4.627515, 4.771355, 4.883232, 4.939029, 4.924598, 4.842271, 4.716929, 
    4.590865, 4.509266, 4.470721, 4.484496, 4.53761, 4.617585, 4.715239, 
    4.824254, 4.940064, 5.058887, 5.17696, 5.289956, 5.392478, 5.47778, 
    5.537942, 5.564931, 5.552924, 5.501613, 5.41886, 5.320036, 5.22286,
  // totalHeight(6,23, 0-49)
    5.005608, 5.010423, 5.018781, 5.032283, 5.052613, 5.081013, 5.117546, 
    5.160475, 5.206153, 5.249742, 5.28655, 5.313443, 5.329684, 5.337036, 
    5.339309, 30, 3.936208, 3.979444, 4.05963, 4.173486, 4.31631, 4.465572, 
    4.636799, 4.799335, 4.926097, 4.994142, 4.988685, 4.909207, 4.776904, 
    4.635037, 4.536873, 4.476786, 4.473642, 4.514404, 4.585753, 4.677729, 
    4.783483, 4.898127, 5.017705, 5.138398, 5.255899, 5.364881, 5.458617, 
    5.528984, 5.567272, 5.566283, 5.52371, 5.445437, 5.345931, 5.243716,
  // totalHeight(6,24, 0-49)
    5.005395, 5.009989, 5.017999, 5.030992, 5.050661, 5.078343, 5.114321, 
    5.157181, 5.203599, 5.248916, 5.288375, 5.318546, 5.338296, 5.349046, 
    5.354481, 30, 3.885182, 3.932935, 4.020948, 4.145664, 4.301788, 4.463101, 
    4.646461, 4.818689, 4.952569, 5.026831, 5.027077, 4.951261, 4.817554, 
    4.668488, 4.561754, 4.487683, 4.472909, 4.504726, 4.569493, 4.656837, 
    4.759587, 4.872656, 4.991975, 5.113683, 5.233487, 5.346098, 5.444815, 
    5.521412, 5.566805, 5.572984, 5.536391, 5.461555, 5.362166, 5.257078,
  // totalHeight(6,25, 0-49)
    5.005977, 5.010957, 5.019516, 5.033198, 5.053604, 5.081876, 5.118042, 
    5.160445, 5.205666, 5.249183, 5.286569, 5.314772, 5.332943, 5.342594, 
    5.347287, 30, 3.875384, 3.92374, 4.013379, 4.140702, 4.30019, 4.464015, 
    4.64996, 4.823952, 4.9589, 5.034354, 5.036249, 4.962126, 4.829005, 
    4.67878, 4.570251, 4.491889, 4.473286, 4.501997, 4.564393, 4.650023, 
    4.75163, 4.864066, 4.983222, 5.105221, 5.225766, 5.339579, 5.439962, 
    5.518659, 5.566463, 5.575105, 5.5406, 5.46701, 5.367731, 5.261695,
  // totalHeight(6,26, 0-49)
    5.007358, 5.013331, 5.023318, 5.038845, 5.061301, 5.09135, 5.128307, 
    5.169772, 5.211891, 5.250265, 5.281169, 5.302535, 5.31439, 5.318717, 
    5.319005, 30, 3.907399, 3.952108, 4.036621, 4.157588, 4.309739, 4.466147, 
    4.645107, 4.813356, 4.943969, 5.016002, 5.015329, 4.94009, 4.808348, 
    4.662022, 4.557912, 4.485681, 4.471959, 4.5043, 4.569307, 4.656758, 
    4.759554, 4.872642, 4.991968, 5.113681, 5.233484, 5.346098, 5.444815, 
    5.521413, 5.566805, 5.572984, 5.53639, 5.461555, 5.362166, 5.257078,
  // totalHeight(6,27, 0-49)
    5.009464, 5.016989, 5.029191, 5.047569, 5.07317, 5.105905, 5.143998, 
    5.18394, 5.221245, 5.251712, 5.272612, 5.283283, 5.285047, 5.280668, 
    5.273688, 30, 3.984281, 4.020194, 4.092436, 4.198112, 4.332588, 4.472099, 
    4.634583, 4.789214, 4.909461, 4.973031, 4.965724, 4.887423, 4.759062, 
    4.622608, 4.529527, 4.472963, 4.471822, 4.513583, 4.585392, 4.677572, 
    4.783415, 4.898097, 5.017692, 5.138393, 5.255897, 5.36488, 5.458617, 
    5.528984, 5.567272, 5.566283, 5.52371, 5.445437, 5.345931, 5.243716,
  // totalHeight(6,28, 0-49)
    5.012121, 5.021662, 5.036722, 5.058746, 5.08832, 5.12436, 5.163691, 
    5.201473, 5.232535, 5.253003, 5.261386, 5.258695, 5.247797, 5.232471, 
    5.216447, 30, 4.109945, 4.130611, 4.183319, 4.265604, 4.37358, 4.487952, 
    4.624791, 4.757003, 4.859302, 4.908553, 4.891548, 4.811182, 4.691791, 
    4.573579, 4.499115, 4.465442, 4.481968, 4.536459, 4.617074, 4.715014, 
    4.824155, 4.940021, 5.058867, 5.176952, 5.289953, 5.392476, 5.477779, 
    5.537941, 5.564931, 5.552924, 5.501613, 5.41886, 5.320036, 5.22286,
  // totalHeight(6,29, 0-49)
    5.01504, 5.026921, 5.045306, 5.071594, 5.1058, 5.145628, 5.186234, 
    5.221255, 5.244844, 5.253647, 5.247667, 5.229831, 5.204763, 5.177385, 
    5.151611, 30, 4.284205, 4.28185, 4.307784, 4.359859, 4.434813, 4.518023, 
    4.622173, 4.724629, 4.802577, 4.8335, 4.806474, 4.727848, 4.624166, 
    4.531176, 4.480493, 4.472147, 4.507318, 4.574645, 4.663714, 4.766834, 
    4.878564, 4.994786, 5.11189, 5.226105, 5.332955, 5.426862, 5.501004, 
    5.547768, 5.560138, 5.534248, 5.47243, 5.384888, 5.287694, 5.197131,
  // totalHeight(6,30, 0-49)
    5.01805, 5.03292, 5.056044, 5.089447, 5.133391, 5.184988, 5.237677, 
    5.28241, 5.310273, 5.315083, 5.294526, 5.249707, 5.183735, 5.100007, 
    5.000019, 4.8457, 4.545903, 4.460265, 4.430046, 4.441324, 4.48198, 
    4.537408, 4.612211, 4.688424, 4.746189, 4.764202, 4.733611, 4.662929, 
    4.579001, 4.51218, 4.48446, 4.498162, 4.54897, 4.626636, 4.722182, 
    4.82893, 4.941996, 5.057481, 5.171744, 5.280814, 5.379909, 5.463158, 
    5.523697, 5.554443, 5.54987, 5.508664, 5.436234, 5.345024, 5.251167, 
    5.168735,
  // totalHeight(6,31, 0-49)
    5.019023, 5.03479, 5.059389, 5.094986, 5.141794, 5.196579, 5.252171, 
    5.298905, 5.32757, 5.332101, 5.310494, 5.263934, 5.195178, 5.107091, 
    5.00141, 4.883553, 4.684901, 4.605775, 4.566805, 4.557559, 4.570552, 
    4.598731, 4.639916, 4.681739, 4.709561, 4.707233, 4.671093, 4.611933, 
    4.553517, 4.517052, 4.514324, 4.54877, 4.613411, 4.699682, 4.800136, 
    4.909025, 5.021885, 5.134902, 5.244286, 5.345759, 5.434185, 5.503451, 
    5.546865, 5.558331, 5.534452, 5.477069, 5.394795, 5.301735, 5.213065, 
    5.139863,
  // totalHeight(6,32, 0-49)
    5.018395, 5.033809, 5.058214, 5.094069, 5.14203, 5.199332, 5.259036, 
    5.311258, 5.346146, 5.356833, 5.340679, 5.298523, 5.232965, 5.146788, 
    5.041823, 4.942011, 4.822749, 4.747123, 4.69965, 4.673524, 4.664025, 
    4.668962, 4.681037, 4.693107, 4.696065, 4.679071, 4.64244, 4.597218, 
    4.562731, 4.552108, 4.569833, 4.620241, 4.694829, 4.786526, 4.889145, 
    4.997667, 5.107924, 5.216065, 5.318056, 5.409244, 5.484132, 5.536515, 
    5.560241, 5.550798, 5.507571, 5.435857, 5.34702, 5.255654, 5.174771, 
    5.111942,
  // totalHeight(6,33, 0-49)
    5.016522, 5.030602, 5.0534, 5.087697, 5.134883, 5.193241, 5.256811, 
    5.316042, 5.360482, 5.382006, 5.376657, 5.344406, 5.287577, 5.209101, 
    5.111249, 5.021931, 4.958303, 4.88466, 4.830286, 4.790932, 4.763344, 
    4.748603, 4.736362, 4.723997, 4.707599, 4.681181, 4.647666, 4.616824, 
    4.603018, 4.612907, 4.64622, 4.708125, 4.789161, 4.883449, 4.985752, 
    5.091572, 5.196871, 5.297654, 5.389551, 5.46751, 5.525791, 5.558421, 
    5.560375, 5.529471, 5.46844, 5.385913, 5.294955, 5.209147, 5.138294, 
    5.086379,
  // totalHeight(6,34, 0-49)
    5.013892, 5.025993, 5.046119, 5.077284, 5.121665, 5.178928, 5.244718, 
    5.310551, 5.365828, 5.401097, 5.410602, 5.392849, 5.349452, 5.283387, 
    5.197491, 5.117618, 5.088926, 5.017687, 4.958633, 4.909221, 4.867121, 
    4.835982, 4.804241, 4.772992, 4.742702, 4.71132, 4.683036, 4.66551, 
    4.668421, 4.693704, 4.738229, 4.807829, 4.892317, 4.98671, 5.086431, 
    5.187284, 5.285219, 5.375988, 5.454842, 5.516418, 5.555013, 5.565441, 
    5.544586, 5.493335, 5.417953, 5.329622, 5.241532, 5.164762, 5.10537, 
    5.064186,
  // totalHeight(6,35, 0-49)
    5.010988, 5.020812, 5.037631, 5.064511, 5.10425, 5.157928, 5.223202, 
    5.293424, 5.358673, 5.408595, 5.435466, 5.43575, 5.409719, 5.359928, 
    5.289591, 5.220821, 5.212025, 5.144827, 5.083393, 5.026625, 4.973094, 
    4.928782, 4.882309, 4.837645, 4.798489, 4.765621, 4.743443, 4.737309, 
    4.752937, 4.789107, 4.841118, 4.915183, 5.000496, 5.092699, 5.187614, 
    5.281154, 5.369122, 5.446951, 5.509573, 5.55156, 5.56776, 5.554558, 
    5.511581, 5.443218, 5.358788, 5.270534, 5.190001, 5.124745, 5.077209, 
    5.045891,
  // totalHeight(6,36, 0-49)
    5.008206, 5.015754, 5.029075, 5.051062, 5.084832, 5.132618, 5.194133, 
    5.265147, 5.33742, 5.400627, 5.445424, 5.465913, 5.46032, 5.430084, 
    5.378282, 5.323157, 5.325123, 5.264044, 5.202501, 5.140908, 5.078958, 
    5.024843, 4.968314, 4.915356, 4.871645, 4.839771, 4.823688, 4.826664, 
    4.851294, 4.894493, 4.950805, 5.026462, 5.110141, 5.197854, 5.285599, 
    5.369229, 5.444311, 5.505991, 5.549098, 5.568619, 5.560713, 5.524215, 
    5.462106, 5.382053, 5.295115, 5.212708, 5.143295, 5.09066, 5.054367, 
    5.031552,
  // totalHeight(6,37, 0-49)
    5.005801, 5.011303, 5.021308, 5.038361, 5.065549, 5.105801, 5.160549, 
    5.228139, 5.302862, 5.375661, 5.436546, 5.477478, 5.494156, 5.486094, 
    5.455472, 5.416793, 5.425346, 5.372597, 5.313364, 5.249673, 5.182581, 
    5.122284, 5.060222, 5.003567, 4.958797, 4.929513, 4.918928, 4.928662, 
    4.958955, 5.005849, 5.063618, 5.138137, 5.217677, 5.298407, 5.37631, 
    5.447072, 5.506024, 5.548225, 5.568847, 5.564021, 5.532116, 5.475121, 
    5.399345, 5.314625, 5.231855, 5.159892, 5.10349, 5.063205, 5.036771, 
    5.020852,
  // totalHeight(6,38, 0-49)
    5.003891, 5.007699, 5.014834, 5.027377, 5.048105, 5.080132, 5.126007, 
    5.186297, 5.258187, 5.335034, 5.407619, 5.466704, 5.505548, 5.521119, 
    5.513827, 5.494351, 5.508985, 5.466975, 5.412887, 5.350326, 5.281836, 
    5.219258, 5.155951, 5.099565, 5.056434, 5.03064, 5.024622, 5.038822, 
    5.071777, 5.119378, 5.175891, 5.246482, 5.319166, 5.390081, 5.455081, 
    5.509673, 5.549134, 5.568857, 5.565062, 5.535907, 5.482723, 5.41076, 
    5.32871, 5.246728, 5.17364, 5.114793, 5.071546, 5.042262, 5.023884, 
    5.013244,
  // totalHeight(6,39, 0-49)
    5.002481, 5.004988, 5.009824, 5.01858, 5.03355, 5.057617, 5.093771, 
    5.144087, 5.20835, 5.282921, 5.360754, 5.432937, 5.491165, 5.529831, 
    5.546874, 5.548873, 5.571401, 5.542856, 5.497346, 5.439801, 5.37418, 
    5.313456, 5.252906, 5.200124, 5.160659, 5.138759, 5.136208, 5.152687, 
    5.185562, 5.231051, 5.283538, 5.347201, 5.409976, 5.467864, 5.516581, 
    5.55163, 5.568645, 5.56403, 5.53591, 5.485222, 5.416424, 5.337203, 
    5.256864, 5.183889, 5.12386, 5.078702, 5.04735, 5.027104, 5.014899, 
    5.008082,
  // totalHeight(6,40, 0-49)
    5.001506, 5.003077, 5.006195, 5.012006, 5.022259, 5.039356, 5.066173, 
    5.105471, 5.158852, 5.225492, 5.301316, 5.379313, 5.451182, 5.50957, 
    5.549834, 5.574276, 5.607434, 5.595249, 5.56227, 5.514218, 5.45616, 
    5.401567, 5.34748, 5.301089, 5.266817, 5.248916, 5.24868, 5.265357, 
    5.295565, 5.336142, 5.381646, 5.435097, 5.484591, 5.526011, 5.555113, 
    5.567804, 5.56073, 5.532122, 5.482724, 5.416423, 5.340039, 5.261992, 
    5.190205, 5.130182, 5.084167, 5.051551, 5.03001, 5.016677, 5.008926, 
    5.004739,
  // totalHeight(6,41, 0-49)
    5.000872, 5.001811, 5.003726, 5.007394, 5.014062, 5.025565, 5.044321, 
    5.073099, 5.114377, 5.169344, 5.236801, 5.312582, 5.390053, 5.461687, 
    5.521057, 5.566554, 5.612437, 5.619046, 5.602568, 5.568698, 5.523036, 
    5.478834, 5.434624, 5.396982, 5.369114, 5.355171, 5.356116, 5.371006, 
    5.396053, 5.428863, 5.464231, 5.504002, 5.536785, 5.558545, 5.565493, 
    5.554577, 5.524221, 5.475122, 5.410758, 5.337202, 5.261991, 5.192336, 
    5.133424, 5.087586, 5.054531, 5.032286, 5.018225, 5.009846, 5.005136, 
    5.00267,
  // totalHeight(6,42, 0-49)
    5.000481, 5.001017, 5.00214, 5.004345, 5.008471, 5.015812, 5.028213, 
    5.048029, 5.077842, 5.119837, 5.174886, 5.241633, 5.316115, 5.392297, 
    5.463521, 5.525497, 5.583997, 5.61024, 5.613234, 5.597641, 5.568791, 
    5.538901, 5.507612, 5.480733, 5.460288, 5.450224, 5.451291, 5.462511, 
    5.480014, 5.502224, 5.524326, 5.547166, 5.560371, 5.560421, 5.544595, 
    5.511576, 5.462096, 5.399337, 5.328705, 5.25686, 5.190202, 5.133424, 
    5.088748, 5.056075, 5.033725, 5.019349, 5.010611, 5.00558, 5.002838, 
    5.001445,
  // totalHeight(6,43, 0-49)
    5.000254, 5.000546, 5.001174, 5.002439, 5.00487, 5.009325, 5.017095, 
    5.029969, 5.050164, 5.080025, 5.121449, 5.175093, 5.239628, 5.311485, 
    5.385376, 5.456191, 5.523962, 5.567801, 5.590858, 5.595832, 5.586867, 
    5.574288, 5.558316, 5.543778, 5.53159, 5.525327, 5.525582, 5.531467, 
    5.539334, 5.548489, 5.55477, 5.558441, 5.550801, 5.52943, 5.493284, 
    5.443173, 5.382017, 5.3146, 5.246713, 5.18388, 5.130176, 5.087583, 
    5.056074, 5.034219, 5.019936, 5.011107, 5.005926, 5.003036, 5.001507, 
    5.000752,
  // totalHeight(6,44, 0-49)
    5.000128, 5.000281, 5.000617, 5.00131, 5.002675, 5.005249, 5.009875, 
    5.017793, 5.030678, 5.050543, 5.079468, 5.119081, 5.169894, 5.230724, 
    5.298507, 5.369052, 5.439737, 5.495649, 5.53579, 5.560483, 5.571956, 
    5.577868, 5.578365, 5.576972, 5.573505, 5.570918, 5.569647, 5.568985, 
    5.565864, 5.560555, 5.549966, 5.534374, 5.507415, 5.468267, 5.417797, 
    5.358663, 5.295023, 5.231793, 5.1736, 5.123836, 5.084153, 5.054524, 
    5.033722, 5.019935, 5.011277, 5.006111, 5.003177, 5.001587, 5.000769, 
    5.000376,
  // totalHeight(6,45, 0-49)
    5.000063, 5.000138, 5.000311, 5.000674, 5.001407, 5.002824, 5.005446, 
    5.010069, 5.017841, 5.03027, 5.049132, 5.07621, 5.112875, 5.159539, 
    5.21521, 5.277477, 5.343553, 5.403429, 5.454043, 5.493758, 5.522719, 
    5.545506, 5.561567, 5.57276, 5.57775, 5.578548, 5.575379, 5.567812, 
    5.55373, 5.5345, 5.508538, 5.476731, 5.435433, 5.385492, 5.329256, 
    5.270243, 5.212493, 5.159744, 5.114697, 5.078644, 5.051517, 5.032265, 
    5.019338, 5.011102, 5.00611, 5.003224, 5.001634, 5.000797, 5.000378, 
    5.000181,
  // totalHeight(6,46, 0-49)
    5.000031, 5.000067, 5.00015, 5.000331, 5.000709, 5.001454, 5.002869, 
    5.005435, 5.009881, 5.017223, 5.02877, 5.046025, 5.070468, 5.103213, 
    5.144585, 5.193819, 5.249195, 5.304764, 5.3573, 5.404286, 5.444343, 
    5.479204, 5.507306, 5.528643, 5.540705, 5.544287, 5.539324, 5.525741, 
    5.502674, 5.472641, 5.435821, 5.39402, 5.3461, 5.29405, 5.24074, 
    5.189366, 5.142821, 5.103158, 5.071325, 5.047211, 5.029928, 5.018178, 
    5.010585, 5.005913, 5.00317, 5.001631, 5.000807, 5.000385, 5.000178, 
    5.000086,
  // totalHeight(6,47, 0-49)
    5.000016, 5.000032, 5.000071, 5.000156, 5.000339, 5.000712, 5.00144, 
    5.002793, 5.0052, 5.009297, 5.015947, 5.026236, 5.041384, 5.062566, 
    5.090646, 5.125872, 5.167685, 5.213145, 5.259974, 5.305874, 5.348906, 
    5.388846, 5.423281, 5.450551, 5.467137, 5.472547, 5.466381, 5.448959, 
    5.420728, 5.385215, 5.34418, 5.300195, 5.253817, 5.207319, 5.163136, 
    5.123419, 5.089652, 5.062486, 5.041776, 5.026793, 5.016487, 5.009737, 
    5.005519, 5.003005, 5.001571, 5.000789, 5.000381, 5.000178, 5.000082, 
    5.00004,
  // totalHeight(6,48, 0-49)
    5.00001, 5.000016, 5.000032, 5.00007, 5.000153, 5.000327, 5.000675, 
    5.00134, 5.002559, 5.004692, 5.008262, 5.013968, 5.022671, 5.035318, 
    5.052807, 5.075786, 5.104437, 5.137691, 5.174414, 5.213105, 5.252073, 
    5.290257, 5.324902, 5.35331, 5.371335, 5.377446, 5.370953, 5.352503, 
    5.323604, 5.288409, 5.249669, 5.210224, 5.171314, 5.134784, 5.102191, 
    5.074564, 5.052313, 5.035273, 5.022853, 5.014224, 5.008505, 5.004887, 
    5.002697, 5.001432, 5.000731, 5.000358, 5.00017, 5.000078, 5.000036, 
    5.000019,
  // totalHeight(6,49, 0-49)
    5.000003, 5.000005, 5.00001, 5.000021, 5.000048, 5.000105, 5.000226, 
    5.000469, 5.000938, 5.001801, 5.003329, 5.005904, 5.010058, 5.016455, 
    5.025851, 5.039001, 5.056527, 5.078323, 5.104247, 5.133745, 5.165843, 
    5.199856, 5.232936, 5.261728, 5.280608, 5.287194, 5.280442, 5.261369, 
    5.232347, 5.199001, 5.164706, 5.132356, 5.102732, 5.076899, 5.055445, 
    5.038478, 5.025686, 5.016487, 5.010173, 5.006035, 5.00344, 5.001884, 
    5.000993, 5.000504, 5.000246, 5.000115, 5.000053, 5.000024, 5.000012, 
    5.000007,
  // totalHeight(7,0, 0-49)
    5.000065, 5.000127, 5.000259, 5.000518, 5.001007, 5.001891, 5.003428, 
    5.005995, 5.010108, 5.016434, 5.025755, 5.038896, 5.056596, 5.079338, 
    5.107157, 5.139503, 5.175241, 5.211763, 5.247095, 5.279533, 5.307879, 
    5.331899, 5.350907, 5.364714, 5.372608, 5.374767, 5.371186, 5.361848, 
    5.346594, 5.326201, 5.300992, 5.271825, 5.239199, 5.204507, 5.169468, 
    5.135854, 5.105211, 5.078644, 5.05671, 5.039443, 5.026458, 5.017118, 
    5.010684, 5.006434, 5.003739, 5.002098, 5.001138, 5.000597, 5.000308, 
    5.000164,
  // totalHeight(7,1, 0-49)
    5.000121, 5.000238, 5.00048, 5.000947, 5.001812, 5.003347, 5.005964, 
    5.010249, 5.016973, 5.027078, 5.041602, 5.061525, 5.087564, 5.119916, 
    5.158052, 5.20067, 5.245986, 5.289452, 5.328742, 5.362245, 5.389309, 
    5.411021, 5.42722, 5.438537, 5.444373, 5.445482, 5.441986, 5.433731, 
    5.419994, 5.40147, 5.377745, 5.349227, 5.315303, 5.277005, 5.236064, 
    5.194644, 5.154975, 5.118989, 5.08803, 5.062733, 5.043062, 5.028478, 
    5.018152, 5.011154, 5.00661, 5.003779, 5.002086, 5.001116, 5.000584, 
    5.000315,
  // totalHeight(7,2, 0-49)
    5.000235, 5.000459, 5.00091, 5.001763, 5.003306, 5.005982, 5.010434, 
    5.017533, 5.028368, 5.04416, 5.066104, 5.095097, 5.131435, 5.174539, 
    5.222845, 5.274029, 5.325931, 5.371635, 5.409235, 5.437857, 5.457925, 
    5.47228, 5.481415, 5.48696, 5.488639, 5.487854, 5.484875, 5.479411, 
    5.470135, 5.457471, 5.440103, 5.41785, 5.388554, 5.352391, 5.310528, 
    5.264997, 5.218402, 5.17348, 5.132623, 5.097514, 5.068947, 5.046889, 
    5.030686, 5.019336, 5.011737, 5.006867, 5.003877, 5.00212, 5.001133, 
    5.000619,
  // totalHeight(7,3, 0-49)
    5.000447, 5.000865, 5.001686, 5.003202, 5.005878, 5.010405, 5.017734, 
    5.029084, 5.045851, 5.069425, 5.100871, 5.14055, 5.18778, 5.240693, 
    5.296419, 5.351787, 5.405229, 5.447082, 5.476982, 5.495352, 5.503921, 
    5.507381, 5.506683, 5.504385, 5.500591, 5.497306, 5.494962, 5.493176, 
    5.490098, 5.485869, 5.478354, 5.466926, 5.447763, 5.419919, 5.383484, 
    5.339691, 5.290837, 5.239985, 5.190429, 5.145115, 5.106135, 5.074507, 
    5.050228, 5.032541, 5.020276, 5.012163, 5.007035, 5.003933, 5.00215, 
    5.001194,
  // totalHeight(7,4, 0-49)
    5.00083, 5.001577, 5.003015, 5.005607, 5.010071, 5.01742, 5.028973, 
    5.046284, 5.070925, 5.104134, 5.146344, 5.196767, 5.253208, 5.312281, 
    5.370041, 5.423226, 5.472451, 5.504696, 5.522296, 5.52714, 5.522073, 
    5.513369, 5.501997, 5.491229, 5.481532, 5.475423, 5.473501, 5.47537, 
    5.478836, 5.483813, 5.487583, 5.489424, 5.484031, 5.469409, 5.444396, 
    5.408932, 5.364272, 5.312967, 5.258545, 5.204911, 5.155597, 5.11315, 
    5.078824, 5.052646, 5.033748, 5.020789, 5.012327, 5.007061, 5.003947, 
    5.002234,
  // totalHeight(7,5, 0-49)
    5.00148, 5.002769, 5.005187, 5.009442, 5.016574, 5.027974, 5.045319, 
    5.070355, 5.104497, 5.148292, 5.200894, 5.259817, 5.321171, 5.380404, 
    5.433293, 5.477595, 5.517872, 5.536584, 5.539735, 5.53039, 5.512024, 
    5.492009, 5.470812, 5.452157, 5.436851, 5.427817, 5.425859, 5.430663, 
    5.439898, 5.453335, 5.467922, 5.483245, 5.492867, 5.494058, 5.484577, 
    5.462999, 5.429098, 5.384137, 5.330914, 5.273443, 5.216244, 5.163455, 
    5.118066, 5.081542, 5.053911, 5.034173, 5.020812, 5.012223, 5.006996, 
    5.004036,
  // totalHeight(7,6, 0-49)
    5.002537, 5.004672, 5.008571, 5.015256, 5.026145, 5.042995, 5.067703, 
    5.101876, 5.146226, 5.199944, 5.260352, 5.323129, 5.38313, 5.435542, 
    5.476911, 5.507005, 5.535779, 5.539415, 5.528361, 5.50633, 5.476847, 
    5.447856, 5.418829, 5.393694, 5.373574, 5.361693, 5.35911, 5.365716, 
    5.379266, 5.39945, 5.423106, 5.450462, 5.474294, 5.491517, 5.499191, 
    5.494801, 5.476672, 5.444415, 5.399313, 5.344433, 5.284281, 5.224, 
    5.16831, 5.120595, 5.082476, 5.053929, 5.033796, 5.020385, 5.011956, 
    5.007038,
  // totalHeight(7,7, 0-49)
    5.004174, 5.007567, 5.013592, 5.023635, 5.039485, 5.063149, 5.09643, 
    5.140269, 5.194015, 5.254954, 5.318458, 5.378851, 5.430717, 5.47008, 
    5.495052, 5.507923, 5.524962, 5.513952, 5.490565, 5.458614, 5.421184, 
    5.386325, 5.352101, 5.322395, 5.298602, 5.284111, 5.280297, 5.287394, 
    5.303493, 5.328266, 5.358603, 5.39561, 5.431551, 5.463284, 5.487547, 
    5.501169, 5.501382, 5.486283, 5.455358, 5.409954, 5.353441, 5.290848, 
    5.227934, 5.169954, 5.120609, 5.081582, 5.052734, 5.032722, 5.019694, 
    5.011834,
  // totalHeight(7,8, 0-49)
    5.006591, 5.011756, 5.020663, 5.035065, 5.057024, 5.088521, 5.130782, 
    5.183451, 5.243975, 5.307598, 5.368227, 5.41984, 5.457864, 5.479952, 
    5.486041, 5.480951, 5.487695, 5.463608, 5.430469, 5.391768, 5.349826, 
    5.31244, 5.275925, 5.243874, 5.217835, 5.201171, 5.195599, 5.201853, 
    5.21865, 5.245731, 5.280169, 5.3241, 5.369467, 5.413232, 5.452092, 
    5.482594, 5.501349, 5.505374, 5.492573, 5.462371, 5.416243, 5.357937, 
    5.29305, 5.227945, 5.16834, 5.118135, 5.078969, 5.050519, 5.031245, 
    5.019186,
  // totalHeight(7,9, 0-49)
    5.009975, 5.017505, 5.030089, 5.049776, 5.078679, 5.118333, 5.168806, 
    5.227921, 5.291047, 5.351834, 5.403693, 5.44137, 5.461924, 5.464885, 
    5.451752, 5.429615, 5.428216, 5.392973, 5.352669, 5.310205, 5.26699, 
    5.230297, 5.194464, 5.162518, 5.135951, 5.117805, 5.110119, 5.114284, 
    5.12995, 5.157085, 5.193079, 5.241197, 5.293196, 5.346199, 5.396987, 
    5.442087, 5.477869, 5.500757, 5.507577, 5.49611, 5.465787, 5.418324, 
    5.357944, 5.290869, 5.224051, 5.163567, 5.113378, 5.074952, 5.047724, 
    5.029982,
  // totalHeight(7,10, 0-49)
    5.01446, 5.02496, 5.041936, 5.067563, 5.103665, 5.150827, 5.207461, 
    5.269351, 5.330144, 5.382782, 5.421267, 5.441902, 5.443639, 5.42762, 
    5.396376, 5.358976, 5.351389, 5.30677, 5.26151, 5.217797, 5.176116, 
    5.143035, 5.110799, 5.081596, 5.056532, 5.03793, 5.028039, 5.029017, 
    5.041786, 5.066779, 5.101882, 5.151564, 5.207518, 5.267011, 5.326935, 
    5.383892, 5.434252, 5.474237, 5.500106, 5.508534, 5.497243, 5.465786, 
    5.416254, 5.353475, 5.284362, 5.216415, 5.155936, 5.106784, 5.070136, 
    5.045145,
  // totalHeight(7,11, 0-49)
    5.020058, 5.034059, 5.055914, 5.087668, 5.130448, 5.183438, 5.24315, 
    5.303562, 5.357356, 5.397788, 5.420244, 5.422883, 5.40632, 5.37279, 
    5.325267, 5.274648, 5.261842, 5.209301, 5.160816, 5.117825, 5.079991, 
    5.053068, 5.027225, 5.003541, 4.982328, 4.9647, 4.952865, 4.949788, 
    4.957981, 4.978666, 5.010483, 5.059205, 5.116598, 5.180028, 5.246441, 
    5.312511, 5.374698, 5.429252, 5.472255, 5.499822, 5.50852, 5.4961, 
    5.46238, 5.410001, 5.344549, 5.27369, 5.205394, 5.146018, 5.099126, 
    5.065478,
  // totalHeight(7,12, 0-49)
    5.026608, 5.044453, 5.071303, 5.108771, 5.156913, 5.213257, 5.272523, 
    5.327488, 5.37078, 5.396759, 5.402548, 5.387994, 5.354888, 5.305989, 
    5.244225, 5.182299, 5.163545, 5.104256, 5.053853, 5.013101, 4.980991, 
    4.962399, 4.945583, 4.930279, 4.915555, 4.900771, 4.887709, 4.880032, 
    4.882082, 4.896287, 4.922391, 4.967634, 5.024047, 5.089039, 5.159525, 
    5.232173, 5.303509, 5.369896, 5.427476, 5.472199, 5.500046, 5.507537, 
    5.492572, 5.455415, 5.399471, 5.33125, 5.259198, 5.191624, 5.134699, 
    5.091459,
  // totalHeight(7,13, 0-49)
    5.033735, 5.05548, 5.086987, 5.129162, 5.180753, 5.237656, 5.293234, 
    5.339825, 5.370763, 5.381915, 5.372065, 5.342326, 5.295123, 5.233254, 
    5.159248, 5.08756, 5.059693, 4.994692, 4.943421, 4.906126, 4.881305, 
    4.872905, 4.867583, 4.863523, 4.858131, 4.848498, 4.835467, 4.823103, 
    4.817653, 4.823181, 4.841021, 4.880143, 4.933115, 4.997382, 5.069714, 
    5.146647, 5.224686, 5.300283, 5.36973, 5.429057, 5.474072, 5.500647, 
    5.505333, 5.486337, 5.44461, 5.384568, 5.313798, 5.241476, 5.176003, 
    5.123024,
  // totalHeight(7,14, 0-49)
    5.040861, 5.066214, 5.101596, 5.147029, 5.199935, 5.254867, 5.304424, 
    5.34119, 5.35965, 5.357197, 5.333939, 5.29176, 5.233256, 5.160916, 
    5.076638, 4.99614, 4.952772, 4.88308, 4.831912, 4.799187, 4.783082, 
    4.786512, 4.794985, 4.804932, 4.811784, 4.809976, 4.798848, 4.782353, 
    4.768427, 4.763132, 4.769983, 4.80008, 4.846959, 4.908147, 4.980169, 
    5.059281, 5.141819, 5.224236, 5.302959, 5.374205, 5.433871, 5.477612, 
    5.501223, 5.501401, 5.476885, 5.429611, 5.365265, 5.292587, 5.221282, 
    5.159416,
  // totalHeight(7,15, 0-49)
    5.04727, 5.075588, 5.113734, 5.160819, 5.213135, 5.26433, 5.306828, 
    5.333897, 5.341276, 5.327645, 5.294003, 5.242578, 5.175807, 5.095669, 
    5.003297, 4.913842, 4.844732, 4.771318, 4.721283, 4.694343, 4.688432, 
    4.705205, 4.729593, 4.756072, 4.777933, 4.786829, 4.780121, 4.760928, 
    4.738266, 4.720271, 4.713288, 4.731091, 4.768864, 4.824393, 4.893883, 
    4.973128, 5.058129, 5.145205, 5.230836, 5.311429, 5.383089, 5.441543, 
    5.482284, 5.501088, 5.494987, 5.46355, 5.410028, 5.341596, 5.268045, 
    5.19916,
  // totalHeight(7,16, 0-49)
    5.052221, 5.082582, 5.122238, 5.169528, 5.219952, 5.266737, 5.302544, 
    5.321485, 5.320392, 5.298859, 5.258375, 5.201202, 5.129457, 5.044556, 
    4.946846, 4.846074, 4.737124, 4.660678, 4.612901, 4.593229, 4.599227, 
    4.630776, 4.672967, 4.718068, 4.757268, 4.779699, 4.780499, 4.761142, 
    4.730637, 4.698801, 4.675304, 4.677201, 4.702387, 4.749299, 4.813816, 
    4.891094, 4.976588, 5.066315, 5.156695, 5.244262, 5.325356, 5.395911, 
    5.45143, 5.487248, 5.499257, 5.485078, 5.445483, 5.385374, 5.313462, 
    5.240213,
  // totalHeight(7,17, 0-49)
    5.055084, 5.086399, 5.126359, 5.172816, 5.22089, 5.263784, 5.294598, 
    5.308188, 5.302143, 5.27656, 5.233084, 5.173849, 5.100662, 5.014484, 
    4.914962, 4.796424, 4.630887, 4.5516, 4.507199, 4.496636, 4.516641, 
    4.564325, 4.625845, 4.690973, 4.749099, 4.787496, 4.799221, 4.783396, 
    4.747558, 4.702156, 4.66026, 4.64256, 4.651261, 4.686162, 4.742951, 
    4.81599, 4.899972, 4.990417, 5.083542, 5.175914, 5.264064, 5.344178, 
    5.411934, 5.462564, 5.491307, 5.494365, 5.470315, 5.421548, 5.354854, 
    5.280277,
  // totalHeight(7,18, 0-49)
    5.055455, 5.086561, 5.125804, 5.170914, 5.217056, 5.257705, 5.286389, 
    5.298403, 5.291608, 5.26616, 5.223593, 5.165879, 5.094666, 5.010685, 
    4.912883, 4.764289, 4.52522, 4.443193, 4.403152, 4.403866, 4.440429, 
    4.50552, 4.587378, 4.673081, 4.750764, 4.806866, 4.832855, 4.825094, 
    4.788147, 4.731499, 4.671028, 4.630623, 4.61889, 4.638094, 4.684124, 
    4.750472, 4.830854, 4.920098, 5.014065, 5.109241, 5.202271, 5.289577, 
    5.367074, 5.430085, 5.473558, 5.492756, 5.484509, 5.448822, 5.390132, 
    5.31718,
  // totalHeight(7,19, 0-49)
    5.053221, 5.082938, 5.120615, 5.164308, 5.209677, 5.250699, 5.281166, 
    5.296271, 5.293453, 5.272348, 5.234126, 5.180676, 5.113756, 5.033909, 
    4.938658, 4.742922, 4.415196, 4.33217, 4.297563, 4.311978, 4.368104, 
    4.45188, 4.554541, 4.660558, 4.75763, 4.832474, 4.875569, 4.880461, 
    4.847667, 4.784114, 4.707324, 4.64267, 4.607326, 4.607371, 4.639596, 
    4.696743, 4.771411, 4.857562, 4.950556, 5.046688, 5.142635, 5.234991, 
    5.319911, 5.392896, 5.448824, 5.4824, 5.489161, 5.467055, 5.418115, 
    5.349228,
  // totalHeight(7,20, 0-49)
    5.047519, 5.072911, 5.105344, 5.143125, 5.182673, 5.219129, 5.247638, 
    5.264693, 5.268921, 5.261077, 5.243481, 5.219299, 5.191885, 5.164235, 
    5.138397, 30, 4.114454, 4.114334, 4.146542, 4.211831, 4.306983, 4.4182, 
    4.544752, 4.671088, 4.786033, 4.877743, 4.936459, 4.953573, 4.925799, 
    4.857228, 4.766321, 4.677095, 4.616313, 4.594654, 4.610526, 4.65621, 
    4.723191, 4.804475, 4.894822, 4.990243, 5.087366, 5.182891, 5.273173, 
    5.353907, 5.420018, 5.465905, 5.486187, 5.477157, 5.438637, 5.375458,
  // totalHeight(7,21, 0-49)
    5.042906, 5.065928, 5.096264, 5.132921, 5.173195, 5.212954, 5.247571, 
    5.273136, 5.287375, 5.289968, 5.282302, 5.266943, 5.247061, 5.225951, 
    5.206573, 30, 3.960332, 3.978011, 4.033281, 4.12433, 4.2451, 4.375662, 
    4.518851, 4.658369, 4.784651, 4.88853, 4.961393, 4.993842, 4.979385, 
    4.918301, 4.827318, 4.723927, 4.643672, 4.602317, 4.601614, 4.634759, 
    4.692778, 4.76789, 4.85425, 4.947518, 5.044199, 5.141039, 5.234534, 
    5.320562, 5.394155, 5.449563, 5.480793, 5.482881, 5.453789, 5.39637,
  // totalHeight(7,22, 0-49)
    5.039219, 5.060489, 5.089365, 5.125412, 5.166588, 5.209273, 5.24895, 
    5.281309, 5.303318, 5.313817, 5.313527, 5.304658, 5.290368, 5.274252, 
    5.259961, 30, 3.835406, 3.868202, 3.942687, 4.05515, 4.197188, 4.343217, 
    4.499814, 4.650155, 4.786009, 4.900363, 4.985329, 5.030774, 5.027747, 
    4.973923, 4.885179, 4.770913, 4.6747, 4.616134, 4.600175, 4.62134, 
    4.670562, 4.739481, 4.821707, 4.912546, 5.008337, 5.105797, 5.201505, 
    5.291459, 5.370781, 5.433647, 5.473652, 5.484908, 5.46392, 5.41185,
  // totalHeight(7,23, 0-49)
    5.037024, 5.057234, 5.085255, 5.120999, 5.162849, 5.207517, 5.250546, 
    5.287356, 5.314402, 5.329967, 5.334363, 5.329612, 5.318913, 5.30611, 
    5.295335, 30, 3.75083, 3.794178, 3.882296, 4.009888, 4.166729, 4.322514, 
    4.487185, 4.643687, 4.784962, 4.90581, 4.999001, 5.054017, 5.060269, 
    5.013733, 4.929824, 4.809685, 4.70313, 4.632049, 4.604081, 4.615284, 
    4.656912, 4.720334, 4.798786, 4.887294, 4.982037, 5.079676, 5.176805, 
    5.269478, 5.352865, 5.421083, 5.467453, 5.485446, 5.470525, 5.42257,
  // totalHeight(7,24, 0-49)
    5.036716, 5.05663, 5.084397, 5.120026, 5.162042, 5.207297, 5.25141, 
    5.289758, 5.318656, 5.336201, 5.342546, 5.339622, 5.330624, 5.319474, 
    5.310493, 30, 3.710093, 3.758837, 3.854186, 3.98978, 4.154303, 4.314251, 
    4.482039, 4.640524, 4.783451, 4.906882, 5.004126, 5.064573, 5.076762, 
    5.03577, 4.956805, 4.834767, 4.72329, 4.645191, 4.609799, 4.614413, 
    4.65074, 4.710127, 4.785641, 4.872161, 4.96578, 5.063129, 5.160812, 
    5.254916, 5.340633, 5.41205, 5.462324, 5.484553, 5.473571, 5.428463,
  // totalHeight(7,25, 0-49)
    5.038471, 5.058876, 5.086976, 5.122606, 5.164133, 5.208367, 5.251034, 
    5.287758, 5.315138, 5.33149, 5.337061, 5.33376, 5.324667, 5.313553, 
    5.304569, 30, 3.712392, 3.76137, 3.857336, 3.993675, 4.158824, 4.318006, 
    4.484923, 4.642324, 4.784227, 4.907133, 5.004549, 5.065886, 5.079467, 
    5.040195, 4.963305, 4.841302, 4.72898, 4.649186, 4.611698, 4.614275, 
    4.648862, 4.706868, 4.781345, 4.867144, 4.960334, 5.057543, 5.155376, 
    5.249931, 5.336409, 5.408885, 5.460465, 5.484119, 5.474478, 5.430358,
  // totalHeight(7,26, 0-49)
    5.042217, 5.063863, 5.092844, 5.128556, 5.168951, 5.210625, 5.24946, 
    5.281579, 5.304241, 5.31635, 5.31849, 5.312615, 5.301614, 5.288908, 
    5.278151, 30, 3.755883, 3.80003, 3.890133, 4.020155, 4.179138, 4.333121, 
    4.495686, 4.649438, 4.788105, 4.907743, 5.001677, 5.059398, 5.069646, 
    5.02778, 4.949212, 4.828493, 4.718805, 4.642381, 4.608218, 4.613591, 
    4.650334, 4.709931, 4.785549, 4.872119, 4.96576, 5.06312, 5.160808, 
    5.254914, 5.340632, 5.412049, 5.462324, 5.484553, 5.473571, 5.428463,
  // totalHeight(7,27, 0-49)
    5.047648, 5.071205, 5.101556, 5.137453, 5.176219, 5.214128, 5.247229, 
    5.272307, 5.287539, 5.292675, 5.288845, 5.278172, 5.26337, 5.247412, 
    5.233242, 30, 3.837907, 3.872372, 3.950503, 4.067498, 4.213774, 4.358329, 
    4.513062, 4.660518, 4.793601, 4.907108, 4.993864, 5.043576, 5.046104, 
    4.997985, 4.914999, 4.797587, 4.69459, 4.626752, 4.60112, 4.613746, 
    4.65615, 4.719967, 4.798612, 4.887213, 4.981999, 5.079659, 5.176796, 
    5.269475, 5.352864, 5.421082, 5.467452, 5.485446, 5.470524, 5.42257,
  // totalHeight(7,28, 0-49)
    5.054279, 5.08032, 5.1125, 5.148775, 5.185695, 5.219107, 5.245215, 
    5.261521, 5.267226, 5.263089, 5.25097, 5.233331, 5.212831, 5.192018, 
    5.172996, 30, 3.95486, 3.975625, 4.036456, 4.134297, 4.261631, 4.392307, 
    4.535101, 4.672795, 4.797129, 4.90109, 4.976916, 5.014869, 5.006731, 
    4.951005, 4.863965, 4.753953, 4.662951, 4.608952, 4.596192, 4.619275, 
    4.669537, 4.738986, 4.821471, 4.912435, 5.008284, 5.105772, 5.201493, 
    5.291453, 5.370779, 5.433645, 5.473652, 5.484908, 5.46392, 5.41185,
  // totalHeight(7,29, 0-49)
    5.061519, 5.090569, 5.125088, 5.162135, 5.197347, 5.22602, 5.244443, 
    5.250815, 5.245413, 5.230116, 5.207698, 5.181172, 5.153317, 5.126302, 
    5.101217, 30, 4.100039, 4.105047, 4.144559, 4.218102, 4.320959, 4.433148, 
    4.559563, 4.683653, 4.795854, 4.887011, 4.948723, 4.97219, 4.951942, 
    4.889277, 4.801144, 4.70358, 4.629909, 4.594042, 4.597061, 4.6324, 
    4.6916, 4.767314, 4.853972, 4.947385, 5.044137, 5.141009, 5.23452, 
    5.320555, 5.394152, 5.449561, 5.480793, 5.482881, 5.453789, 5.396369,
  // totalHeight(7,30, 0-49)
    5.069942, 5.104444, 5.145037, 5.188226, 5.228665, 5.260446, 5.278681, 
    5.280539, 5.265384, 5.23421, 5.188872, 5.131349, 5.06307, 4.983942, 
    4.890614, 4.694397, 4.378685, 4.306954, 4.281877, 4.30549, 4.370964, 
    4.459809, 4.568273, 4.679267, 4.780853, 4.860884, 4.909776, 4.919673, 
    4.888474, 4.82117, 4.735869, 4.654694, 4.601761, 4.586124, 4.605887, 
    4.653808, 4.721985, 4.803879, 4.89453, 4.990101, 5.087297, 5.182858, 
    5.273158, 5.353899, 5.420014, 5.465903, 5.486187, 5.477157, 5.438637, 
    5.375458,
  // totalHeight(7,31, 0-49)
    5.073872, 5.110393, 5.153061, 5.197888, 5.238931, 5.269813, 5.28551, 
    5.283435, 5.26344, 5.227028, 5.17638, 5.113566, 5.040033, 4.956133, 
    4.860312, 4.711382, 4.476999, 4.403505, 4.371749, 4.381316, 4.427418, 
    4.499416, 4.589086, 4.681817, 4.765648, 4.827684, 4.859194, 4.855018, 
    4.817186, 4.75356, 4.681082, 4.623222, 4.59458, 4.599795, 4.6354, 
    4.694525, 4.770272, 4.856986, 4.950268, 5.046546, 5.142564, 5.234956, 
    5.319895, 5.392888, 5.448821, 5.482398, 5.48916, 5.467055, 5.418115, 
    5.349227,
  // totalHeight(7,32, 0-49)
    5.074563, 5.111968, 5.156186, 5.203183, 5.24673, 5.279979, 5.297396, 
    5.296023, 5.275575, 5.23764, 5.184599, 5.118748, 5.041742, 4.954269, 
    4.855663, 4.736937, 4.571723, 4.498174, 4.459996, 4.456672, 4.485158, 
    4.540483, 4.610906, 4.684608, 4.750361, 4.79529, 4.81181, 4.797491, 
    4.758013, 4.70317, 4.647774, 4.613843, 4.608014, 4.631615, 4.680494, 
    4.748522, 4.829835, 4.919573, 5.013799, 5.109106, 5.202204, 5.289543, 
    5.367058, 5.430077, 5.473555, 5.492754, 5.484507, 5.448821, 5.390131, 
    5.31718,
  // totalHeight(7,33, 0-49)
    5.072055, 5.109157, 5.154137, 5.203316, 5.250513, 5.288494, 5.311002, 
    5.31429, 5.297483, 5.261912, 5.210007, 5.14432, 5.066876, 4.978845, 
    4.880323, 4.778907, 4.66792, 4.594558, 4.550687, 4.536237, 4.549191, 
    4.588276, 4.639575, 4.693966, 4.741624, 4.770691, 4.775239, 4.755387, 
    4.719284, 4.677091, 4.640542, 4.628673, 4.642346, 4.680838, 4.739939, 
    4.814349, 4.8991, 4.989961, 5.083307, 5.175795, 5.264003, 5.344147, 
    5.411918, 5.462556, 5.491303, 5.494362, 5.470314, 5.421547, 5.354854, 
    5.280277,
  // totalHeight(7,34, 0-49)
    5.066685, 5.102252, 5.146866, 5.197575, 5.248649, 5.292713, 5.322759, 
    5.333969, 5.324487, 5.295034, 5.247876, 5.185752, 5.11112, 5.025746, 
    4.930516, 4.839296, 4.766814, 4.694075, 4.645786, 4.622183, 4.62171, 
    4.645421, 4.67846, 4.714131, 4.744484, 4.759594, 4.755527, 4.734432, 
    4.705405, 4.677551, 4.65919, 4.666082, 4.695303, 4.745059, 4.811397, 
    4.889759, 4.975869, 5.065935, 5.156497, 5.244161, 5.325305, 5.395886, 
    5.451417, 5.487242, 5.499254, 5.485077, 5.445483, 5.385374, 5.313462, 
    5.240213,
  // totalHeight(7,35, 0-49)
    5.059091, 5.091941, 5.134801, 5.18574, 5.23992, 5.290249, 5.329171, 
    5.350695, 5.351656, 5.331776, 5.292833, 5.237574, 5.16882, 5.088939, 
    4.999584, 4.915709, 4.867932, 4.796804, 4.745568, 4.71463, 4.70265, 
    4.712214, 4.728501, 4.746943, 4.761694, 4.765309, 4.755863, 4.73676, 
    4.716686, 4.702873, 4.700494, 4.722412, 4.763369, 4.821098, 4.89199, 
    4.972076, 5.057559, 5.144899, 5.230677, 5.311346, 5.383048, 5.441524, 
    5.482273, 5.501082, 5.494984, 5.463549, 5.410028, 5.341596, 5.268045, 
    5.19916,
  // totalHeight(7,36, 0-49)
    5.050116, 5.079262, 5.118917, 5.168323, 5.223925, 5.279467, 5.327296, 
    5.360398, 5.374112, 5.366771, 5.339256, 5.293997, 5.233984, 5.162076, 
    5.080613, 5.003589, 4.970191, 4.901921, 4.849092, 4.81234, 4.790542, 
    4.787408, 4.788884, 4.792263, 4.793777, 4.788606, 4.776517, 4.761394, 
    4.750595, 4.749277, 4.760054, 4.793442, 4.842779, 4.90564, 4.978724, 
    5.058472, 5.141376, 5.223999, 5.302834, 5.37414, 5.433838, 5.477597, 
    5.501214, 5.501397, 5.476884, 5.429609, 5.365265, 5.292587, 5.221282, 
    5.159416,
  // totalHeight(7,37, 0-49)
    5.040674, 5.065457, 5.100637, 5.146596, 5.201307, 5.259878, 5.315217, 
    5.359754, 5.387404, 5.394824, 5.381534, 5.34921, 5.300679, 5.239072, 
    5.167283, 5.097776, 5.072126, 5.007897, 4.954634, 4.913358, 4.883272, 
    4.869039, 4.857895, 4.848771, 4.839742, 4.828416, 4.815767, 4.805543, 
    4.803319, 4.812391, 4.833456, 4.87515, 4.92999, 4.995509, 5.06863, 
    5.146039, 5.224351, 5.300103, 5.369635, 5.429007, 5.474048, 5.500636, 
    5.505328, 5.486333, 5.444608, 5.384567, 5.313798, 5.241476, 5.176003, 
    5.123024,
  // totalHeight(7,38, 0-49)
    5.031587, 5.051754, 5.081593, 5.122414, 5.173713, 5.232343, 5.292474, 
    5.346719, 5.387997, 5.411265, 5.414304, 5.39752, 5.363111, 5.314147, 
    5.253855, 5.193147, 5.17178, 5.112633, 5.059998, 5.015416, 4.978568, 
    4.954986, 4.933573, 4.914676, 4.897844, 4.882706, 4.870935, 4.86574, 
    4.870833, 4.888049, 4.916724, 4.963934, 5.021742, 5.087658, 5.158724, 
    5.231721, 5.303259, 5.369761, 5.427405, 5.472163, 5.500027, 5.507529, 
    5.492567, 5.455412, 5.39947, 5.33125, 5.259198, 5.191624, 5.134699, 
    5.091459,
  // totalHeight(7,39, 0-49)
    5.023478, 5.03917, 5.063326, 5.09785, 5.143517, 5.198998, 5.260269, 
    5.32098, 5.373845, 5.412485, 5.432821, 5.433532, 5.415639, 5.38168, 
    5.334877, 5.284673, 5.266556, 5.213517, 5.162659, 5.11611, 5.074186, 
    5.043216, 5.01401, 4.988095, 4.966056, 4.949053, 4.939028, 4.938462, 
    4.949347, 4.97249, 5.0063, 5.056495, 5.114914, 5.179015, 5.245848, 
    5.312171, 5.374506, 5.429146, 5.472199, 5.499791, 5.508503, 5.496091, 
    5.462376, 5.409999, 5.344549, 5.273689, 5.205394, 5.146018, 5.099126, 
    5.065478,
  // totalHeight(7,40, 0-49)
    5.01671, 5.028383, 5.047037, 5.074806, 5.113331, 5.162851, 5.22134, 
    5.284199, 5.344914, 5.396571, 5.433529, 5.452536, 5.452931, 5.436152, 
    5.404949, 5.367265, 5.35313, 5.307418, 5.259766, 5.2129, 5.167883, 
    5.131764, 5.097353, 5.067103, 5.04221, 5.024868, 5.016986, 5.020291, 
    5.035318, 5.062237, 5.098837, 5.149593, 5.206281, 5.266251, 5.326477, 
    5.383618, 5.434089, 5.474142, 5.500051, 5.508503, 5.497226, 5.465776, 
    5.416249, 5.353471, 5.28436, 5.216414, 5.155935, 5.106784, 5.070136, 
    5.045145,
  // totalHeight(7,41, 0-49)
    5.011393, 5.019699, 5.033443, 5.054687, 5.08547, 5.127131, 5.179427, 
    5.239829, 5.303455, 5.363914, 5.414792, 5.451157, 5.470404, 5.472347, 
    5.458686, 5.435668, 5.427438, 5.390626, 5.348041, 5.302955, 5.257243, 
    5.218533, 5.181604, 5.149585, 5.123898, 5.107349, 5.101637, 5.107809, 
    5.125257, 5.153823, 5.190883, 5.239744, 5.292246, 5.345578, 5.396583, 
    5.44182, 5.477694, 5.500643, 5.507504, 5.496064, 5.465759, 5.418307, 
    5.357935, 5.290864, 5.224049, 5.163566, 5.113376, 5.074951, 5.047723, 
    5.029982,
  // totalHeight(7,42, 0-49)
    5.007448, 5.013103, 5.022773, 5.03824, 5.061559, 5.094617, 5.138445, 
    5.192428, 5.253744, 5.317492, 5.377594, 5.428209, 5.465016, 5.485915, 
    5.491031, 5.484582, 5.484806, 5.458848, 5.423669, 5.382972, 5.339408, 
    5.300989, 5.264325, 5.232959, 5.208259, 5.193301, 5.189502, 5.197357, 
    5.215441, 5.243477, 5.278582, 5.322964, 5.368637, 5.412613, 5.451626, 
    5.482244, 5.501094, 5.50519, 5.492446, 5.462286, 5.416188, 5.357902, 
    5.293029, 5.227933, 5.168333, 5.118133, 5.078968, 5.050518, 5.031245, 
    5.019185,
  // totalHeight(7,43, 0-49)
    5.004671, 5.00836, 5.014862, 5.025596, 5.042367, 5.06715, 5.101645, 
    5.146619, 5.201205, 5.262506, 5.325803, 5.385471, 5.436242, 5.474329, 
    5.498009, 5.509168, 5.520347, 5.507353, 5.482279, 5.449014, 5.41083, 
    5.375861, 5.342307, 5.313881, 5.291713, 5.278893, 5.276544, 5.284764, 
    5.301612, 5.326838, 5.35743, 5.394591, 5.430645, 5.462481, 5.486856, 
    5.500595, 5.500926, 5.485937, 5.455106, 5.409778, 5.353324, 5.290773, 
    5.22789, 5.169929, 5.120594, 5.081575, 5.05273, 5.03272, 5.019693, 
    5.011834,
  // totalHeight(7,44, 0-49)
    5.002813, 5.005119, 5.009302, 5.016413, 5.027887, 5.045482, 5.071043, 
    5.106079, 5.151144, 5.205262, 5.265625, 5.327862, 5.386883, 5.437991, 
    5.477863, 5.506032, 5.529777, 5.531497, 5.519186, 5.496544, 5.467158, 
    5.438933, 5.411334, 5.388013, 5.36974, 5.359428, 5.357933, 5.365097, 
    5.378753, 5.398783, 5.422194, 5.449341, 5.473051, 5.490255, 5.498004, 
    5.493757, 5.475805, 5.443734, 5.398806, 5.344073, 5.284039, 5.223843, 
    5.168211, 5.120537, 5.082442, 5.053911, 5.033787, 5.020379, 5.011954, 
    5.007036,
  // totalHeight(7,45, 0-49)
    5.001627, 5.00301, 5.005588, 5.010087, 5.017568, 5.029425, 5.047313, 
    5.072919, 5.10756, 5.151648, 5.204203, 5.262649, 5.32308, 5.380993, 
    5.432267, 5.474555, 5.510695, 5.527712, 5.530097, 5.520863, 5.503451, 
    5.485116, 5.466168, 5.449955, 5.436787, 5.429237, 5.42793, 5.432586, 
    5.441073, 5.453529, 5.467171, 5.481771, 5.49093, 5.491922, 5.482465, 
    5.461075, 5.427461, 5.382823, 5.329916, 5.272722, 5.215748, 5.163129, 
    5.11786, 5.081418, 5.053839, 5.034134, 5.020792, 5.012212, 5.00699, 
    5.004033,
  // totalHeight(7,46, 0-49)
    5.000904, 5.001698, 5.003219, 5.005941, 5.01059, 5.018181, 5.030026, 
    5.047634, 5.072513, 5.105799, 5.147814, 5.197673, 5.25313, 5.310821, 
    5.366889, 5.418075, 5.464053, 5.494967, 5.512374, 5.518117, 5.514961, 
    5.509031, 5.500986, 5.493574, 5.486524, 5.481907, 5.480128, 5.480912, 
    5.48242, 5.485212, 5.486995, 5.487328, 5.480935, 5.465807, 5.440713, 
    5.405491, 5.361278, 5.310514, 5.256648, 5.203514, 5.154617, 5.112494, 
    5.078404, 5.052387, 5.033595, 5.020703, 5.01228, 5.007036, 5.003934, 
    5.002227,
  // totalHeight(7,47, 0-49)
    5.000479, 5.000916, 5.001769, 5.003335, 5.006079, 5.010685, 5.018091, 
    5.029477, 5.046185, 5.069523, 5.100471, 5.139313, 5.185328, 5.236683, 
    5.29062, 5.344086, 5.395159, 5.436237, 5.466683, 5.48693, 5.498612, 
    5.506318, 5.510494, 5.51297, 5.512695, 5.511067, 5.508265, 5.504123, 
    5.497348, 5.489172, 5.47811, 5.463986, 5.442956, 5.414068, 5.377319, 
    5.333785, 5.285583, 5.235593, 5.186958, 5.142507, 5.104268, 5.07323, 
    5.049392, 5.032015, 5.019961, 5.011981, 5.006932, 5.003879, 5.00212, 
    5.001179,
  // totalHeight(7,48, 0-49)
    5.000237, 5.00046, 5.000906, 5.001745, 5.003255, 5.005858, 5.010167, 
    5.017009, 5.027408, 5.04252, 5.063472, 5.091123, 5.125785, 5.16698, 
    5.213346, 5.262811, 5.313305, 5.359091, 5.398305, 5.430139, 5.45493, 
    5.475578, 5.491802, 5.50423, 5.510761, 5.511994, 5.507837, 5.49834, 
    5.482945, 5.46386, 5.440705, 5.414022, 5.381519, 5.343398, 5.300726, 
    5.255343, 5.209594, 5.165942, 5.126526, 5.092831, 5.06552, 5.044494, 
    5.029083, 5.018308, 5.011105, 5.006493, 5.003665, 5.002002, 5.00107, 
    5.000583,
  // totalHeight(7,49, 0-49)
    5.000078, 5.000158, 5.000323, 5.000648, 5.001265, 5.002378, 5.004317, 
    5.007565, 5.012781, 5.020815, 5.032668, 5.049388, 5.071904, 5.100811, 
    5.136148, 5.177304, 5.223419, 5.26947, 5.313471, 5.353898, 5.39002, 
    5.424407, 5.454918, 5.480593, 5.49589, 5.500593, 5.494115, 5.476953, 
    5.449314, 5.416775, 5.380487, 5.34278, 5.30167, 5.258408, 5.214767, 
    5.172745, 5.1342, 5.100561, 5.072627, 5.050539, 5.033884, 5.021892, 
    5.013636, 5.008191, 5.004746, 5.002652, 5.001432, 5.00075, 5.000383, 
    5.000201,
  // totalHeight(8,0, 0-49)
    5.001369, 5.00236, 5.004135, 5.007111, 5.011874, 5.019187, 5.02997, 
    5.045208, 5.065813, 5.092411, 5.125103, 5.163265, 5.205472, 5.249606, 
    5.293155, 5.333694, 5.369721, 5.397316, 5.416229, 5.42692, 5.430637, 
    5.429839, 5.425939, 5.420931, 5.415915, 5.412307, 5.410614, 5.410615, 
    5.41119, 5.411488, 5.409767, 5.404738, 5.39423, 5.377171, 5.353137, 
    5.322467, 5.286308, 5.246513, 5.205389, 5.165338, 5.128472, 5.096318, 
    5.069674, 5.048647, 5.032804, 5.021383, 5.013495, 5.008281, 5.005001, 
    5.003084,
  // totalHeight(8,1, 0-49)
    5.002229, 5.003803, 5.006566, 5.011106, 5.018226, 5.028921, 5.044301, 
    5.065442, 5.093146, 5.127659, 5.168413, 5.213895, 5.261753, 5.309123, 
    5.353121, 5.391528, 5.424201, 5.445468, 5.456513, 5.458668, 5.453891, 
    5.445782, 5.435674, 5.425931, 5.417472, 5.412071, 5.410341, 5.412109, 
    5.416037, 5.421542, 5.426564, 5.429821, 5.428074, 5.419613, 5.403261, 
    5.378569, 5.345982, 5.306887, 5.263489, 5.218513, 5.174774, 5.134702, 
    5.100015, 5.071559, 5.049369, 5.032875, 5.021171, 5.013241, 5.008139, 
    5.005085,
  // totalHeight(8,2, 0-49)
    5.003713, 5.006243, 5.010573, 5.017516, 5.028118, 5.043579, 5.065092, 
    5.093582, 5.12938, 5.171907, 5.219525, 5.269629, 5.319023, 5.3645, 
    5.403409, 5.434417, 5.459604, 5.47129, 5.472511, 5.465329, 5.452096, 
    5.437172, 5.421472, 5.407487, 5.395916, 5.388781, 5.386798, 5.389922, 
    5.39677, 5.407083, 5.418703, 5.430604, 5.438771, 5.441057, 5.435635, 
    5.421216, 5.397282, 5.364281, 5.323711, 5.278013, 5.230247, 5.183597, 
    5.140839, 5.103923, 5.073798, 5.050491, 5.033351, 5.021364, 5.013425, 
    5.008539,
  // totalHeight(8,3, 0-49)
    5.006076, 5.010056, 5.016683, 5.027022, 5.042336, 5.063916, 5.092799, 
    5.129389, 5.173098, 5.222139, 5.273632, 5.324032, 5.36979, 5.408006, 
    5.436888, 5.456504, 5.471837, 5.472431, 5.463517, 5.447612, 5.427128, 
    5.40682, 5.386859, 5.369648, 5.355633, 5.346969, 5.344492, 5.348353, 
    5.357283, 5.371386, 5.388593, 5.408371, 5.426187, 5.439701, 5.446662, 
    5.445097, 5.433551, 5.411355, 5.378881, 5.337667, 5.290347, 5.24031, 
    5.191145, 5.146004, 5.107107, 5.075537, 5.051323, 5.033752, 5.021726, 
    5.014085,
  // totalHeight(8,4, 0-49)
    5.009637, 5.015692, 5.025481, 5.040294, 5.061502, 5.09025, 5.127049, 
    5.171336, 5.221224, 5.273581, 5.324505, 5.370071, 5.407087, 5.433594, 
    5.449055, 5.455122, 5.460109, 5.449643, 5.431532, 5.408463, 5.382619, 
    5.358882, 5.336395, 5.317299, 5.301744, 5.291907, 5.288743, 5.292657, 
    5.302639, 5.319189, 5.340461, 5.366611, 5.392787, 5.416655, 5.435787, 
    5.447778, 5.450466, 5.442185, 5.42209, 5.39045, 5.348847, 5.300132, 
    5.24806, 5.196651, 5.149448, 5.108942, 5.07633, 5.051642, 5.034104, 
    5.022564,
  // totalHeight(8,5, 0-49)
    5.01475, 5.023616, 5.037497, 5.057807, 5.085801, 5.12212, 5.166306, 
    5.216456, 5.269265, 5.320505, 5.365861, 5.401783, 5.426079, 5.438101, 
    5.438597, 5.430701, 5.42629, 5.4058, 5.380095, 5.351824, 5.322756, 
    5.297715, 5.274599, 5.255134, 5.239125, 5.228632, 5.224696, 5.228026, 
    5.237998, 5.255537, 5.279135, 5.309788, 5.342454, 5.374955, 5.404862, 
    5.429592, 5.446565, 5.453413, 5.448264, 5.430104, 5.399138, 5.357038, 
    5.306925, 5.252957, 5.199602, 5.15078, 5.109215, 5.07619, 5.051716, 
    5.034968,
  // totalHeight(8,6, 0-49)
    5.021751, 5.034218, 5.053062, 5.079626, 5.114713, 5.158042, 5.207815, 
    5.260664, 5.312117, 5.35747, 5.39277, 5.415498, 5.424806, 5.421356, 
    5.406937, 5.385913, 5.373868, 5.3448, 5.313278, 5.281764, 5.251529, 
    5.227237, 5.205383, 5.187147, 5.171925, 5.161469, 5.156841, 5.159067, 
    5.168033, 5.185125, 5.209272, 5.242446, 5.279513, 5.318528, 5.357177, 
    5.392874, 5.422873, 5.444416, 5.454944, 5.452408, 5.435674, 5.404944, 
    5.362053, 5.310448, 5.254735, 5.199829, 5.15, 5.108155, 5.075609, 5.052327,
  // totalHeight(8,7, 0-49)
    5.03087, 5.047679, 5.07213, 5.105202, 5.146861, 5.19554, 5.247961, 
    5.299513, 5.345158, 5.38049, 5.402569, 5.410242, 5.403994, 5.385534, 
    5.357308, 5.324667, 5.306974, 5.270771, 5.235045, 5.202008, 5.172415, 
    5.150715, 5.131906, 5.116521, 5.103456, 5.093926, 5.088892, 5.089666, 
    5.096759, 5.112054, 5.135026, 5.168761, 5.208121, 5.251438, 5.296572, 
    5.341026, 5.38205, 5.416742, 5.442186, 5.45566, 5.454984, 5.438967, 
    5.407883, 5.363819, 5.310629, 5.253408, 5.197519, 5.147527, 5.106443, 
    5.075536,
  // totalHeight(8,8, 0-49)
    5.042141, 5.063857, 5.094147, 5.13329, 5.180078, 5.231492, 5.282947, 
    5.329145, 5.365218, 5.387711, 5.395039, 5.387403, 5.366355, 5.334259, 
    5.293848, 5.251297, 5.229727, 5.187588, 5.148976, 5.115803, 5.088339, 
    5.070806, 5.056664, 5.045733, 5.036299, 5.028781, 5.023865, 5.023066, 
    5.027584, 5.039847, 5.060001, 5.092403, 5.132013, 5.177479, 5.226856, 
    5.277767, 5.32753, 5.373251, 5.411896, 5.440407, 5.455941, 5.456232, 
    5.440107, 5.408016, 5.362398, 5.307615, 5.249297, 5.193226, 5.14417, 
    5.105097,
  // totalHeight(8,9, 0-49)
    5.055322, 5.08219, 5.118004, 5.162039, 5.21173, 5.262723, 5.309602, 
    5.347069, 5.371074, 5.379469, 5.372033, 5.35006, 5.315778, 5.271844, 
    5.22097, 5.170115, 5.145872, 5.098701, 5.058197, 5.025952, 5.0018, 
    4.989735, 4.981704, 4.976761, 4.972498, 4.968266, 4.964252, 4.962024, 
    4.963476, 4.971612, 4.987387, 5.016612, 5.05449, 5.100041, 5.151529, 
    5.206686, 5.262909, 5.317366, 5.367041, 5.408783, 5.439424, 5.456029, 
    5.456311, 5.439203, 5.405454, 5.357993, 5.301782, 5.243008, 5.187781, 
    5.140861,
  // totalHeight(8,10, 0-49)
    5.069841, 5.101693, 5.142138, 5.189268, 5.239218, 5.286673, 5.326009, 
    5.352551, 5.363453, 5.357918, 5.336849, 5.30226, 5.256696, 5.202795, 
    5.143048, 5.085224, 5.058656, 5.007109, 4.965445, 4.934928, 4.915015, 
    4.909478, 4.908812, 4.911294, 4.913756, 4.914239, 4.912184, 4.908985, 
    4.907153, 4.910244, 4.920147, 4.944366, 4.97854, 5.022159, 5.07372, 
    5.131052, 5.191589, 5.252552, 5.310984, 5.363772, 5.407672, 5.439425, 
    5.456047, 5.4553, 5.436343, 5.400368, 5.35093, 5.293661, 5.235225, 
    5.181823,
  // totalHeight(8,11, 0-49)
    5.084838, 5.121063, 5.164775, 5.212887, 5.260504, 5.301888, 5.331789, 
    5.346568, 5.34467, 5.326456, 5.293612, 5.248514, 5.193708, 5.13161, 
    5.064352, 5.000533, 4.970798, 4.915408, 4.873148, 4.844985, 4.83006, 
    4.831906, 4.839677, 4.850883, 4.861561, 4.868284, 4.869509, 4.866175, 
    4.861197, 4.858579, 4.861226, 4.878594, 4.907023, 4.946648, 4.996276, 
    5.053806, 5.116663, 5.182054, 5.247064, 5.308654, 5.363636, 5.408683, 
    5.44047, 5.45601, 5.453212, 5.431593, 5.392934, 5.341518, 5.283602, 
    5.226091,
  // totalHeight(8,12, 0-49)
    5.099267, 5.138888, 5.184268, 5.231308, 5.274516, 5.308251, 5.328059, 
    5.331479, 5.318122, 5.289199, 5.246833, 5.19346, 5.131418, 5.062748, 
    4.989133, 4.919843, 4.884488, 4.825829, 4.783488, 4.758223, 4.748928, 
    4.758839, 4.775925, 4.796943, 4.817178, 4.831673, 4.837736, 4.835538, 
    4.828052, 4.819459, 4.813668, 4.822335, 4.842855, 4.876289, 4.92189, 
    4.977654, 5.040928, 5.108822, 5.178389, 5.246644, 5.310491, 5.366675, 
    5.411796, 5.442484, 5.455814, 5.449941, 5.424872, 5.383087, 5.32959, 
    5.271071,
  // totalHeight(8,13, 0-49)
    5.112081, 5.153917, 5.199409, 5.243758, 5.281303, 5.306915, 5.317125, 
    5.310584, 5.287816, 5.250561, 5.201094, 5.141697, 5.07436, 5.000659, 
    4.921747, 4.846888, 4.801401, 4.740222, 4.698379, 4.676562, 4.673483, 
    4.691962, 4.719002, 4.750622, 4.781459, 4.80514, 4.817774, 4.818466, 
    4.809773, 4.795585, 4.780596, 4.77881, 4.789131, 4.813954, 4.853247, 
    4.905177, 4.966969, 5.035536, 5.107794, 5.180731, 5.25133, 5.316455, 
    5.372781, 5.41683, 5.445218, 5.455135, 5.445074, 5.415627, 5.37001, 
    5.313847,
  // totalHeight(8,14, 0-49)
    5.122416, 5.165294, 5.209671, 5.250387, 5.28198, 5.300036, 5.302077, 
    5.287667, 5.25795, 5.214927, 5.160814, 5.097618, 5.026911, 4.949761, 
    4.8667, 4.785186, 4.722669, 4.659978, 4.619365, 4.601606, 4.605288, 
    4.632604, 4.669907, 4.712483, 4.754512, 4.788497, 4.809477, 4.815284, 
    4.807504, 4.789055, 4.764913, 4.75128, 4.749103, 4.762674, 4.793109, 
    4.838937, 4.897255, 4.964674, 5.037851, 5.11364, 5.18903, 5.260995, 
    5.326344, 5.381658, 5.423375, 5.448099, 5.453174, 5.437504, 5.402347, 
    5.351675,
  // totalHeight(8,15, 0-49)
    5.129766, 5.172712, 5.215269, 5.252206, 5.278469, 5.290407, 5.286373, 
    5.266594, 5.232567, 5.18635, 5.129982, 5.065152, 4.993019, 4.914148, 
    4.828405, 4.73751, 4.64882, 4.585863, 4.547379, 4.534361, 4.545287, 
    4.581367, 4.628794, 4.682116, 4.735318, 4.780255, 4.811194, 4.824649, 
    4.820728, 4.800571, 4.768612, 4.74255, 4.725894, 4.725502, 4.744281, 
    4.781486, 4.83417, 4.898561, 4.970917, 5.047832, 5.126202, 5.203052, 
    5.275322, 5.339731, 5.392716, 5.430585, 5.449921, 5.448276, 5.425073, 
    5.382407,
  // totalHeight(8,16, 0-49)
    5.134052, 5.176439, 5.217067, 5.250836, 5.273164, 5.281045, 5.27343, 
    5.250941, 5.215213, 5.16822, 5.111789, 5.047322, 4.975654, 4.896925, 
    4.81037, 4.704902, 4.579583, 4.517775, 4.48243, 4.474857, 4.49339, 
    4.537728, 4.59462, 4.65787, 4.721575, 4.777524, 4.819635, 4.843246, 
    4.846655, 4.828532, 4.791764, 4.754059, 4.721835, 4.705099, 4.70937, 
    4.735244, 4.779961, 4.839344, 4.909132, 4.985513, 5.065176, 5.145107, 
    5.222342, 5.293738, 5.355831, 5.404837, 5.436883, 5.448555, 5.437765, 
    5.404779,
  // totalHeight(8,17, 0-49)
    5.13558, 5.177178, 5.216339, 5.248187, 5.268536, 5.274807, 5.266268, 
    5.243672, 5.208608, 5.162899, 5.108179, 5.045659, 4.975985, 4.899038, 
    4.813493, 4.685416, 4.513347, 4.454445, 4.423234, 4.421718, 4.448077, 
    4.499756, 4.565007, 4.636907, 4.70996, 4.776448, 4.830373, 4.866174, 
    4.880282, 4.868591, 4.831599, 4.784774, 4.737452, 4.702971, 4.690291, 
    4.702183, 4.736541, 4.78889, 4.854359, 4.928604, 5.007979, 5.08934, 
    5.169746, 5.246167, 5.315263, 5.37328, 5.416127, 5.43977, 5.440993, 
    5.418493,
  // totalHeight(8,18, 0-49)
    5.134904, 5.175833, 5.214426, 5.246045, 5.266733, 5.274041, 5.267223, 
    5.246889, 5.214422, 5.171445, 5.119457, 5.059613, 4.99252, 4.917845, 
    4.833514, 4.673349, 4.446044, 4.392892, 4.366827, 4.371818, 4.406159, 
    4.46414, 4.53652, 4.615712, 4.696862, 4.773158, 4.838974, 4.888155, 
    4.915483, 4.914273, 4.88238, 4.830496, 4.7705, 4.718554, 4.687547, 
    4.683339, 4.705169, 4.748554, 4.808033, 4.878636, 4.956275, 5.037578, 
    5.119546, 5.199218, 5.273369, 5.338331, 5.389959, 5.423878, 5.43611, 
    5.42413,
  // totalHeight(8,19, 0-49)
    5.132595, 5.173156, 5.21232, 5.245671, 5.269256, 5.280378, 5.277858, 
    5.261819, 5.23324, 5.193517, 5.144123, 5.086297, 5.020607, 4.946133, 
    4.858912, 4.659686, 4.369835, 4.327592, 4.308208, 4.320153, 4.362873, 
    4.426592, 4.505294, 4.590879, 4.679287, 4.764817, 4.84228, 4.905135, 
    4.946831, 4.958759, 4.936626, 4.884299, 4.815693, 4.74858, 4.699572, 
    4.678265, 4.686046, 4.71891, 4.770968, 4.836618, 4.91126, 4.991214, 
    5.073359, 5.154741, 5.232225, 5.30225, 5.360712, 5.4031, 5.424982, 
    5.422957,
  // totalHeight(8,20, 0-49)
    5.126199, 5.16312, 5.199585, 5.231456, 5.255075, 5.268044, 5.269554, 
    5.260229, 5.241733, 5.216325, 5.186499, 5.154742, 5.123319, 5.093983, 
    5.067405, 30, 4.110707, 4.123703, 4.162252, 4.22343, 4.302578, 4.387699, 
    4.480834, 4.576489, 4.673163, 4.767192, 4.854263, 4.927924, 4.980938, 
    5.003913, 4.991771, 4.940973, 4.867107, 4.788014, 4.72289, 4.684924, 
    4.678152, 4.699588, 4.743227, 4.802933, 4.873587, 4.951164, 5.032368, 
    5.114204, 5.193589, 5.267064, 5.330619, 5.379736, 5.409759, 5.416706,
  // totalHeight(8,21, 0-49)
    5.123293, 5.160292, 5.19839, 5.233569, 5.261959, 5.280674, 5.288291, 
    5.284894, 5.271763, 5.25098, 5.225037, 5.196559, 5.168098, 5.141923, 
    5.119676, 30, 4.030297, 4.047019, 4.093606, 4.164876, 4.254046, 4.343937, 
    4.441362, 4.540665, 4.641256, 4.74086, 4.835884, 4.920084, 4.985749, 
    5.023064, 5.026696, 4.98524, 4.915319, 4.832731, 4.757448, 4.705839, 
    4.685367, 4.695097, 4.729599, 4.782505, 4.848262, 4.922476, 5.001632, 
    5.082644, 5.162446, 5.237658, 5.304375, 5.358139, 5.394198, 5.408191,
  // totalHeight(8,22, 0-49)
    5.121522, 5.158882, 5.19856, 5.236558, 5.268754, 5.291821, 5.30385, 
    5.304541, 5.29497, 5.277183, 5.253765, 5.227507, 5.201188, 5.177412, 
    5.158434, 30, 3.962537, 3.984438, 4.038232, 4.117738, 4.215069, 4.308348, 
    4.409274, 4.511858, 4.616008, 4.720365, 4.821665, 4.913651, 4.988194, 
    5.035557, 5.051208, 5.016985, 4.95165, 4.868662, 4.787441, 4.726087, 
    4.694775, 4.694649, 4.721154, 4.767963, 4.829233, 4.900268, 4.97734, 
    5.057264, 5.136958, 5.2131, 5.281876, 5.338915, 5.379454, 5.398909,
  // totalHeight(8,23, 0-49)
    5.120916, 5.158588, 5.199337, 5.239162, 5.273767, 5.299524, 5.314222, 
    5.31733, 5.309831, 5.293787, 5.271873, 5.247006, 5.222109, 5.199984, 
    5.183231, 30, 3.917093, 3.943388, 4.002137, 4.086914, 4.189435, 4.283938, 
    4.386425, 4.49054, 4.59648, 4.703573, 4.808774, 4.905783, 4.986151, 
    5.040359, 5.064946, 5.036311, 4.975649, 4.894337, 4.810658, 4.743364, 
    4.704498, 4.696982, 4.71723, 4.759143, 4.816749, 4.885137, 4.960407, 
    5.039274, 5.118623, 5.195158, 5.265129, 5.324236, 5.367732, 5.390903,
  // totalHeight(8,24, 0-49)
    5.121484, 5.15919, 5.200179, 5.240473, 5.275757, 5.302342, 5.317935, 
    5.321938, 5.315293, 5.30006, 5.278937, 5.254865, 5.230805, 5.209631, 
    5.194072, 30, 3.898081, 3.926662, 3.987599, 4.074533, 4.179204, 4.273223, 
    4.375597, 4.479658, 4.58575, 4.69365, 4.800478, 4.89992, 4.983319, 
    5.04135, 5.071414, 5.046269, 4.989053, 4.909707, 4.825484, 4.755218, 
    4.711973, 4.699844, 4.715989, 4.754571, 4.8096, 4.876063, 4.949962, 
    5.027952, 5.106898, 5.183519, 5.254107, 5.31441, 5.359709, 5.385231,
  // totalHeight(8,25, 0-49)
    5.12319, 5.160546, 5.200797, 5.240048, 5.274151, 5.299625, 5.314344, 
    5.317798, 5.31093, 5.295742, 5.274842, 5.251086, 5.227356, 5.206459, 
    5.191058, 30, 3.905595, 3.934001, 3.99451, 4.080811, 4.184822, 4.277218, 
    4.378278, 4.481149, 4.586186, 4.693312, 4.799687, 4.89899, 4.982497, 
    5.040989, 5.072271, 5.047817, 4.991623, 4.913149, 4.829183, 4.758409, 
    4.714091, 4.70067, 4.715574, 4.753094, 4.807269, 4.873075, 4.946495, 
    5.024164, 5.102949, 5.179572, 5.250342, 5.311027, 5.356915, 5.383218,
  // totalHeight(8,26, 0-49)
    5.125965, 5.16261, 5.201203, 5.237979, 5.269135, 5.291635, 5.303749, 
    5.305204, 5.296997, 5.28103, 5.259737, 5.235774, 5.211836, 5.190529, 
    5.174261, 30, 3.937386, 3.963501, 4.021425, 4.104737, 4.20558, 4.295581, 
    4.394385, 4.495152, 4.598157, 4.703125, 4.807133, 4.903847, 4.984638, 
    5.040278, 5.0684, 5.04177, 4.983876, 4.904703, 4.821317, 4.752176, 
    4.709991, 4.698662, 4.715331, 4.75422, 4.809419, 4.87597, 4.949917, 
    5.027929, 5.106887, 5.183514, 5.254105, 5.314409, 5.359708, 5.385231,
  // totalHeight(8,27, 0-49)
    5.129717, 5.165435, 5.201689, 5.23486, 5.261594, 5.279465, 5.287314, 
    5.285252, 5.274403, 5.256595, 5.234052, 5.209174, 5.184377, 5.16194, 
    5.143804, 30, 3.989284, 4.01185, 4.065571, 4.143941, 4.239443, 4.326462, 
    4.422174, 4.519982, 4.619985, 4.72141, 4.821146, 4.912863, 4.98817, 
    5.037752, 5.058598, 5.027196, 4.965382, 4.884583, 4.802653, 4.737598, 
    4.700779, 4.694783, 4.716008, 4.758492, 4.81641, 4.884964, 4.96032, 
    5.03923, 5.118601, 5.195146, 5.265124, 5.324234, 5.36773, 5.390903,
  // totalHeight(8,28, 0-49)
    5.134365, 5.169187, 5.202791, 5.231663, 5.252913, 5.264796, 5.266833, 
    5.25964, 5.244601, 5.223562, 5.198596, 5.171845, 5.145388, 5.121049, 
    5.100052, 30, 4.056873, 4.075941, 4.124346, 4.195992, 4.284093, 4.367258, 
    4.458745, 4.55243, 4.648153, 4.744445, 4.837958, 4.922404, 4.989758, 
    5.030591, 5.041007, 5.003144, 4.936561, 4.854705, 4.776264, 4.7182, 
    4.689766, 4.691714, 4.719532, 4.767098, 4.828782, 4.900036, 4.977222, 
    5.057204, 5.136929, 5.213084, 5.281867, 5.338911, 5.379453, 5.398908,
  // totalHeight(8,29, 0-49)
    5.139871, 5.174164, 5.205247, 5.229603, 5.244735, 5.249564, 5.244349, 
    5.230343, 5.209353, 5.183419, 5.154596, 5.124834, 5.095839, 5.068839, 
    5.043989, 30, 4.134919, 4.152247, 4.194923, 4.258248, 4.336938, 4.414831, 
    4.500596, 4.588754, 4.67878, 4.768302, 4.853632, 4.928486, 4.985303, 
    5.014688, 5.012098, 4.966738, 4.896005, 4.815494, 4.744064, 4.696627, 
    4.679617, 4.691761, 4.727758, 4.781523, 4.847747, 4.922211, 5.001495, 
    5.082574, 5.16241, 5.23764, 5.304365, 5.358133, 5.394195, 5.408189,
  // totalHeight(8,30, 0-49)
    5.149293, 5.187366, 5.220729, 5.245617, 5.259345, 5.260664, 5.249608, 
    5.227057, 5.194283, 5.152627, 5.103288, 5.047123, 4.984291, 4.913467, 
    4.830404, 4.635087, 4.366791, 4.33845, 4.330659, 4.350416, 4.397135, 
    4.457949, 4.533136, 4.614896, 4.700094, 4.78401, 4.861721, 4.926516, 
    4.971288, 4.987126, 4.969789, 4.916682, 4.843794, 4.76844, 4.708371, 
    4.675247, 4.67223, 4.696182, 4.74135, 4.801925, 4.873054, 4.950885, 
    5.032222, 5.114128, 5.19355, 5.267044, 5.330608, 5.37973, 5.409755, 
    5.416704,
  // totalHeight(8,31, 0-49)
    5.154108, 5.192601, 5.225134, 5.247748, 5.25784, 5.254495, 5.238242, 
    5.21049, 5.172945, 5.127208, 5.074561, 5.015869, 4.951433, 4.880641, 
    4.801196, 4.644937, 4.432422, 4.392949, 4.379121, 4.393623, 4.43407, 
    4.491832, 4.56249, 4.638905, 4.717442, 4.792549, 4.859183, 4.911111, 
    4.942367, 4.945229, 4.916481, 4.861229, 4.793419, 4.729975, 4.685867, 
    4.669163, 4.680465, 4.715677, 4.769167, 4.835639, 4.910736, 4.990936, 
    5.073214, 5.154664, 5.232185, 5.30223, 5.360701, 5.403094, 5.424978, 
    5.422956,
  // totalHeight(8,32, 0-49)
    5.157407, 5.197023, 5.230282, 5.252917, 5.262111, 5.256892, 5.237898, 
    5.206759, 5.165463, 5.115866, 5.059437, 4.997152, 4.929425, 4.855934, 
    4.775219, 4.651386, 4.489683, 4.443143, 4.423618, 4.431955, 4.465497, 
    4.519353, 4.584921, 4.655719, 4.727498, 4.793783, 4.849238, 4.888139, 
    4.905953, 4.896959, 4.860013, 4.806783, 4.748804, 4.70111, 4.675007, 
    4.67511, 4.700132, 4.745621, 4.806382, 4.877728, 4.955783, 5.037313, 
    5.119405, 5.199143, 5.273329, 5.33831, 5.389947, 5.423872, 5.436106, 
    5.424129,
  // totalHeight(8,33, 0-49)
    5.158516, 5.199754, 5.23505, 5.259749, 5.270575, 5.266178, 5.24701, 
    5.214706, 5.171402, 5.119178, 5.05975, 4.994316, 4.923507, 4.847308, 
    4.764863, 4.663693, 4.545833, 4.494422, 4.469296, 4.470886, 4.496832, 
    4.54519, 4.604345, 4.668429, 4.732591, 4.78956, 4.833763, 4.860198, 
    4.866086, 4.848289, 4.808124, 4.76158, 4.717298, 4.687345, 4.679305, 
    4.695044, 4.732172, 4.786329, 4.852901, 4.927793, 5.007535, 5.089099, 
    5.169616, 5.246097, 5.315227, 5.37326, 5.416117, 5.439764, 5.44099, 
    5.418491,
  // totalHeight(8,34, 0-49)
    5.156674, 5.199654, 5.237898, 5.26634, 5.281066, 5.280095, 5.263408, 
    5.232435, 5.189331, 5.136365, 5.075525, 5.008317, 4.935713, 4.858127, 
    4.77535, 4.688264, 4.605028, 4.550157, 4.519898, 4.514716, 4.532631, 
    4.573838, 4.625031, 4.68093, 4.736253, 4.78332, 4.816595, 4.832085, 
    4.828914, 4.806611, 4.768563, 4.732501, 4.703937, 4.691649, 4.700083, 
    4.72925, 4.776286, 4.837176, 4.907887, 4.984814, 5.064787, 5.144894, 
    5.222227, 5.293676, 5.355797, 5.404819, 5.436873, 5.448549, 5.437762, 
    5.404777,
  // totalHeight(8,35, 0-49)
    5.151281, 5.195655, 5.237204, 5.270538, 5.291034, 5.29586, 5.284276, 
    5.257265, 5.216847, 5.165399, 5.10517, 5.038023, 4.965342, 4.888039, 
    4.806555, 4.727874, 4.66922, 4.612257, 4.577751, 4.566242, 4.576077, 
    4.608909, 4.650864, 4.69726, 4.742668, 4.779547, 4.802795, 4.809654, 
    4.800983, 4.778551, 4.746922, 4.72342, 4.710607, 4.714301, 4.736648, 
    4.776581, 4.831155, 4.89677, 4.969879, 5.047243, 5.125873, 5.202868, 
    5.275223, 5.339676, 5.392687, 5.430571, 5.449914, 5.448271, 5.425071, 
    5.382406,
  // totalHeight(8,36, 0-49)
    5.142104, 5.187049, 5.231609, 5.270293, 5.297827, 5.310411, 5.306343, 
    5.285905, 5.250766, 5.203276, 5.145887, 5.080808, 5.009852, 4.934427, 
    4.85556, 4.782229, 4.739129, 4.681488, 4.643786, 4.626654, 4.628716, 
    4.652565, 4.684572, 4.720676, 4.75562, 4.782554, 4.797193, 4.798059, 
    4.787327, 4.768233, 4.745573, 4.734941, 4.736442, 4.753576, 4.786968, 
    4.834998, 4.894826, 4.963222, 5.037002, 5.113153, 5.188756, 5.260842, 
    5.326259, 5.381612, 5.423351, 5.448085, 5.453167, 5.4375, 5.402345, 
    5.351675,
  // totalHeight(8,37, 0-49)
    5.129393, 5.173698, 5.220318, 5.263993, 5.299031, 5.320687, 5.326133, 
    5.314678, 5.287379, 5.246348, 5.194114, 5.133163, 5.065706, 4.993609, 
    4.918402, 4.849136, 4.814672, 4.757637, 4.717738, 4.695762, 4.690593, 
    4.705426, 4.727391, 4.753076, 4.777669, 4.795451, 4.803186, 4.800547, 
    4.790458, 4.776838, 4.763995, 4.765265, 4.778885, 4.806695, 4.848376, 
    4.902049, 4.965028, 5.034365, 5.107103, 5.18033, 5.251101, 5.316327, 
    5.372707, 5.41679, 5.445196, 5.455124, 5.445068, 5.415625, 5.370009, 
    5.313847,
  // totalHeight(8,38, 0-49)
    5.113876, 5.156118, 5.203286, 5.250753, 5.292802, 5.323964, 5.340252, 
    5.339784, 5.322693, 5.290582, 5.245847, 5.191123, 5.128939, 5.06156, 
    4.990949, 4.92551, 4.895123, 4.839703, 4.798448, 4.772382, 4.760661, 
    4.766866, 4.779205, 4.794943, 4.809895, 4.819722, 4.822293, 4.81818, 
    4.810492, 4.803233, 4.799835, 4.811351, 4.83469, 4.870549, 4.918038, 
    4.975163, 5.039362, 5.107861, 5.17781, 5.2463, 5.31029, 5.36656, 
    5.411729, 5.442446, 5.455794, 5.449931, 5.424867, 5.383084, 5.329588, 
    5.27107,
  // totalHeight(8,39, 0-49)
    5.096656, 5.135428, 5.181291, 5.230628, 5.278194, 5.318223, 5.345743, 
    5.35758, 5.352668, 5.331766, 5.29685, 5.250499, 5.195425, 5.134211, 
    5.069193, 5.00797, 4.979156, 4.926097, 4.884192, 4.854754, 4.837235, 
    4.835485, 4.838983, 4.845691, 4.852136, 4.855419, 4.85442, 4.850298, 
    4.845923, 4.844999, 4.849974, 4.869821, 4.900551, 4.94209, 4.99318, 
    5.051761, 5.115341, 5.181213, 5.246534, 5.308325, 5.363435, 5.408561, 
    5.440397, 5.455967, 5.453187, 5.43158, 5.392928, 5.341514, 5.283599, 
    5.22609,
  // totalHeight(8,40, 0-49)
    5.079001, 5.113148, 5.155824, 5.20466, 5.255383, 5.302495, 5.340465, 
    5.364939, 5.373489, 5.365705, 5.342792, 5.306976, 5.260952, 5.2075, 
    5.149253, 5.093055, 5.064897, 5.0148, 4.972912, 4.940837, 4.918354, 
    4.909531, 4.905233, 4.904131, 4.903456, 4.901661, 4.898442, 4.895254, 
    4.894445, 4.899253, 4.911187, 4.93741, 4.973363, 5.018431, 5.071098, 
    5.129232, 5.190343, 5.251703, 5.310411, 5.363389, 5.407419, 5.439262, 
    5.455943, 5.455236, 5.436306, 5.400346, 5.350918, 5.293653, 5.235221, 
    5.181822,
  // totalHeight(8,41, 0-49)
    5.062121, 5.090923, 5.128824, 5.174737, 5.225716, 5.277128, 5.323496, 
    5.359679, 5.381943, 5.388488, 5.379393, 5.356171, 5.321213, 5.27729, 
    5.227234, 5.177218, 5.149961, 5.103456, 5.062327, 5.028457, 5.001982, 
    4.98717, 4.976339, 4.968845, 4.962564, 4.957095, 4.952728, 4.950969, 
    4.953513, 4.963099, 4.980418, 5.011087, 5.050213, 5.096777, 5.149055, 
    5.204819, 5.261506, 5.316321, 5.366274, 5.40823, 5.439034, 5.455762, 
    5.456133, 5.439089, 5.405383, 5.35795, 5.301758, 5.242993, 5.187772, 
    5.140857,
  // totalHeight(8,42, 0-49)
    5.046977, 5.07022, 5.102299, 5.143245, 5.191529, 5.243844, 5.29543, 
    5.341003, 5.375879, 5.396879, 5.402698, 5.393766, 5.371802, 5.339299, 
    5.299088, 5.256725, 5.231469, 5.189376, 5.149957, 5.115338, 5.086065, 
    5.066585, 5.050688, 5.038368, 5.028037, 5.02018, 5.015453, 5.015247, 
    5.020588, 5.033757, 5.054786, 5.087964, 5.128242, 5.174273, 5.224139, 
    5.275482, 5.32564, 5.371724, 5.410694, 5.439491, 5.455265, 5.455751, 
    5.439777, 5.407797, 5.36226, 5.307529, 5.249246, 5.193198, 5.144154, 
    5.105088,
  // totalHeight(8,43, 0-49)
    5.034163, 5.052107, 5.077977, 5.1126, 5.155713, 5.205489, 5.25843, 
    5.309834, 5.354713, 5.388844, 5.409515, 5.415804, 5.408386, 5.389111, 
    5.360541, 5.327561, 5.306041, 5.269506, 5.233062, 5.199059, 5.168477, 
    5.145934, 5.126657, 5.111196, 5.098354, 5.089241, 5.084676, 5.085835, 
    5.093141, 5.108504, 5.131452, 5.165137, 5.204473, 5.247838, 5.293118, 
    5.337825, 5.379192, 5.41429, 5.440164, 5.454059, 5.453766, 5.438076, 
    5.407258, 5.363396, 5.310354, 5.253236, 5.197416, 5.147466, 5.106408, 
    5.075515,
  // totalHeight(8,44, 0-49)
    5.023893, 5.037152, 5.057038, 5.08481, 5.121122, 5.165492, 5.215907, 
    5.268845, 5.319784, 5.364102, 5.398016, 5.419214, 5.427063, 5.422406, 
    5.407182, 5.385447, 5.369846, 5.3404, 5.308588, 5.276946, 5.246899, 
    5.223215, 5.202463, 5.185639, 5.171791, 5.162381, 5.15825, 5.160318, 
    5.168521, 5.184505, 5.207436, 5.239498, 5.275653, 5.314039, 5.352384, 
    5.388091, 5.418369, 5.440388, 5.451512, 5.449613, 5.433495, 5.403317, 
    5.360887, 5.309646, 5.254205, 5.199492, 5.149795, 5.108033, 5.075538, 
    5.052284,
  // totalHeight(8,45, 0-49)
    5.016068, 5.025445, 5.040023, 5.06117, 5.090047, 5.127151, 5.171838, 
    5.22204, 5.274341, 5.324514, 5.368355, 5.402508, 5.425014, 5.435463, 
    5.434813, 5.426049, 5.418765, 5.398278, 5.373139, 5.345995, 5.318683, 
    5.296079, 5.275944, 5.259601, 5.246169, 5.237257, 5.233617, 5.23592, 
    5.243749, 5.258614, 5.279437, 5.307597, 5.338169, 5.369109, 5.398049, 
    5.4224, 5.439507, 5.446893, 5.442554, 5.425341, 5.395344, 5.354149, 
    5.304817, 5.251482, 5.198609, 5.150136, 5.108815, 5.075948, 5.051572, 
    5.034879,
  // totalHeight(8,46, 0-49)
    5.010371, 5.016713, 5.026895, 5.042174, 5.063859, 5.092983, 5.129908, 
    5.173916, 5.222999, 5.273985, 5.323053, 5.366474, 5.401325, 5.425965, 
    5.440145, 5.44553, 5.448809, 5.439283, 5.423095, 5.402858, 5.380724, 
    5.361625, 5.344312, 5.33029, 5.318596, 5.310812, 5.307542, 5.309251, 
    5.315293, 5.327178, 5.343702, 5.365603, 5.388121, 5.409129, 5.4263, 
    5.437255, 5.439753, 5.431987, 5.41292, 5.382617, 5.342471, 5.295172, 
    5.244368, 5.194016, 5.147643, 5.107752, 5.075573, 5.051174, 5.03382, 
    5.022387,
  // totalHeight(8,47, 0-49)
    5.006379, 5.010458, 5.017199, 5.027631, 5.042955, 5.064367, 5.092776, 
    5.128459, 5.170724, 5.217763, 5.2668, 5.314528, 5.357748, 5.393965, 
    5.421778, 5.441412, 5.456867, 5.46001, 5.454927, 5.44398, 5.429455, 
    5.416289, 5.403948, 5.393989, 5.385193, 5.379011, 5.375869, 5.37608, 
    5.378881, 5.385936, 5.396016, 5.409431, 5.421616, 5.430514, 5.434071, 
    5.430398, 5.418005, 5.396079, 5.364757, 5.325294, 5.280035, 5.23211, 
    5.184909, 5.141459, 5.10393, 5.073397, 5.049934, 5.032877, 5.021182, 
    5.013739,
  // totalHeight(8,48, 0-49)
    5.003644, 5.006086, 5.010241, 5.016864, 5.02692, 5.041507, 5.061704, 
    5.088339, 5.121694, 5.161249, 5.20556, 5.252367, 5.298956, 5.342635, 
    5.381233, 5.413701, 5.441738, 5.458355, 5.465828, 5.466006, 5.46107, 
    5.455938, 5.450424, 5.446013, 5.441033, 5.436764, 5.433451, 5.431307, 
    5.42953, 5.430123, 5.431936, 5.435133, 5.435347, 5.430807, 5.42, 
    5.401847, 5.375895, 5.342507, 5.302944, 5.259302, 5.21424, 5.17055, 
    5.13068, 5.096348, 5.068379, 5.046762, 5.030877, 5.019772, 5.012416, 
    5.007883,
  // totalHeight(8,49, 0-49)
    5.001472, 5.002565, 5.00451, 5.007768, 5.012981, 5.020984, 5.032765, 
    5.049376, 5.071753, 5.100489, 5.135601, 5.176348, 5.22122, 5.268123, 
    5.314735, 5.359285, 5.403051, 5.435205, 5.457379, 5.470873, 5.477746, 
    5.48514, 5.4914, 5.497845, 5.49962, 5.498258, 5.49363, 5.486034, 
    5.474223, 5.463232, 5.452115, 5.442515, 5.428285, 5.40822, 5.38172, 
    5.348891, 5.31062, 5.268536, 5.22482, 5.181884, 5.141978, 5.106841, 
    5.077487, 5.054176, 5.036537, 5.023789, 5.01498, 5.009157, 5.005493, 
    5.003342,
  // totalHeight(9,0, 0-49)
    5.013042, 5.019694, 5.029954, 5.044734, 5.064919, 5.091146, 5.123545, 
    5.161498, 5.203522, 5.247341, 5.290179, 5.329203, 5.361989, 5.386886, 
    5.403194, 5.411325, 5.413615, 5.407965, 5.397056, 5.382667, 5.366389, 
    5.350346, 5.335258, 5.322433, 5.312547, 5.306667, 5.305348, 5.308775, 
    5.316498, 5.328191, 5.342663, 5.358954, 5.37482, 5.38847, 5.398046, 
    5.401766, 5.398109, 5.386037, 5.365193, 5.336077, 5.300086, 5.259408, 
    5.216734, 5.174833, 5.136135, 5.102393, 5.074556, 5.052821, 5.03683, 
    5.025922,
  // totalHeight(9,1, 0-49)
    5.018539, 5.027684, 5.041417, 5.060682, 5.086233, 5.118349, 5.15655, 
    5.19942, 5.244636, 5.289235, 5.330095, 5.364451, 5.390327, 5.406764, 
    5.413841, 5.412899, 5.408258, 5.395083, 5.37753, 5.357601, 5.33689, 
    5.31798, 5.300873, 5.28678, 5.275898, 5.269395, 5.267859, 5.271605, 
    5.28021, 5.293866, 5.31147, 5.332596, 5.354544, 5.375515, 5.393538, 
    5.406585, 5.412741, 5.410409, 5.398545, 5.376884, 5.346107, 5.307889, 
    5.264752, 5.219728, 5.175877, 5.135812, 5.10137, 5.073483, 5.052285, 
    5.037354,
  // totalHeight(9,2, 0-49)
    5.026684, 5.039216, 5.057403, 5.082047, 5.113499, 5.151348, 5.194202, 
    5.239692, 5.284729, 5.326012, 5.360569, 5.386237, 5.401902, 5.407519, 
    5.403984, 5.393466, 5.38223, 5.362339, 5.339471, 5.315671, 5.292365, 
    5.272373, 5.254879, 5.240854, 5.229998, 5.223449, 5.221773, 5.225418, 
    5.234077, 5.248452, 5.26766, 5.291913, 5.318253, 5.345037, 5.370354, 
    5.392126, 5.40825, 5.416761, 5.416035, 5.405025, 5.383495, 5.35221, 
    5.312987, 5.268557, 5.222194, 5.177207, 5.136419, 5.101797, 5.074339, 
    5.054193,
  // totalHeight(9,3, 0-49)
    5.037796, 5.054545, 5.077931, 5.108358, 5.145469, 5.18788, 5.233158, 
    5.278073, 5.319133, 5.353187, 5.377922, 5.392138, 5.395739, 5.389587, 
    5.375238, 5.355539, 5.338708, 5.313167, 5.286374, 5.260293, 5.236083, 
    5.216662, 5.200305, 5.187636, 5.177845, 5.171894, 5.170265, 5.173514, 
    5.181518, 5.195473, 5.21482, 5.240509, 5.269487, 5.300368, 5.331426, 
    5.360679, 5.385998, 5.405237, 5.416381, 5.417744, 5.408212, 5.3875, 
    5.356378, 5.316756, 5.271558, 5.224334, 5.17869, 5.137706, 5.103526, 
    5.07722,
  // totalHeight(9,4, 0-49)
    5.052035, 5.073641, 5.102532, 5.138441, 5.180034, 5.224841, 5.269492, 
    5.310276, 5.3438, 5.367561, 5.380238, 5.381697, 5.372798, 5.355103, 
    5.330607, 5.30267, 5.281563, 5.251438, 5.221951, 5.194925, 5.171211, 
    5.153751, 5.139843, 5.129701, 5.121983, 5.117336, 5.116074, 5.11881, 
    5.125641, 5.138234, 5.156425, 5.182015, 5.211965, 5.245227, 5.280334, 
    5.31548, 5.34862, 5.37757, 5.400111, 5.414134, 5.417838, 5.409997, 
    5.390258, 5.359409, 5.319504, 5.273733, 5.225988, 5.18022, 5.139762, 
    5.106874,
  // totalHeight(9,5, 0-49)
    5.06927, 5.096024, 5.130133, 5.170412, 5.21444, 5.258764, 5.299453, 
    5.332823, 5.356091, 5.367723, 5.367478, 5.356185, 5.335419, 5.307194, 
    5.273708, 5.238726, 5.214715, 5.180921, 5.149723, 5.122785, 5.100636, 
    5.086227, 5.075836, 5.069233, 5.064543, 5.061961, 5.061525, 5.063834, 
    5.069201, 5.079716, 5.095667, 5.119814, 5.149218, 5.18323, 5.220694, 
    5.260019, 5.299302, 5.336403, 5.369049, 5.394906, 5.411742, 5.417627, 
    5.411244, 5.392218, 5.361438, 5.321201, 5.275047, 5.227249, 5.182064, 
    5.142961,
  // totalHeight(9,6, 0-49)
    5.088974, 5.120697, 5.159075, 5.201886, 5.245714, 5.28647, 5.320168, 
    5.343662, 5.355105, 5.354039, 5.341181, 5.318075, 5.28674, 5.249392, 
    5.208251, 5.167442, 5.141766, 5.105011, 5.072841, 5.046739, 5.026933, 
    5.016384, 5.01034, 5.008129, 5.007359, 5.007643, 5.008629, 5.010802, 
    5.014644, 5.022597, 5.035425, 5.056958, 5.084433, 5.117664, 5.155847, 
    5.197634, 5.241279, 5.284737, 5.325753, 5.361929, 5.390816, 5.410064, 
    5.417652, 5.412226, 5.393486, 5.362525, 5.321963, 5.275724, 5.22841, 
    5.184418,
  // totalHeight(9,7, 0-49)
    5.110209, 5.146196, 5.187303, 5.230341, 5.2712, 5.305634, 5.330105, 
    5.342353, 5.341588, 5.328314, 5.30397, 5.270539, 5.230231, 5.185272, 
    5.137776, 5.092242, 5.065883, 5.026673, 4.994061, 4.969322, 4.952398, 
    4.94629, 4.94522, 4.948102, 4.952066, 4.956038, 4.959166, 4.961686, 
    4.96418, 4.969313, 4.978322, 4.996211, 5.020468, 5.051454, 5.088767, 
    5.131334, 5.177573, 5.225541, 5.273042, 5.317697, 5.356995, 5.388387, 
    5.409444, 5.418111, 5.413079, 5.394205, 5.362855, 5.321998, 5.275874, 
    5.22923,
  // totalHeight(9,8, 0-49)
    5.131696, 5.170769, 5.212703, 5.253581, 5.289032, 5.315145, 5.329186, 
    5.329929, 5.317555, 5.293313, 5.25909, 5.217057, 5.16942, 5.118283, 
    5.06558, 5.016235, 4.989789, 4.94848, 4.915803, 4.892795, 4.879127, 
    4.877858, 4.882214, 4.890742, 4.900167, 4.908644, 4.914731, 4.918277, 
    4.919837, 4.922133, 4.926813, 4.940151, 4.959956, 4.987245, 5.022112, 
    5.063804, 5.110915, 5.161597, 5.213713, 5.264927, 5.312754, 5.354599, 
    5.387856, 5.410053, 5.419156, 5.413955, 5.394502, 5.362439, 5.321009, 
    5.274606,
  // totalHeight(9,9, 0-49)
    5.152001, 5.192673, 5.233472, 5.270114, 5.29842, 5.315174, 5.318628, 
    5.308538, 5.285864, 5.252336, 5.21005, 5.161165, 5.107756, 5.051719, 
    4.994766, 4.942291, 4.915819, 4.872682, 4.84023, 4.81922, 4.809059, 
    4.812881, 4.822952, 4.837524, 4.85301, 4.866771, 4.876707, 4.882144, 
    4.883457, 4.883184, 4.883249, 4.891264, 4.905428, 4.927546, 4.95835, 
    4.997493, 5.043778, 5.095445, 5.150386, 5.2063, 5.260748, 5.311169, 
    5.354927, 5.389367, 5.412012, 5.420855, 5.414785, 5.39402, 5.360405, 
    5.317352,
  // totalHeight(9,10, 0-49)
    5.169785, 5.210491, 5.248452, 5.279398, 5.299693, 5.307023, 5.300615, 
    5.281043, 5.249805, 5.208882, 5.160379, 5.106323, 5.048559, 4.988734, 
    4.928304, 4.873112, 4.845929, 4.801261, 4.769295, 4.750492, 4.743991, 
    4.753007, 4.768904, 4.789725, 4.811697, 4.831421, 4.846126, 4.854508, 
    4.856575, 4.854371, 4.849869, 4.852006, 4.859412, 4.874855, 4.899894, 
    4.934735, 4.978467, 5.029416, 5.085478, 5.144336, 5.203576, 5.260691, 
    5.313084, 5.358071, 5.392953, 5.41521, 5.422825, 5.414724, 5.391241, 
    5.354405,
  // totalHeight(9,11, 0-49)
    5.184051, 5.223395, 5.257313, 5.281863, 5.294163, 5.292828, 5.27793, 
    5.25065, 5.212797, 5.166412, 5.113485, 5.055821, 4.994998, 4.932372, 
    4.869107, 4.811265, 4.781673, 4.735917, 4.704734, 4.688303, 4.685516, 
    4.699636, 4.72124, 4.748251, 4.776879, 4.803067, 4.823434, 4.835981, 
    4.840165, 4.837159, 4.828632, 4.824708, 4.824437, 4.831717, 4.849192, 
    4.877854, 4.917208, 4.965708, 5.021219, 5.081358, 5.143673, 5.205681, 
    5.264839, 5.318503, 5.363908, 5.398248, 5.41888, 5.423704, 5.411665, 
    5.383304,
  // totalHeight(9,12, 0-49)
    5.194335, 5.231282, 5.260574, 5.278791, 5.28386, 5.275225, 5.253618, 
    5.220604, 5.178126, 5.128154, 5.072487, 5.012671, 4.949991, 4.885493, 
    4.82, 4.759103, 4.724104, 4.677974, 4.647959, 4.634027, 4.634865, 
    4.653734, 4.680614, 4.713413, 4.74852, 4.781399, 4.808202, 4.826231, 
    4.834251, 4.832163, 4.82086, 4.811296, 4.802845, 4.800652, 4.808741, 
    4.829211, 4.862217, 4.906439, 4.959705, 5.019504, 5.083271, 5.148478, 
    5.212607, 5.273064, 5.327098, 5.371778, 5.404087, 5.421196, 5.420952, 
    5.402519,
  // totalHeight(9,13, 0-49)
    5.20077, 5.234771, 5.259482, 5.27208, 5.271227, 5.25703, 5.230669, 
    5.19392, 5.148717, 5.09689, 5.04002, 4.97939, 4.916002, 4.850582, 
    4.783556, 4.718486, 4.673654, 4.628222, 4.599886, 4.588519, 4.592689, 
    4.615596, 4.646937, 4.684716, 4.725712, 4.765153, 4.798926, 4.823727, 
    4.837541, 4.838665, 4.826695, 4.812769, 4.796377, 4.783873, 4.780921, 
    4.791139, 4.815689, 4.853671, 4.902922, 4.960753, 5.024401, 5.091208, 
    5.158616, 5.22405, 5.284799, 5.337901, 5.380161, 5.408309, 5.419418, 
    5.411558,
  // totalHeight(9,14, 0-49)
    5.204044, 5.235059, 5.255784, 5.26395, 5.258807, 5.240928, 5.211757, 
    5.173126, 5.126891, 5.074712, 5.01796, 4.9577, 4.894693, 4.829371, 
    4.761736, 4.690343, 4.630024, 4.586733, 4.560706, 4.551862, 4.558817, 
    4.584635, 4.619225, 4.660789, 4.706684, 4.75217, 4.793106, 4.82573, 
    4.84728, 4.85427, 4.84457, 4.828547, 4.805531, 4.782758, 4.767636, 
    4.765727, 4.779678, 4.809348, 4.852722, 4.90692, 4.968901, 5.035783, 
    5.104878, 5.173582, 5.2392, 5.2988, 5.349137, 5.386735, 5.408215, 5.410872,
  // totalHeight(9,15, 0-49)
    5.205245, 5.233704, 5.251448, 5.256646, 5.248955, 5.229216, 5.198977, 
    5.160035, 5.114126, 5.062756, 5.007135, 4.948183, 4.886503, 4.822322, 
    4.75529, 4.674098, 4.592133, 4.552732, 4.529696, 4.523179, 4.532108, 
    4.559325, 4.595654, 4.639558, 4.689092, 4.739789, 4.787691, 4.828758, 
    4.859601, 4.875039, 4.871017, 4.856003, 4.828897, 4.797172, 4.769747, 
    4.754407, 4.755836, 4.775146, 4.810735, 4.859603, 4.918382, 4.983872, 
    5.053164, 5.123552, 5.192328, 5.2566, 5.31316, 5.358506, 5.389058, 5.40165,
  // totalHeight(9,16, 0-49)
    5.205641, 5.232349, 5.248367, 5.25215, 5.243571, 5.223566, 5.193663, 
    5.155571, 5.1109, 5.061044, 5.007129, 4.950017, 4.890282, 4.828084, 
    4.762897, 4.667199, 4.558082, 4.524595, 4.505179, 4.500589, 4.510473, 
    4.537367, 4.573853, 4.618652, 4.670533, 4.725457, 4.779788, 4.82938, 
    4.870381, 4.896234, 4.90115, 4.890569, 4.862889, 4.82492, 4.786451, 
    4.75743, 4.745025, 4.7522, 4.7782, 4.820086, 4.874176, 4.936878, 
    5.004986, 5.075613, 5.145999, 5.21328, 5.274343, 5.325768, 5.363969, 
    5.385563,
  // totalHeight(9,17, 0-49)
    5.206429, 5.23244, 5.24809, 5.25195, 5.243927, 5.22491, 5.196322, 
    5.159752, 5.116711, 5.068528, 5.016322, 4.960996, 4.903182, 4.84309, 
    4.780164, 4.665139, 4.525096, 4.499957, 4.484663, 4.481379, 4.491128, 
    4.516054, 4.551351, 4.595904, 4.649085, 4.707342, 4.767391, 4.825082, 
    4.876275, 4.913509, 4.929801, 4.926649, 4.902213, 4.861757, 4.814963, 
    4.77341, 4.746902, 4.740796, 4.755741, 4.789182, 4.837222, 4.895868, 
    4.96155, 5.03114, 5.101774, 5.170614, 5.234653, 5.290627, 5.335063, 
    5.36453,
  // totalHeight(9,18, 0-49)
    5.208497, 5.234978, 5.251599, 5.256881, 5.250602, 5.233477, 5.206757, 
    5.171896, 5.13033, 5.083377, 5.032204, 4.977786, 4.920807, 4.861402, 
    4.798707, 4.662005, 4.489505, 4.475817, 4.465091, 4.462282, 4.47091, 
    4.492671, 4.525987, 4.569733, 4.623669, 4.684685, 4.74978, 4.814837, 
    4.875535, 4.924022, 4.952873, 4.959058, 4.941103, 4.902152, 4.850769, 
    4.799243, 4.759669, 4.740109, 4.743153, 4.767068, 4.80796, 4.861491, 
    4.9237, 4.991181, 5.060933, 5.130117, 5.195842, 5.255026, 5.304377, 
    5.340523,
  // totalHeight(9,19, 0-49)
    5.212205, 5.240322, 5.25919, 5.267125, 5.263608, 5.249043, 5.224416, 
    5.191014, 5.150217, 5.103388, 5.051769, 4.996344, 4.937584, 4.874966, 
    4.806328, 4.651233, 4.447761, 4.448816, 4.443101, 4.439723, 4.446472, 
    4.464695, 4.496089, 4.539269, 4.594101, 4.657805, 4.727543, 4.799196, 
    4.868299, 4.927033, 4.968306, 4.984324, 4.974784, 4.940611, 4.888542, 
    4.830527, 4.780185, 4.748146, 4.739299, 4.753189, 4.786242, 4.833904, 
    4.891861, 4.956418, 5.024415, 5.092998, 5.159379, 5.220663, 5.273758, 
    5.315415,
  // totalHeight(9,20, 0-49)
    5.212728, 5.239095, 5.257136, 5.265122, 5.262591, 5.250175, 5.229265, 
    5.201706, 5.169541, 5.134852, 5.099675, 5.065902, 5.035129, 5.008301, 
    4.984965, 30, 4.281867, 4.296238, 4.319592, 4.349007, 4.384036, 4.42006, 
    4.463272, 4.513869, 4.573604, 4.641306, 4.715052, 4.791258, 4.865699, 
    4.931174, 4.981727, 5.005177, 5.003088, 4.974547, 4.924257, 4.862964, 
    4.804741, 4.762134, 4.742292, 4.746347, 4.771365, 4.812787, 4.866036, 
    4.927151, 4.99281, 5.06013, 5.12641, 5.188928, 5.244792, 5.290888,
  // totalHeight(9,21, 0-49)
    5.21802, 5.246518, 5.267158, 5.277958, 5.278198, 5.26831, 5.249588, 
    5.223853, 5.193182, 5.159711, 5.125531, 5.092601, 5.062645, 5.036921, 
    5.015751, 30, 4.280171, 4.286097, 4.301404, 4.32449, 4.355588, 4.38597, 
    4.42638, 4.475754, 4.535542, 4.604822, 4.681754, 4.762756, 4.84341, 
    4.91684, 4.978211, 5.011083, 5.019394, 5.000573, 4.957034, 4.897546, 
    4.835649, 4.785192, 4.75563, 4.750137, 4.766894, 4.801638, 4.849658, 
    4.906757, 4.969437, 5.034751, 5.100053, 5.162745, 5.22009, 5.269087,
  // totalHeight(9,22, 0-49)
    5.22302, 5.253256, 5.275841, 5.288589, 5.290601, 5.282212, 5.264708, 
    5.239964, 5.210128, 5.177406, 5.143931, 5.111705, 5.082527, 5.057864, 
    5.038573, 30, 4.278119, 4.278525, 4.288034, 4.306596, 4.335303, 4.361061, 
    4.399333, 4.447818, 4.507654, 4.578084, 4.657235, 4.741405, 4.825919, 
    4.904216, 4.972783, 5.011243, 5.026633, 5.015471, 4.978484, 4.922526, 
    4.859972, 4.804983, 4.768548, 4.755605, 4.765541, 4.794574, 4.838022, 
    4.891535, 4.95148, 5.014856, 5.079045, 5.141546, 5.199745, 5.250741,
  // totalHeight(9,23, 0-49)
    5.226744, 5.258028, 5.281734, 5.295559, 5.298512, 5.290893, 5.27401, 
    5.249787, 5.220436, 5.188205, 5.155255, 5.1236, 5.095076, 5.07127, 
    5.053352, 30, 4.279414, 4.276551, 4.281965, 4.297147, 4.32407, 4.345681, 
    4.381749, 4.428933, 4.488155, 4.558842, 4.639098, 4.725091, 4.811872, 
    4.893102, 4.966422, 5.00808, 5.028121, 5.022609, 4.991148, 4.939076, 
    4.877542, 4.820482, 4.779746, 4.76159, 4.766459, 4.791107, 4.830965, 
    4.881619, 4.93934, 5.001071, 5.064211, 5.126318, 5.184858, 5.237008,
  // totalHeight(9,24, 0-49)
    5.228496, 5.259939, 5.283836, 5.297881, 5.301076, 5.293717, 5.277114, 
    5.253204, 5.224204, 5.192366, 5.159845, 5.128648, 5.100616, 5.077384, 
    5.060251, 30, 4.283651, 4.279233, 4.282315, 4.295458, 4.321284, 4.339952, 
    4.374256, 4.42016, 4.47849, 4.548845, 4.629343, 4.716074, 4.803885, 
    4.886553, 4.962506, 5.005624, 5.028133, 5.025902, 4.997901, 4.948527, 
    4.888073, 4.830173, 4.787071, 4.765799, 4.767502, 4.789327, 4.826833, 
    4.875592, 4.931826, 4.992456, 5.054884, 5.116711, 5.175456, 5.228333,
  // totalHeight(9,25, 0-49)
    5.22796, 5.258594, 5.281716, 5.295139, 5.297939, 5.290426, 5.27388, 
    5.250185, 5.221498, 5.190021, 5.157872, 5.127028, 5.099308, 5.07633, 
    5.059365, 30, 4.289196, 4.284725, 4.287505, 4.300285, 4.325872, 4.343461, 
    4.376945, 4.422066, 4.479642, 4.549365, 4.629392, 4.715792, 4.803343, 
    4.885863, 4.962089, 5.004999, 5.027723, 5.026116, 4.998996, 4.950472, 
    4.89053, 4.832613, 4.789001, 4.766916, 4.767715, 4.788686, 4.825451, 
    4.87359, 4.929327, 4.989579, 5.051758, 5.113479, 5.17228, 5.22539,
  // totalHeight(9,26, 0-49)
    5.225247, 5.254143, 5.275551, 5.287515, 5.289261, 5.281141, 5.26438, 
    5.240758, 5.21231, 5.18114, 5.149289, 5.11869, 5.091106, 5.068068, 
    5.050664, 30, 4.295433, 4.292458, 4.29705, 4.311205, 4.33739, 4.355901, 
    4.389616, 4.434559, 4.491645, 4.560555, 4.639478, 4.724538, 4.810594, 
    4.891437, 4.965577, 5.006762, 5.027511, 5.023829, 4.99484, 4.945057, 
    4.88476, 4.827417, 4.78503, 4.764428, 4.766649, 4.788824, 4.826549, 
    4.875436, 4.931742, 4.99241, 5.054859, 5.116698, 5.175449, 5.22833,
  // totalHeight(9,27, 0-49)
    5.220861, 5.247246, 5.266091, 5.275759, 5.275703, 5.266364, 5.248924, 
    5.225036, 5.196589, 5.16555, 5.133861, 5.103376, 5.075775, 5.052415, 
    5.034029, 30, 4.302463, 4.302832, 4.311277, 4.328385, 4.355904, 4.377017, 
    4.411754, 4.456905, 4.513578, 4.58136, 4.658477, 4.741166, 4.824496, 
    4.902151, 4.97192, 5.009845, 5.026492, 5.018219, 4.984942, 4.932204, 
    4.871093, 4.815196, 4.775881, 4.759018, 4.764867, 4.790172, 4.830435, 
    4.881328, 4.939181, 5.000987, 5.064165, 5.126294, 5.184847, 5.237001,
  // totalHeight(9,28, 0-49)
    5.215629, 5.238973, 5.254549, 5.261092, 5.258357, 5.246945, 5.228058, 
    5.203263, 5.174317, 5.143045, 5.111273, 5.080747, 5.053013, 5.029168, 
    5.009374, 30, 4.311146, 4.317119, 4.331298, 4.35264, 4.382026, 4.406691, 
    4.442622, 4.4878, 4.543655, 4.609676, 4.684156, 4.763472, 4.842965, 
    4.916097, 4.979532, 5.0127, 5.023324, 5.008373, 4.969041, 4.912435, 
    4.850762, 4.797608, 4.763256, 4.75213, 4.763408, 4.793327, 4.837316, 
    4.891145, 4.951268, 5.014741, 5.078983, 5.141513, 5.199726, 5.250731,
  // totalHeight(9,29, 0-49)
    5.210575, 5.230656, 5.242446, 5.245065, 5.238635, 5.224026, 5.202578, 
    5.175876, 5.145615, 5.11352, 5.081297, 5.050559, 5.022669, 4.99836, 
    4.977002, 30, 4.32097, 4.335202, 4.357126, 4.384002, 4.415863, 4.444396, 
    4.481161, 4.525657, 4.579839, 4.643129, 4.713893, 4.78861, 4.862862, 
    4.929764, 4.984661, 5.011045, 5.013606, 4.990396, 4.944409, 4.88464, 
    4.824273, 4.776336, 4.749413, 4.746114, 4.764445, 4.80021, 4.84885, 
    4.906308, 4.96919, 5.034617, 5.099981, 5.162707, 5.22007, 5.269075,
  // totalHeight(9,30, 0-49)
    5.211185, 5.232265, 5.243868, 5.245254, 5.236584, 5.218601, 5.192334, 
    5.158899, 5.119413, 5.074954, 5.0265, 4.974833, 4.92029, 4.862335, 
    4.799018, 4.650102, 4.46623, 4.474145, 4.474097, 4.474111, 4.482029, 
    4.496277, 4.523712, 4.562758, 4.613616, 4.67399, 4.741224, 4.811243, 
    4.879523, 4.938704, 4.982891, 5.000132, 4.992626, 4.960247, 4.908324, 
    4.847715, 4.791922, 4.752495, 4.735684, 4.742134, 4.768816, 4.811302, 
    4.865192, 4.926679, 4.992549, 5.059987, 5.126332, 5.188886, 5.244769, 
    5.290876,
  // totalHeight(9,31, 0-49)
    5.20908, 5.227884, 5.236427, 5.234247, 5.221874, 5.200438, 5.171289, 
    5.135762, 5.095062, 5.050255, 5.002267, 4.951888, 4.899677, 4.845722, 
    4.789222, 4.658228, 4.501397, 4.496706, 4.493328, 4.495354, 4.506206, 
    4.525119, 4.554814, 4.594297, 4.643971, 4.701432, 4.764091, 4.828028, 
    4.888942, 4.939219, 4.972041, 4.980291, 4.964257, 4.925714, 4.87197, 
    4.814879, 4.767239, 4.738547, 4.732779, 4.749048, 4.783735, 4.832435, 
    4.89102, 4.955945, 5.024151, 5.092851, 5.159298, 5.220619, 5.273735, 
    5.315403,
  // totalHeight(9,32, 0-49)
    5.209422, 5.227388, 5.234317, 5.229859, 5.214752, 5.190379, 5.15834, 
    5.120173, 5.077215, 5.030576, 4.981167, 4.929723, 4.876769, 4.822464, 
    4.766259, 4.657221, 4.530038, 4.515179, 4.508562, 4.511379, 4.524328, 
    4.547682, 4.579953, 4.620469, 4.669526, 4.724418, 4.782448, 4.839732, 
    4.892161, 4.932154, 4.95264, 4.951416, 4.927637, 4.885253, 4.833202, 
    4.783412, 4.747004, 4.730926, 4.736993, 4.76317, 4.805598, 4.860101, 
    4.922898, 4.990724, 5.060675, 5.129973, 5.195764, 5.254982, 5.304353, 
    5.340511,
  // totalHeight(9,33, 0-49)
    5.211784, 5.230331, 5.23714, 5.231805, 5.215128, 5.188638, 5.154125, 
    5.113319, 5.067709, 5.018507, 4.966658, 4.912882, 4.857656, 4.801088, 
    4.742635, 4.653386, 4.555256, 4.532505, 4.522496, 4.524918, 4.538918, 
    4.565711, 4.600144, 4.641606, 4.68998, 4.742125, 4.795075, 4.84495, 
    4.887879, 4.916761, 4.925084, 4.915268, 4.8861, 4.843475, 4.797151, 
    4.758084, 4.735029, 4.73236, 4.75014, 4.785647, 4.835072, 4.894595, 
    4.960809, 5.030715, 5.101532, 5.170478, 5.234578, 5.290584, 5.33504, 
    5.364517,
  // totalHeight(9,34, 0-49)
    5.215219, 5.235668, 5.243885, 5.23924, 5.222435, 5.195026, 5.158927, 
    5.11603, 5.067999, 5.016191, 4.961662, 4.905194, 4.847309, 4.788183, 
    4.727444, 4.6529, 4.580625, 4.55162, 4.538008, 4.538926, 4.552721, 
    4.581357, 4.616908, 4.658594, 4.70565, 4.754443, 4.80167, 4.843497, 
    4.87642, 4.894343, 4.89206, 4.875939, 4.844918, 4.806159, 4.769204, 
    4.743195, 4.734305, 4.744707, 4.773262, 4.816971, 4.872271, 4.935742, 
    5.004318, 5.075227, 5.145776, 5.213154, 5.274272, 5.325727, 5.363947, 
    5.38555,
  // totalHeight(9,35, 0-49)
    5.218414, 5.241881, 5.252987, 5.250708, 5.235466, 5.208694, 5.172336, 
    5.12841, 5.078754, 5.02491, 4.968103, 4.90927, 4.849085, 4.787934, 
    4.725807, 4.660797, 4.609091, 4.575197, 4.557967, 4.556472, 4.56875, 
    4.597325, 4.632507, 4.673204, 4.717884, 4.762468, 4.803359, 4.83689, 
    4.860095, 4.868361, 4.85827, 4.839107, 4.810142, 4.778883, 4.753745, 
    4.741656, 4.746446, 4.768659, 4.806472, 4.856906, 4.916722, 4.98287, 
    5.052571, 5.123204, 5.192127, 5.256485, 5.313095, 5.358469, 5.389037, 
    5.401639,
  // totalHeight(9,36, 0-49)
    5.219895, 5.247176, 5.262488, 5.264244, 5.252396, 5.228087, 5.193159, 
    5.149686, 5.099665, 5.044836, 4.98664, 4.926233, 4.864524, 4.80219, 
    4.739642, 4.680242, 4.642906, 4.605454, 4.584847, 4.580313, 4.589905, 
    4.616549, 4.649711, 4.687962, 4.729007, 4.768494, 4.802673, 4.828212, 
    4.842849, 4.843726, 4.829322, 4.810611, 4.787079, 4.765726, 4.753314, 
    4.754615, 4.771617, 4.803811, 4.849074, 4.904593, 4.967452, 5.034897, 
    5.104344, 5.173264, 5.239013, 5.29869, 5.349073, 5.3867, 5.408195, 
    5.410862,
  // totalHeight(9,37, 0-49)
    5.218255, 5.249717, 5.27024, 5.277552, 5.270936, 5.25105, 5.219474, 
    5.178236, 5.129437, 5.075015, 5.016646, 4.955743, 4.893483, 4.830852, 
    4.76865, 4.712382, 4.683611, 4.643882, 4.620321, 4.612436, 4.618487, 
    4.641649, 4.671282, 4.705679, 4.741915, 4.775605, 4.803057, 4.82145, 
    4.829312, 4.825551, 4.810279, 4.794975, 4.779095, 4.768571, 4.768416, 
    4.7816, 4.808813, 4.848932, 4.899767, 4.958707, 5.023099, 5.090394, 
    5.158112, 5.223743, 5.284613, 5.33779, 5.380095, 5.408271, 5.419396, 
    5.411546,
  // totalHeight(9,38, 0-49)
    5.212383, 5.247881, 5.274166, 5.288225, 5.288517, 5.274992, 5.248788, 
    5.21174, 5.165967, 5.113562, 5.056436, 4.996264, 4.934503, 4.87243, 
    4.811168, 4.756728, 4.73197, 4.691082, 4.665075, 4.653807, 4.65584, 
    4.674464, 4.699435, 4.72888, 4.759443, 4.786973, 4.808064, 4.820529, 
    4.823663, 4.81791, 4.804527, 4.794577, 4.787253, 4.787226, 4.797941, 
    4.821002, 4.856258, 4.902263, 4.956853, 5.017594, 5.082009, 5.147655, 
    5.212077, 5.272727, 5.326886, 5.371646, 5.404006, 5.421148, 5.420925, 
    5.402503,
  // totalHeight(9,39, 0-49)
    5.20167, 5.240501, 5.272511, 5.294001, 5.302503, 5.297089, 5.278226, 
    5.247378, 5.20655, 5.157911, 5.103568, 5.045445, 4.985273, 4.924599, 
    4.864816, 4.811718, 4.787943, 4.746778, 4.718848, 4.70439, 4.702281, 
    4.715828, 4.73548, 4.759322, 4.783782, 4.805178, 4.82057, 4.828451, 
    4.828772, 4.823126, 4.813404, 4.809672, 4.810735, 4.820044, 4.839785, 
    4.870599, 4.911798, 4.96177, 5.018401, 5.079369, 5.142285, 5.204723, 
    5.264188, 5.318067, 5.363621, 5.398062, 5.418763, 5.423631, 5.411623, 
    5.383276,
  // totalHeight(9,40, 0-49)
    5.186132, 5.22708, 5.264103, 5.293013, 5.310456, 5.314495, 5.304725, 
    5.282016, 5.248078, 5.205032, 5.155106, 5.100437, 5.043005, 4.984615, 
    4.926899, 4.87519, 4.850765, 4.809989, 4.780656, 4.763356, 4.757268, 
    4.765635, 4.779768, 4.797813, 4.816178, 4.8318, 4.84232, 4.846885, 
    4.845916, 4.841768, 4.836526, 4.838995, 4.847562, 4.864634, 4.891436, 
    4.927948, 4.973135, 5.025293, 5.082327, 5.141959, 5.201804, 5.259393, 
    5.312152, 5.357416, 5.392503, 5.414909, 5.422629, 5.414599, 5.391162, 
    5.354355,
  // totalHeight(9,41, 0-49)
    5.166451, 5.207902, 5.248558, 5.28407, 5.310394, 5.324593, 5.325236, 
    5.312375, 5.287194, 5.251593, 5.207793, 5.158082, 5.10465, 5.049539, 
    4.994611, 4.944724, 4.91911, 4.879265, 4.849064, 4.829385, 4.819679, 
    4.823095, 4.831874, 4.844314, 4.856938, 4.867391, 4.873917, 4.876226, 
    4.875024, 4.873092, 4.872416, 4.880478, 4.895287, 4.918398, 4.950332, 
    4.990605, 5.037953, 5.090587, 5.146398, 5.203084, 5.258206, 5.309211, 
    5.353455, 5.388292, 5.41125, 5.42033, 5.414435, 5.393792, 5.360259, 
    5.317256,
  // totalHeight(9,42, 0-49)
    5.143857, 5.184021, 5.226386, 5.266863, 5.301079, 5.325276, 5.336976, 
    5.335222, 5.320437, 5.294066, 5.258155, 5.215016, 5.166993, 5.116336, 
    5.06512, 5.017797, 4.99126, 4.952888, 4.922406, 4.90091, 4.888094, 
    4.887012, 4.890862, 4.898168, 4.905657, 4.911681, 4.915056, 4.915931, 
    4.915131, 4.915613, 4.919096, 4.931798, 4.951411, 4.978819, 5.014019, 
    5.056201, 5.103926, 5.155319, 5.208214, 5.260242, 5.308877, 5.35149, 
    5.38544, 5.408236, 5.417833, 5.413025, 5.393868, 5.362019, 5.320735, 
    5.274421,
  // totalHeight(9,43, 0-49)
    5.119925, 5.157089, 5.198948, 5.24208, 5.282256, 5.315266, 5.337736, 
    5.347641, 5.344442, 5.32887, 5.302574, 5.267717, 5.226689, 5.18188, 
    5.135561, 5.09184, 5.065246, 5.028996, 4.998917, 4.976262, 4.960958, 
    4.95599, 4.955519, 4.958347, 4.961455, 4.963848, 4.964833, 4.96487, 
    4.964771, 4.967505, 4.974444, 4.990649, 5.013561, 5.043531, 5.080167, 
    5.122412, 5.168684, 5.217022, 5.265179, 5.3107, 5.350989, 5.383418, 
    5.405475, 5.415052, 5.410805, 5.392574, 5.361722, 5.321233, 5.275365, 
    5.228883,
  // totalHeight(9,44, 0-49)
    5.096272, 5.129057, 5.168241, 5.211352, 5.254784, 5.29438, 5.326228, 
    5.34737, 5.35621, 5.352563, 5.337418, 5.312571, 5.280278, 5.24296, 
    5.203005, 5.164229, 5.138921, 5.105624, 5.076772, 5.053725, 5.036647, 
    5.028522, 5.024458, 5.023581, 5.023133, 5.022689, 5.021945, 5.021548, 
    5.022201, 5.026792, 5.036315, 5.054803, 5.079486, 5.110286, 5.146511, 
    5.186906, 5.22978, 5.273088, 5.314514, 5.351556, 5.381634, 5.402251, 
    5.411257, 5.407187, 5.389662, 5.359727, 5.319985, 5.274365, 5.22749, 
    5.183779,
  // totalHeight(9,45, 0-49)
    5.074281, 5.101814, 5.136524, 5.17699, 5.220571, 5.263685, 5.302406, 
    5.333194, 5.353523, 5.36219, 5.359307, 5.346044, 5.324288, 5.296298, 
    5.264447, 5.232249, 5.209951, 5.180675, 5.154027, 5.131465, 5.113417, 
    5.102954, 5.096113, 5.092372, 5.089212, 5.08668, 5.084756, 5.084169, 
    5.085434, 5.091334, 5.102482, 5.122004, 5.14693, 5.17682, 5.210737, 
    5.247275, 5.284656, 5.320791, 5.353364, 5.379928, 5.39808, 5.405691, 
    5.401236, 5.384155, 5.355194, 5.316544, 5.271692, 5.224903, 5.180446, 
    5.141823,
  // totalHeight(9,46, 0-49)
    5.0549, 5.07686, 5.105901, 5.141548, 5.18226, 5.22542, 5.26764, 5.305339, 
    5.335418, 5.355771, 5.36553, 5.365007, 5.355437, 5.338662, 5.316822, 
    5.293051, 5.275785, 5.251806, 5.228491, 5.207395, 5.189259, 5.177374, 
    5.168643, 5.162926, 5.157879, 5.153938, 5.151259, 5.150574, 5.152169, 
    5.158724, 5.17048, 5.189789, 5.213448, 5.240694, 5.270373, 5.30097, 
    5.330666, 5.357411, 5.379015, 5.393284, 5.398237, 5.392398, 5.375129, 
    5.346938, 5.309633, 5.26622, 5.22047, 5.176284, 5.136996, 5.104896,
  // totalHeight(9,47, 0-49)
    5.038558, 5.055104, 5.07795, 5.107332, 5.142719, 5.182619, 5.224613, 
    5.265657, 5.302625, 5.332863, 5.354623, 5.367231, 5.371015, 5.367095, 
    5.3571, 5.343633, 5.333583, 5.316318, 5.297566, 5.279008, 5.261748, 
    5.249465, 5.23981, 5.233042, 5.226902, 5.222136, 5.219, 5.218166, 
    5.219665, 5.226124, 5.237422, 5.255292, 5.276211, 5.299119, 5.322676, 
    5.345291, 5.365184, 5.380476, 5.389296, 5.389965, 5.381234, 5.362558, 
    5.334355, 5.298147, 5.256485, 5.212605, 5.169889, 5.131297, 5.098928, 
    5.073874,
  // totalHeight(9,48, 0-49)
    5.025191, 5.036808, 5.053524, 5.076003, 5.104483, 5.138533, 5.17689, 
    5.217495, 5.257764, 5.295023, 5.326963, 5.351994, 5.369394, 5.379289, 
    5.382505, 5.380936, 5.380241, 5.371087, 5.358146, 5.343263, 5.327931, 
    5.316406, 5.306894, 5.300048, 5.293569, 5.288468, 5.285032, 5.28385, 
    5.284679, 5.29018, 5.29989, 5.31511, 5.331882, 5.348882, 5.364614, 
    5.377472, 5.385822, 5.388123, 5.38307, 5.369785, 5.348024, 5.318344, 
    5.282197, 5.241826, 5.199984, 5.1595, 5.122818, 5.091662, 5.06691, 
    5.048687,
  // totalHeight(9,49, 0-49)
    5.012385, 5.018913, 5.028864, 5.043107, 5.062448, 5.087427, 5.118075, 
    5.153737, 5.193004, 5.233839, 5.273879, 5.31083, 5.342823, 5.368688, 
    5.388059, 5.402215, 5.418763, 5.421006, 5.415788, 5.405649, 5.392869, 
    5.385442, 5.379874, 5.377387, 5.372908, 5.368307, 5.363704, 5.359727, 
    5.355256, 5.355647, 5.359989, 5.371101, 5.38187, 5.390671, 5.395897, 
    5.396035, 5.389802, 5.3763, 5.355184, 5.326793, 5.292233, 5.253324, 
    5.212403, 5.171985, 5.134371, 5.101318, 5.073847, 5.052252, 5.036246, 
    5.025198,
  // totalHeight(10,0, 0-49)
    5.063582, 5.085031, 5.112928, 5.146696, 5.184947, 5.225497, 5.265574, 
    5.302221, 5.332746, 5.355133, 5.368267, 5.371976, 5.366912, 5.354355, 
    5.335983, 5.3139, 5.291661, 5.267425, 5.244224, 5.223267, 5.205225, 
    5.190944, 5.179907, 5.172104, 5.167113, 5.164995, 5.165788, 5.169702, 
    5.176876, 5.187829, 5.202584, 5.221438, 5.243492, 5.268015, 5.293913, 
    5.31977, 5.34392, 5.364543, 5.379786, 5.387915, 5.38752, 5.377726, 
    5.358419, 5.3304, 5.295416, 5.256012, 5.215207, 5.176044, 5.141145, 
    5.112394,
  // totalHeight(10,1, 0-49)
    5.079928, 5.105417, 5.137311, 5.174423, 5.214681, 5.255301, 5.293159, 
    5.325284, 5.349298, 5.363727, 5.368092, 5.362825, 5.349079, 5.32849, 
    5.302971, 5.274961, 5.249591, 5.22163, 5.19565, 5.1729, 5.153946, 
    5.139993, 5.129792, 5.123188, 5.119247, 5.117973, 5.119292, 5.123413, 
    5.130458, 5.141384, 5.156361, 5.176321, 5.200119, 5.227235, 5.256737, 
    5.287312, 5.31734, 5.344975, 5.368256, 5.385231, 5.394138, 5.393606, 
    5.382902, 5.362143, 5.332445, 5.295923, 5.255486, 5.214435, 5.175961, 
    5.142664,
  // totalHeight(10,2, 0-49)
    5.100276, 5.12977, 5.1649, 5.203756, 5.243615, 5.281312, 5.313743, 
    5.338332, 5.35337, 5.358143, 5.352868, 5.338513, 5.316582, 5.288897, 
    5.257421, 5.224789, 5.197577, 5.167107, 5.139554, 5.116156, 5.097363, 
    5.084681, 5.076171, 5.071518, 5.069331, 5.069472, 5.071693, 5.076145, 
    5.082903, 5.093283, 5.107612, 5.127469, 5.151559, 5.179631, 5.210985, 
    5.244498, 5.27869, 5.311812, 5.34193, 5.367047, 5.385226, 5.394764, 
    5.394402, 5.383549, 5.362504, 5.332596, 5.296147, 5.256245, 5.216292, 
    5.179459,
  // totalHeight(10,3, 0-49)
    5.123564, 5.156494, 5.193518, 5.232036, 5.268888, 5.30088, 5.325299, 
    5.340286, 5.344973, 5.33944, 5.324524, 5.3016, 5.27236, 5.238668, 
    5.202416, 5.166353, 5.138496, 5.1065, 5.078358, 5.055256, 5.03751, 
    5.026891, 5.020802, 5.018765, 5.018983, 5.021102, 5.024645, 5.029631, 
    5.036055, 5.045497, 5.058444, 5.077137, 5.100204, 5.127726, 5.159303, 
    5.194069, 5.230758, 5.267785, 5.303344, 5.335496, 5.362273, 5.381793, 
    5.39242, 5.392964, 5.382909, 5.362636, 5.33356, 5.298093, 5.259374, 
    5.220767,
  // totalHeight(10,4, 0-49)
    5.148277, 5.183551, 5.220681, 5.256588, 5.288019, 5.312116, 5.326862, 
    5.331258, 5.325281, 5.309696, 5.285806, 5.25523, 5.219736, 5.181118, 
    5.141133, 5.102629, 5.075132, 5.042326, 5.01433, 4.99224, 4.976225, 
    4.968293, 4.965206, 4.966337, 4.969534, 4.974173, 4.979482, 4.985287, 
    4.991461, 4.999736, 5.010735, 5.027388, 5.048301, 5.073945, 5.104287, 
    5.138782, 5.176426, 5.215847, 5.255407, 5.293285, 5.327562, 5.356293, 
    5.377622, 5.389924, 5.392003, 5.383332, 5.364291, 5.336296, 5.301751, 
    5.263733,
  // totalHeight(10,5, 0-49)
    5.17261, 5.208737, 5.244016, 5.275208, 5.299335, 5.314187, 5.318586, 
    5.31239, 5.29629, 5.271561, 5.239791, 5.202709, 5.162052, 5.119503, 
    5.076645, 5.036462, 5.010109, 4.97695, 4.949606, 4.929027, 4.91522, 
    4.910427, 4.91076, 4.915475, 4.92213, 4.929779, 4.937321, 4.944317, 
    4.950469, 4.957533, 4.96622, 4.980175, 4.998003, 5.020619, 5.048433, 
    5.081285, 5.118479, 5.158883, 5.201038, 5.243255, 5.283694, 5.320426, 
    5.351492, 5.375001, 5.389269, 5.393025, 5.385661, 5.367476, 5.339813, 
    5.305001,
  // totalHeight(10,6, 0-49)
    5.194726, 5.230039, 5.261647, 5.286497, 5.302191, 5.307335, 5.301603, 
    5.285583, 5.260492, 5.227921, 5.189589, 5.147222, 5.102467, 5.056863, 
    5.011828, 4.97053, 4.945855, 4.912601, 4.886216, 4.867458, 4.85615, 
    4.854763, 4.858765, 4.867326, 4.877797, 4.888885, 4.899129, 4.907778, 
    4.914294, 4.920318, 4.926564, 4.9374, 4.951415, 4.97002, 4.994144, 
    5.024087, 5.059518, 5.099563, 5.142944, 5.188095, 5.233257, 5.276544, 
    5.315973, 5.349518, 5.375189, 5.391176, 5.396054, 5.389062, 5.370367, 
    5.341236,
  // totalHeight(10,7, 0-49)
    5.213053, 5.245964, 5.27248, 5.290026, 5.296961, 5.292734, 5.27777, 
    5.253204, 5.220595, 5.181672, 5.138168, 5.091727, 5.04387, 4.995987, 
    4.949328, 4.907313, 4.88458, 4.851351, 4.826089, 4.809305, 4.800615, 
    4.802724, 4.810457, 4.822952, 4.837451, 4.852314, 4.865723, 4.876563, 
    4.88401, 4.889411, 4.893355, 4.900923, 4.910622, 4.924387, 4.94375, 
    4.969565, 5.001939, 5.040301, 5.083554, 5.130239, 5.178657, 5.226962, 
    5.27318, 5.315236, 5.350972, 5.378225, 5.394969, 5.399563, 5.391072, 
    5.369621,
  // totalHeight(10,8, 0-49)
    5.226548, 5.255755, 5.276319, 5.286304, 5.284873, 5.272231, 5.249386, 
    5.217844, 5.179329, 5.135591, 5.088283, 5.038926, 4.98889, 4.939411, 
    4.891582, 4.849094, 4.828224, 4.795094, 4.771032, 4.756248, 4.750131, 
    4.755633, 4.766952, 4.783258, 4.801815, 4.820665, 4.837659, 4.851306, 
    4.860435, 4.865911, 4.868018, 4.872491, 4.877636, 4.885912, 4.899523, 
    4.919997, 4.947987, 4.983297, 5.02504, 5.071846, 5.122056, 5.173835, 
    5.225216, 5.274106, 5.318265, 5.355324, 5.38286, 5.39859, 5.40069, 
    5.388237,
  // totalHeight(10,9, 0-49)
    5.234836, 5.259479, 5.273821, 5.276622, 5.26777, 5.248077, 5.218955, 
    5.182111, 5.139313, 5.09224, 5.042422, 4.991228, 4.93987, 4.889423, 
    4.840813, 4.797938, 4.778379, 4.745469, 4.722646, 4.709779, 4.706027, 
    4.714598, 4.729111, 4.748862, 4.77128, 4.794157, 4.815078, 4.832183, 
    4.843925, 4.850475, 4.851599, 4.853556, 4.854271, 4.856665, 4.863659, 
    4.877585, 4.899804, 4.930608, 4.969382, 5.014863, 5.0654, 5.119133, 
    5.17407, 5.228092, 5.27892, 5.324071, 5.360898, 5.386709, 5.399065, 
    5.396215,
  // totalHeight(10,10, 0-49)
    5.238247, 5.257951, 5.266341, 5.262815, 5.247848, 5.222678, 5.188955, 
    5.148462, 5.102916, 5.053882, 5.002743, 4.950707, 4.898828, 4.848012, 
    4.798991, 4.755602, 4.736162, 4.703743, 4.682203, 4.671069, 4.66929, 
    4.68035, 4.697388, 4.71993, 4.745744, 4.772466, 4.797513, 4.818703, 
    4.834116, 4.843032, 4.844454, 4.844961, 4.841871, 4.838394, 4.838163, 
    4.844429, 4.859446, 4.88419, 4.918439, 4.961081, 5.01046, 5.064648, 
    5.121579, 5.17908, 5.234825, 5.286284, 5.330706, 5.365195, 5.38696, 
    5.393692,
  // totalHeight(10,11, 0-49)
    5.237722, 5.252574, 5.255694, 5.247005, 5.227397, 5.198365, 5.161659, 
    5.119038, 5.072123, 5.022343, 4.970935, 4.918961, 4.86732, 4.81674, 
    4.767717, 4.723385, 4.702055, 4.670654, 4.650481, 4.64079, 4.640394, 
    4.653071, 4.671667, 4.696053, 4.724506, 4.754633, 4.783804, 4.809594, 
    4.829752, 4.842523, 4.845928, 4.846569, 4.840914, 4.832191, 4.824595, 
    4.822354, 4.828823, 4.845907, 4.873978, 4.912177, 4.958867, 5.012014, 
    5.069425, 5.128822, 5.187816, 5.243847, 5.294146, 5.335773, 5.365799, 
    5.381611,
  // totalHeight(10,12, 0-49)
    5.234626, 5.245103, 5.243909, 5.231354, 5.20858, 5.177192, 5.138937, 
    5.095491, 5.048359, 4.998839, 4.948044, 4.896914, 4.84622, 4.796515, 
    4.748018, 4.701878, 4.675796, 4.646248, 4.627597, 4.618956, 4.619151, 
    4.632289, 4.651206, 4.676237, 4.706321, 4.739155, 4.772195, 4.802876, 
    4.828703, 4.846828, 4.854155, 4.856939, 4.85062, 4.838054, 4.82369, 
    4.812641, 4.809513, 4.817426, 4.837632, 4.869717, 4.912129, 4.962729, 
    5.019142, 5.078934, 5.139617, 5.198605, 5.253157, 5.300396, 5.33741, 
    5.361478,
  // totalHeight(10,13, 0-49)
    5.230535, 5.237388, 5.232965, 5.21782, 5.193212, 5.160748, 5.122097, 
    5.078829, 5.032333, 4.983805, 4.934273, 4.884608, 4.835494, 4.787343, 
    4.740097, 4.690714, 4.656355, 4.629813, 4.612917, 4.604844, 4.60468, 
    4.616896, 4.634736, 4.65907, 4.689609, 4.724247, 4.760649, 4.796208, 
    4.828288, 4.853024, 4.866192, 4.873289, 4.868722, 4.854521, 4.834921, 
    4.81561, 4.802438, 4.8, 4.810771, 4.835072, 4.871596, 4.918133, 4.972108, 
    5.030878, 5.091822, 5.152305, 5.209641, 5.261067, 5.303789, 5.335109,
  // totalHeight(10,14, 0-49)
    5.22699, 5.231134, 5.224566, 5.207964, 5.182598, 5.150006, 5.111754, 
    5.069297, 5.023933, 4.976803, 4.928903, 4.881094, 4.834053, 4.788131, 
    4.743088, 4.688396, 4.642111, 4.619964, 4.605116, 4.597078, 4.595531, 
    4.605345, 4.620689, 4.643006, 4.672795, 4.708239, 4.747289, 4.787376, 
    4.82584, 4.857959, 4.878545, 4.891905, 4.89165, 4.878604, 4.856218, 
    4.830238, 4.807499, 4.794166, 4.79429, 4.80929, 4.838372, 4.879369, 
    4.929523, 4.985952, 5.04586, 5.106551, 5.16538, 5.219721, 5.266939, 
    5.304432,
  // totalHeight(10,15, 0-49)
    5.225293, 5.227697, 5.219958, 5.202792, 5.177416, 5.145269, 5.107808, 
    5.066401, 5.02229, 4.976607, 4.930377, 4.88452, 4.839792, 4.79663, 
    4.75483, 4.69235, 4.631154, 4.614925, 4.602443, 4.593904, 4.58998, 
    4.595966, 4.607544, 4.62669, 4.65465, 4.689934, 4.730808, 4.7748, 
    4.819294, 4.85896, 4.887938, 4.908922, 4.915213, 4.906217, 4.884106, 
    4.854033, 4.823288, 4.799448, 4.788349, 4.792909, 4.813193, 4.847295, 
    4.892347, 4.94524, 5.002972, 5.062758, 5.12198, 5.17813, 5.228736, 
    5.271329,
  // totalHeight(10,16, 0-49)
    5.226336, 5.227925, 5.219817, 5.202703, 5.177724, 5.146221, 5.109568, 
    5.06908, 5.025991, 4.981462, 4.936589, 4.892404, 4.84983, 4.809532, 
    4.771629, 4.699264, 4.621652, 4.61295, 4.603134, 4.593575, 4.586397, 
    4.587306, 4.594104, 4.609207, 4.634496, 4.668808, 4.710706, 4.757823, 
    4.807619, 4.854417, 4.892068, 4.921228, 4.935552, 4.933044, 4.914313, 
    4.883314, 4.847099, 4.81419, 4.792173, 4.785765, 4.796284, 4.822381, 
    4.861237, 4.909564, 4.964163, 5.022121, 5.08082, 5.137845, 5.190862, 
    5.237532,
  // totalHeight(10,17, 0-49)
    5.230514, 5.23212, 5.224253, 5.207549, 5.183083, 5.152126, 5.116007, 
    5.076031, 5.033445, 4.989463, 4.945265, 4.902009, 4.860803, 4.822589, 
    4.787977, 4.705591, 4.612271, 4.612747, 4.605839, 4.594719, 4.583512, 
    4.578328, 4.579618, 4.590136, 4.612224, 4.645008, 4.687278, 4.736743, 
    4.790919, 4.844021, 4.890014, 4.927098, 4.949994, 4.955523, 4.94271, 
    4.913936, 4.875333, 4.835699, 4.804019, 4.7869, 4.787251, 4.804621, 
    4.836472, 4.879438, 4.930146, 4.985555, 5.04301, 5.100143, 5.154733, 
    5.204546,
  // totalHeight(10,18, 0-49)
    5.237718, 5.240082, 5.232924, 5.216834, 5.19283, 5.162156, 5.126127, 
    5.086053, 5.043212, 4.998859, 4.954231, 4.910549, 4.86899, 4.830619, 
    4.796376, 4.707914, 4.602833, 4.613844, 4.60993, 4.59652, 4.580455, 
    4.568354, 4.563672, 4.569397, 4.588124, 4.619167, 4.66143, 4.712628, 
    4.770273, 4.82866, 4.882247, 4.92637, 4.957467, 4.971514, 4.966166, 
    4.942143, 4.904187, 4.860658, 4.821369, 4.794617, 4.785073, 4.793501, 
    4.817908, 4.85501, 4.901318, 4.953671, 5.009349, 5.066003, 5.121474, 
    5.173612,
  // totalHeight(10,19, 0-49)
    5.247415, 5.251267, 5.245289, 5.230013, 5.20642, 5.175728, 5.139245, 
    5.098292, 5.054173, 5.008155, 4.961453, 4.915181, 4.870294, 4.827582, 
    4.788054, 4.702839, 4.595904, 4.617163, 4.615731, 4.598713, 4.576507, 
    4.556717, 4.545831, 4.546948, 4.562612, 4.592149, 4.634409, 4.687026, 
    4.747424, 4.810097, 4.870316, 4.920206, 4.958426, 4.980475, 4.982996, 
    4.965231, 4.930353, 4.885727, 4.841322, 4.806689, 4.788195, 4.788025, 
    4.80498, 4.836047, 4.87772, 4.926739, 4.980312, 5.036072, 5.091892, 
    5.14567,
  // totalHeight(10,20, 0-49)
    5.253863, 5.255918, 5.248505, 5.232355, 5.208736, 5.179231, 5.145556, 
    5.109469, 5.072702, 5.036943, 5.003791, 4.974656, 4.950539, 4.931577, 
    4.916345, 30, 4.529047, 4.533604, 4.533447, 4.529254, 4.524078, 4.517531, 
    4.516744, 4.524277, 4.543463, 4.574782, 4.617994, 4.671397, 4.732827, 
    4.797443, 4.86176, 4.91475, 4.957507, 4.985386, 4.994432, 4.982762, 
    4.952068, 4.908407, 4.861261, 4.820816, 4.794822, 4.786893, 4.796811, 
    4.82201, 4.859082, 4.904712, 4.956047, 5.010677, 5.066474, 5.121367,
  // totalHeight(10,21, 0-49)
    5.263675, 5.267076, 5.260616, 5.245088, 5.221847, 5.192562, 5.159019, 
    5.122997, 5.086214, 5.050299, 5.016766, 4.986938, 4.961788, 4.941614, 
    4.925509, 30, 4.57267, 4.567389, 4.555607, 4.539651, 4.524162, 4.505689, 
    4.496675, 4.498558, 4.514233, 4.543977, 4.587254, 4.642064, 4.705884, 
    4.773979, 4.843802, 4.901035, 4.949372, 4.984136, 5.000959, 4.997036, 
    4.972662, 4.932421, 4.884916, 4.840544, 4.808241, 4.793121, 4.796153, 
    4.815408, 4.847692, 4.889668, 4.938398, 4.991401, 5.046501, 5.101614,
  // totalHeight(10,22, 0-49)
    5.271476, 5.27575, 5.269802, 5.254496, 5.231293, 5.201962, 5.168361, 
    5.132299, 5.095483, 5.059496, 5.025783, 4.995612, 4.969961, 4.949296, 
    4.933185, 30, 4.606127, 4.593786, 4.574115, 4.550414, 4.528358, 4.500781, 
    4.48548, 4.482813, 4.495416, 4.523509, 4.566337, 4.621633, 4.686522, 
    4.756358, 4.829571, 4.888551, 4.939791, 4.978797, 5.001094, 5.003343, 
    4.984809, 4.94875, 4.902673, 4.85667, 4.820312, 4.799883, 4.797452, 
    4.8118, 4.840026, 4.878856, 4.925291, 4.976785, 5.031116, 5.086174,
  // totalHeight(10,23, 0-49)
    5.276399, 5.281113, 5.275375, 5.260115, 5.236866, 5.207469, 5.173829, 
    5.13778, 5.101011, 5.065071, 5.031356, 5.001098, 4.975291, 4.954518, 
    4.93868, 30, 4.630615, 4.613832, 4.58922, 4.560673, 4.534565, 4.500163, 
    4.480029, 4.473634, 4.483511, 4.509951, 4.552076, 4.607405, 4.672744, 
    4.743471, 4.818842, 4.878325, 4.930957, 4.972464, 4.998406, 5.005173, 
    4.991349, 4.959182, 4.915194, 4.868976, 4.830346, 4.80637, 4.800004, 
    4.810667, 4.83577, 4.87212, 4.916699, 4.966904, 5.020463, 5.075243,
  // totalHeight(10,24, 0-49)
    5.277895, 5.282643, 5.276915, 5.261662, 5.238444, 5.20912, 5.175599, 
    5.139707, 5.103124, 5.067368, 5.033813, 5.003671, 4.977938, 4.957258, 
    4.941692, 30, 4.644578, 4.625749, 4.598795, 4.567974, 4.540061, 4.501756, 
    4.478832, 4.470163, 4.478271, 4.503554, 4.545105, 4.600323, 4.665806, 
    4.736924, 4.813501, 4.87292, 4.926011, 4.96866, 4.996484, 5.005741, 
    4.994654, 4.964887, 4.922336, 4.876217, 4.836404, 4.810391, 4.801668, 
    4.810068, 4.83323, 4.868037, 4.911464, 4.96088, 5.013984, 5.068623,
  // totalHeight(10,25, 0-49)
    5.275751, 5.280137, 5.274252, 5.259029, 5.235986, 5.20693, 5.173734, 
    5.138188, 5.10195, 5.066529, 5.033287, 5.003433, 4.977952, 4.957484, 
    4.942075, 30, 4.646362, 4.627713, 4.600918, 4.57033, 4.542782, 4.504051, 
    4.480865, 4.47187, 4.479598, 4.504527, 4.545787, 4.600784, 4.666057, 
    4.736995, 4.813643, 4.872583, 4.925354, 4.967914, 4.995914, 5.005612, 
    4.995152, 4.966033, 4.923948, 4.877962, 4.837917, 4.81139, 4.802017, 
    4.809758, 4.832334, 4.866657, 4.909718, 4.958877, 5.011829, 5.066416,
  // totalHeight(10,26, 0-49)
    5.270087, 5.273705, 5.267471, 5.252261, 5.229498, 5.200881, 5.168194, 
    5.133167, 5.097431, 5.062489, 5.029718, 5.00033, 4.975293, 4.955161, 
    4.939804, 30, 4.636261, 4.619933, 4.595723, 4.567776, 4.542617, 4.506954, 
    4.486037, 4.478699, 4.487489, 4.512912, 4.554196, 4.60886, 4.67358, 
    4.743774, 4.819333, 4.877504, 4.92928, 4.970582, 4.997083, 5.005145, 
    4.993102, 4.962729, 4.919972, 4.874004, 4.834575, 4.809024, 4.800726, 
    4.809459, 4.832855, 4.867812, 4.911335, 4.960805, 5.013942, 5.0686,
  // totalHeight(10,27, 0-49)
    5.261351, 5.26376, 5.256897, 5.241565, 5.219057, 5.190928, 5.158837, 
    5.124437, 5.089321, 5.054998, 5.022872, 4.994169, 4.969829, 4.950259, 
    4.934984, 30, 4.616155, 4.604306, 4.585077, 4.56209, 4.541208, 4.511642, 
    4.495096, 4.490992, 4.501941, 4.528447, 4.569895, 4.624023, 4.687788, 
    4.756649, 4.829976, 4.887001, 4.937045, 4.975907, 4.999275, 5.003732, 
    4.988097, 4.954829, 4.910524, 4.864675, 4.826832, 4.803771, 4.798227, 
    4.809523, 4.835066, 4.871701, 4.916456, 4.966763, 5.020384, 5.0752,
  // totalHeight(10,28, 0-49)
    5.250287, 5.251001, 5.243098, 5.227319, 5.204828, 5.177031, 5.145455, 
    5.111665, 5.077218, 5.043633, 5.012346, 4.984618, 4.961354, 4.942771, 
    4.927911, 30, 4.589266, 4.58401, 4.572131, 4.556344, 4.541521, 4.520256, 
    4.509414, 4.509357, 4.5229, 4.55061, 4.592104, 4.645408, 4.707838, 
    4.774844, 4.844988, 4.900376, 4.947849, 4.983022, 5.001625, 5.000618, 
    4.979618, 4.942165, 4.895842, 4.850533, 4.815399, 4.796301, 4.795027, 
    4.81025, 4.839077, 4.87829, 4.924963, 4.976596, 5.031007, 5.086114,
  // totalHeight(10,29, 0-49)
    5.237892, 5.236384, 5.226872, 5.210082, 5.187092, 5.159198, 5.127821, 
    5.094449, 5.060609, 5.027836, 4.997607, 4.971239, 4.949625, 4.9328, 
    4.919292, 30, 4.557674, 4.560971, 4.558987, 4.552932, 4.546215, 4.534846, 
    4.530406, 4.534475, 4.550333, 4.578779, 4.61976, 4.671615, 4.73202, 
    4.796323, 4.862085, 4.914719, 4.958258, 4.988181, 5.000409, 4.992544, 
    4.965331, 4.923674, 4.876193, 4.832937, 4.80229, 4.788859, 4.793301, 
    4.813599, 4.846585, 4.889009, 4.938014, 4.991178, 5.046374, 5.101542,
  // totalHeight(10,30, 0-49)
    5.229731, 5.229138, 5.220243, 5.203627, 5.180113, 5.150661, 5.116294, 
    5.078084, 5.037141, 4.994608, 4.951617, 4.909244, 4.868432, 4.829989, 
    4.794954, 4.714292, 4.616234, 4.637926, 4.637839, 4.622587, 4.602194, 
    4.580849, 4.568728, 4.568097, 4.581463, 4.608438, 4.648096, 4.698241, 
    4.756376, 4.817419, 4.877771, 4.926244, 4.964109, 4.986963, 4.99125, 
    4.975613, 4.942276, 4.897612, 4.851018, 4.812195, 4.788252, 4.782269, 
    4.793753, 4.820078, 4.857902, 4.904008, 4.955632, 5.010437, 5.066337, 
    5.121289,
  // totalHeight(10,31, 0-49)
    5.219232, 5.216277, 5.205369, 5.187213, 5.162733, 5.132943, 5.098883, 
    5.061612, 5.022202, 4.98176, 4.94143, 4.902367, 4.865702, 4.832438, 
    4.803414, 4.719196, 4.623185, 4.63613, 4.634095, 4.622359, 4.607735, 
    4.594142, 4.588014, 4.591664, 4.607731, 4.635858, 4.675278, 4.723969, 
    4.779628, 4.836938, 4.891286, 4.934981, 4.966794, 4.982536, 4.979336, 
    4.957036, 4.91935, 4.873874, 4.830328, 4.797622, 4.781393, 4.783288, 
    4.801867, 4.834084, 4.87652, 4.926019, 4.979887, 5.035825, 5.091748, 
    5.145588,
  // totalHeight(10,32, 0-49)
    5.212204, 5.207666, 5.195166, 5.175536, 5.149817, 5.119109, 5.084501, 
    5.047058, 5.007833, 4.967883, 4.928288, 4.890134, 4.854459, 4.822115, 
    4.793561, 4.715725, 4.631017, 4.635134, 4.631091, 4.622012, 4.61214, 
    4.605616, 4.605232, 4.613331, 4.632458, 4.662114, 4.70151, 4.748676, 
    4.801376, 4.854101, 4.901446, 4.939006, 4.963384, 4.970959, 4.959958, 
    4.931739, 4.891537, 4.847791, 4.809901, 4.785426, 4.77831, 4.788849, 
    4.814866, 4.853093, 4.900144, 4.952962, 5.008929, 5.065755, 5.121329, 
    5.173527,
  // totalHeight(10,33, 0-49)
    5.20914, 5.203825, 5.190194, 5.169207, 5.142048, 5.109946, 5.074082, 
    5.035568, 4.995455, 4.954757, 4.914469, 4.875549, 4.838848, 4.804925, 
    4.77372, 4.706617, 4.637273, 4.633828, 4.628059, 4.621222, 4.615577, 
    4.615524, 4.620589, 4.633079, 4.655277, 4.686444, 4.725629, 4.770813, 
    4.819751, 4.866857, 4.906264, 4.936515, 4.952563, 4.951732, 4.933675, 
    4.901386, 4.861358, 4.822259, 4.792506, 4.777924, 4.780762, 4.800201, 
    4.83359, 4.877619, 4.929025, 4.984875, 5.042601, 5.0999, 5.154591, 
    5.204463,
  // totalHeight(10,34, 0-49)
    5.210141, 5.204962, 5.190825, 5.168797, 5.140215, 5.106468, 5.068875, 
    5.028635, 4.986836, 4.944474, 4.902484, 4.861712, 4.82285, 4.786231, 
    4.751455, 4.695054, 4.642087, 4.632432, 4.625143, 4.620174, 4.618269, 
    4.623944, 4.634017, 4.650625, 4.67562, 4.707963, 4.746448, 4.788954, 
    4.833173, 4.873645, 4.904438, 4.926645, 4.934232, 4.925783, 4.902545, 
    4.868981, 4.83229, 4.800661, 4.780991, 4.77725, 4.790213, 4.818267, 
    4.858552, 4.907861, 4.963102, 5.021472, 5.080428, 5.137609, 5.190722, 
    5.237449,
  // totalHeight(10,35, 0-49)
    5.214813, 5.2108, 5.196992, 5.174516, 5.144845, 5.109542, 5.070085, 
    5.0278, 4.983854, 4.939272, 4.894969, 4.851746, 4.810218, 4.770653, 
    4.732632, 4.684653, 4.646751, 4.632051, 4.62333, 4.619743, 4.620919, 
    4.631336, 4.64574, 4.665937, 4.693183, 4.726111, 4.763205, 4.802227, 
    4.84081, 4.873873, 4.895854, 4.909962, 4.909899, 4.895682, 4.870054, 
    4.838493, 4.808202, 4.78625, 4.777755, 4.784982, 4.807583, 4.843489, 
    4.889846, 4.943633, 5.00196, 5.062129, 5.121593, 5.177893, 5.228593, 
    5.271242,
  // totalHeight(10,36, 0-49)
    5.222264, 5.220515, 5.208066, 5.186024, 5.155957, 5.119577, 5.078528, 
    5.03429, 4.988141, 4.941181, 4.894366, 4.848512, 4.804265, 4.76197, 
    4.721433, 4.679046, 4.653185, 4.63448, 4.62433, 4.621491, 4.624862, 
    4.638769, 4.656545, 4.67952, 4.708213, 4.740936, 4.775853, 4.810642, 
    4.842913, 4.868268, 4.881892, 4.888682, 4.882713, 4.865387, 4.840581, 
    4.814148, 4.792623, 4.781571, 4.784374, 4.801928, 4.833148, 4.875787, 
    4.927128, 4.984381, 5.044846, 5.105902, 5.164972, 5.219464, 5.266778, 
    5.30433,
  // totalHeight(10,37, 0-49)
    5.231169, 5.232775, 5.222847, 5.202373, 5.172933, 5.13634, 5.094387, 
    5.048704, 5.000711, 4.951622, 4.902481, 4.854186, 4.807487, 4.762895, 
    4.720541, 4.681284, 4.663596, 4.641848, 4.63024, 4.627433, 4.631958, 
    4.647927, 4.667863, 4.692542, 4.721674, 4.753293, 4.785275, 4.815282, 
    4.840997, 4.858955, 4.865395, 4.866431, 4.85696, 4.839487, 4.818485, 
    4.799541, 4.78807, 4.788061, 4.801427, 4.82809, 4.86656, 4.914594, 
    4.969669, 5.029223, 5.090712, 5.15157, 5.209159, 5.260755, 5.303586, 
    5.334973,
  // totalHeight(10,38, 0-49)
    5.239892, 5.24584, 5.239644, 5.222045, 5.194521, 5.158906, 5.117092, 
    5.070849, 5.021742, 4.971128, 4.920183, 4.869933, 4.821266, 4.774899, 
    4.73128, 4.693408, 4.680095, 4.656179, 4.643091, 4.639637, 4.644267, 
    4.660845, 4.6816, 4.706756, 4.735232, 4.764845, 4.793278, 4.818267, 
    4.837685, 4.849177, 4.850168, 4.847516, 4.837119, 4.822165, 4.80716, 
    4.796963, 4.795705, 4.805967, 4.828554, 4.862772, 4.906951, 4.958941, 
    5.016412, 5.076992, 5.138256, 5.197663, 5.252513, 5.29996, 5.337116, 
    5.361272,
  // totalHeight(10,39, 0-49)
    5.246655, 5.257724, 5.256416, 5.243073, 5.218928, 5.18572, 5.145367, 
    5.099737, 5.050538, 4.999286, 4.947315, 4.895807, 4.845814, 4.798248, 
    4.753822, 4.71631, 4.704317, 4.678978, 4.664438, 4.659803, 4.663629, 
    4.679513, 4.699796, 4.724214, 4.750978, 4.777809, 4.802306, 4.822383, 
    4.83622, 4.842612, 4.840141, 4.835948, 4.826879, 4.816355, 4.808491, 
    4.8072, 4.815392, 4.83454, 4.864683, 4.904767, 4.953069, 5.007549, 
    5.066037, 5.126289, 5.185953, 5.242501, 5.293189, 5.335102, 5.365329, 
    5.381271,
  // totalHeight(10,40, 0-49)
    5.249744, 5.266394, 5.270947, 5.263197, 5.243958, 5.214726, 5.177338, 
    5.133704, 5.085651, 5.034855, 4.982824, 4.930913, 4.880349, 4.832219, 
    4.787439, 4.749863, 4.737173, 4.711016, 4.69513, 4.68898, 4.691325, 
    4.705497, 4.724216, 4.746839, 4.771021, 4.794501, 4.81493, 4.830498, 
    4.839759, 4.842586, 4.838536, 4.834641, 4.828501, 4.823401, 4.822832, 
    4.829747, 4.846045, 4.872379, 4.908298, 4.952549, 5.003408, 5.058919, 
    5.117007, 5.175501, 5.232083, 5.284229, 5.329195, 5.364105, 5.386174, 
    5.393111,
  // totalHeight(10,41, 0-49)
    5.247719, 5.269979, 5.281053, 5.280043, 5.267168, 5.243511, 5.210688, 
    5.170568, 5.125053, 5.075967, 5.024994, 4.973671, 4.923398, 4.875422, 
    4.830817, 4.79321, 4.778804, 4.752316, 4.735268, 4.727466, 4.727908, 
    4.739669, 4.756018, 4.776052, 4.797035, 4.816849, 4.833313, 4.844961, 
    4.85074, 4.851439, 4.847338, 4.845059, 4.842711, 4.843216, 4.849365, 
    4.863264, 4.886032, 4.917758, 4.95768, 5.004436, 5.056305, 5.111372, 
    5.167601, 5.222831, 5.274746, 5.320846, 5.358463, 5.384906, 5.397736, 
    5.395216,
  // totalHeight(10,42, 0-49)
    5.239619, 5.267014, 5.284798, 5.291317, 5.286037, 5.269451, 5.242799, 
    5.207787, 5.166325, 5.120343, 5.071693, 5.02209, 4.973096, 4.926105, 
    4.88232, 4.845045, 4.828703, 4.802299, 4.784326, 4.774885, 4.773208, 
    4.78215, 4.795608, 4.812541, 4.829976, 4.846041, 4.858818, 4.867209, 
    4.870528, 4.870278, 4.867199, 4.867313, 4.869003, 4.87472, 4.886584, 
    4.906005, 4.933528, 4.968866, 5.01106, 5.058681, 5.109999, 5.1631, 
    5.215928, 5.266298, 5.311891, 5.350265, 5.378949, 5.395628, 5.398466, 
    5.386536,
  // totalHeight(10,43, 0-49)
    5.225125, 5.256631, 5.280723, 5.295022, 5.298166, 5.289894, 5.270908, 
    5.242608, 5.206801, 5.165462, 5.120562, 5.073971, 5.027399, 4.982369, 
    4.940185, 4.903838, 4.885886, 4.85994, 4.841307, 4.830328, 4.826455, 
    4.832383, 4.842665, 4.856229, 4.869998, 4.882415, 4.891881, 4.897665, 
    4.899386, 4.899063, 4.897659, 4.900507, 4.90607, 4.916288, 4.932685, 
    4.956121, 4.986723, 5.023946, 5.066707, 5.113532, 5.16267, 5.212178, 
    5.259955, 5.303786, 5.34137, 5.370416, 5.388793, 5.394788, 5.38742, 
    5.366787,
  // totalHeight(10,44, 0-49)
    5.204635, 5.238729, 5.268057, 5.289697, 5.30149, 5.302343, 5.292276, 
    5.272214, 5.243718, 5.20869, 5.169145, 5.127045, 5.08421, 5.042264, 
    5.0026, 4.967926, 4.949046, 4.92391, 4.904885, 4.892501, 4.88643, 
    4.88929, 4.896282, 4.906398, 4.916552, 4.925547, 4.932125, 4.93589, 
    4.936687, 4.936886, 4.937493, 4.94312, 4.952159, 4.966044, 4.985777, 
    5.011779, 5.043863, 5.081303, 5.122929, 5.167236, 5.212452, 5.256604, 
    5.297564, 5.333117, 5.361072, 5.379413, 5.386541, 5.381553, 5.364513, 
    5.336632,
  // totalHeight(10,45, 0-49)
    5.179212, 5.214012, 5.246877, 5.274645, 5.294554, 5.304733, 5.304421, 
    5.293918, 5.274354, 5.247395, 5.214958, 5.179004, 5.14139, 5.103791, 
    5.067675, 5.035524, 5.016601, 4.992625, 4.973468, 4.959824, 4.951601, 
    4.951439, 4.955157, 4.961893, 4.9686, 4.974474, 4.978585, 4.980832, 
    4.981196, 4.982283, 4.985005, 4.993274, 5.005284, 5.021986, 5.043922, 
    5.071142, 5.103206, 5.139245, 5.178025, 5.218019, 5.257449, 5.294353, 
    5.326642, 5.352213, 5.369123, 5.375821, 5.371424, 5.355994, 5.330694, 
    5.29772,
  // totalHeight(10,46, 0-49)
    5.15041, 5.183906, 5.218145, 5.250115, 5.276795, 5.295731, 5.305416, 
    5.305406, 5.296213, 5.27905, 5.255547, 5.227502, 5.196701, 5.164815, 
    5.133346, 5.104626, 5.08668, 5.064239, 5.04522, 5.03049, 5.020214, 
    5.017181, 5.017759, 5.021304, 5.024827, 5.027922, 5.029962, 5.031085, 
    5.031336, 5.033477, 5.038228, 5.048871, 5.063292, 5.081979, 5.10506, 
    5.132253, 5.162891, 5.19597, 5.230196, 5.264036, 5.295753, 5.323472, 
    5.345274, 5.359347, 5.364205, 5.358969, 5.343636, 5.319263, 5.287948, 
    5.25254,
  // totalHeight(10,47, 0-49)
    5.119985, 5.150326, 5.183611, 5.217366, 5.248749, 5.275069, 5.294239, 
    5.305062, 5.307268, 5.30139, 5.288529, 5.270121, 5.247734, 5.222944, 
    5.197252, 5.1729, 5.157071, 5.136595, 5.11804, 5.102479, 5.090351, 
    5.084734, 5.082446, 5.08311, 5.083791, 5.084471, 5.08479, 5.085076, 
    5.085362, 5.088531, 5.095047, 5.107666, 5.123862, 5.143695, 5.166904, 
    5.192897, 5.220782, 5.249414, 5.27744, 5.303342, 5.32549, 5.342224, 
    5.351979, 5.353467, 5.345912, 5.329299, 5.304561, 5.273603, 5.239101, 
    5.204047,
  // totalHeight(10,48, 0-49)
    5.089595, 5.115337, 5.145545, 5.178566, 5.212147, 5.243782, 5.271115, 
    5.29231, 5.306252, 5.312603, 5.311698, 5.304386, 5.291848, 5.275453, 
    5.25664, 5.23762, 5.225192, 5.207209, 5.189566, 5.173572, 5.159956, 
    5.152224, 5.147508, 5.145734, 5.143994, 5.142636, 5.141529, 5.141139, 
    5.141435, 5.145405, 5.153227, 5.167259, 5.184483, 5.204558, 5.226863, 
    5.250508, 5.274375, 5.297177, 5.317502, 5.333895, 5.344922, 5.349295, 
    5.346019, 5.33458, 5.315123, 5.288604, 5.256801, 5.222151, 5.187412, 
    5.155191,
  // totalHeight(10,49, 0-49)
    5.053679, 5.072524, 5.096591, 5.125384, 5.157755, 5.191944, 5.225796, 
    5.257071, 5.283777, 5.304451, 5.318295, 5.325191, 5.325613, 5.320494, 
    5.311103, 5.300251, 5.299141, 5.285053, 5.268355, 5.251288, 5.235315, 
    5.227765, 5.223431, 5.222784, 5.22031, 5.217353, 5.213843, 5.210539, 
    5.206765, 5.208167, 5.214479, 5.229855, 5.247833, 5.267559, 5.287977, 
    5.307836, 5.32576, 5.340317, 5.350102, 5.353841, 5.350516, 5.339516, 
    5.320797, 5.295008, 5.263525, 5.228363, 5.191968, 5.156848, 5.125219, 
    5.098701,
  // totalHeight(11,0, 0-49)
    5.173462, 5.206308, 5.240257, 5.272574, 5.300474, 5.321579, 5.334246, 
    5.337715, 5.33208, 5.318138, 5.297173, 5.270765, 5.240604, 5.208375, 
    5.175654, 5.144077, 5.116427, 5.090436, 5.068562, 5.051296, 5.038685, 
    5.030923, 5.027062, 5.026567, 5.028524, 5.032345, 5.037494, 5.043713, 
    5.050945, 5.059712, 5.070448, 5.084126, 5.100892, 5.121141, 5.144976, 
    5.172139, 5.202004, 5.233603, 5.265666, 5.296687, 5.325003, 5.348888, 
    5.366683, 5.376942, 5.378628, 5.371307, 5.355311, 5.331816, 5.302765, 
    5.270608,
  // totalHeight(11,1, 0-49)
    5.194742, 5.228152, 5.26071, 5.289646, 5.312393, 5.32699, 5.332311, 
    5.328114, 5.314935, 5.29389, 5.266475, 5.234376, 5.199319, 5.162972, 
    5.126867, 5.092795, 5.064954, 5.037652, 5.015035, 4.997619, 4.985379, 
    4.97889, 4.976613, 4.977965, 4.981647, 4.987005, 4.993341, 5.000309, 
    5.007703, 5.0163, 5.026547, 5.039942, 5.056371, 5.076459, 5.100532, 
    5.128533, 5.160006, 5.194112, 5.229676, 5.265248, 5.299183, 5.329723, 
    5.355093, 5.373639, 5.383974, 5.385177, 5.376961, 5.359829, 5.335091, 
    5.304753,
  // totalHeight(11,2, 0-49)
    5.215133, 5.247335, 5.276393, 5.299809, 5.315543, 5.322279, 5.319528, 
    5.307566, 5.287278, 5.259983, 5.227242, 5.190721, 5.152076, 5.112883, 
    5.074576, 5.039062, 5.011899, 4.983998, 4.961249, 4.944171, 4.93268, 
    4.927715, 4.927212, 4.93057, 4.936181, 4.943317, 4.951117, 4.959096, 
    4.966879, 4.975387, 4.985026, 4.997762, 5.013227, 5.032263, 5.055445, 
    5.082962, 5.114574, 5.149624, 5.187086, 5.225627, 5.263697, 5.299596, 
    5.33156, 5.357855, 5.376884, 5.387331, 5.388323, 5.37959, 5.3616, 5.335593,
  // totalHeight(11,3, 0-49)
    5.23278, 5.262092, 5.285949, 5.302372, 5.310034, 5.308362, 5.297498, 
    5.278173, 5.251532, 5.218977, 5.182038, 5.142278, 5.101216, 5.060287, 
    5.020789, 4.984736, 4.959036, 4.931108, 4.908727, 4.892389, 4.881948, 
    4.878703, 4.880101, 4.885571, 4.893275, 4.902404, 4.911927, 4.921201, 
    4.929637, 4.9382, 4.947193, 4.959, 4.972971, 4.990158, 5.011407, 
    5.037199, 5.067567, 5.102092, 5.139944, 5.17996, 5.220726, 5.260663, 
    5.298082, 5.331253, 5.358465, 5.378115, 5.388823, 5.389595, 5.380008, 
    5.360395,
  // totalHeight(11,4, 0-49)
    5.246124, 5.271151, 5.28868, 5.297393, 5.296728, 5.286824, 5.26838, 
    5.242476, 5.21042, 5.173625, 5.133534, 5.091561, 5.049062, 5.007304, 
    4.967432, 4.931567, 4.908005, 4.880484, 4.858866, 4.843581, 4.83441, 
    4.833011, 4.836378, 4.843999, 4.853899, 4.86519, 4.876671, 4.887522, 
    4.896918, 4.905757, 4.914163, 4.924904, 4.936983, 4.951648, 4.970031, 
    4.992957, 5.020799, 5.053441, 5.090303, 5.130426, 5.172563, 5.215267, 
    5.256948, 5.295912, 5.330392, 5.358579, 5.378705, 5.389174, 5.388783, 
    5.376987,
  // totalHeight(11,5, 0-49)
    5.254175, 5.273928, 5.284616, 5.285609, 5.277045, 5.259663, 5.234583, 
    5.203132, 5.1667, 5.126667, 5.08436, 5.041042, 4.997897, 4.956021, 
    4.916396, 4.881262, 4.860361, 4.83355, 4.812981, 4.798963, 4.791189, 
    4.79168, 4.796989, 4.80671, 4.818825, 4.832373, 4.846004, 4.858711, 
    4.86942, 4.878846, 4.88686, 4.896566, 4.906542, 4.918179, 4.932914, 
    4.951959, 4.976102, 5.005606, 5.040208, 5.079185, 5.121468, 5.165733, 
    5.210474, 5.254028, 5.294588, 5.330204, 5.358836, 5.378459, 5.387281, 
    5.384035,
  // totalHeight(11,6, 0-49)
    5.256631, 5.270588, 5.274484, 5.268309, 5.25277, 5.229043, 5.198534, 
    5.162709, 5.122982, 5.080671, 5.036992, 4.993062, 4.949906, 4.90846, 
    4.869534, 4.835497, 4.817565, 4.791654, 4.772311, 4.759662, 4.753291, 
    4.755591, 4.762683, 4.77432, 4.788547, 4.804348, 4.820257, 4.835084, 
    4.847507, 4.857955, 4.865939, 4.874877, 4.882786, 4.891138, 4.901649, 
    4.915957, 4.935346, 4.960551, 4.991693, 5.028335, 5.069591, 5.114242, 
    5.160832, 5.2077, 5.252995, 5.294673, 5.33052, 5.358258, 5.375719, 
    5.381134,
  // totalHeight(11,7, 0-49)
    5.253899, 5.261981, 5.259573, 5.247164, 5.225865, 5.197128, 5.162515, 
    5.123538, 5.081592, 5.037923, 4.993641, 4.949739, 4.907105, 4.866518, 
    4.828615, 4.795863, 4.780922, 4.756021, 4.737971, 4.726662, 4.721548, 
    4.72541, 4.733949, 4.747142, 4.763211, 4.781125, 4.799346, 4.816528, 
    4.831117, 4.843144, 4.851673, 4.860385, 4.866592, 4.871735, 4.877743, 
    4.88669, 4.900416, 4.920234, 4.94675, 4.979874, 5.018923, 5.062773, 
    5.109976, 5.158839, 5.207454, 5.253706, 5.295303, 5.329849, 5.355006, 
    5.36871,
  // totalHeight(11,8, 0-49)
    5.246972, 5.249469, 5.241543, 5.224041, 5.198316, 5.165953, 5.128552, 
    5.087615, 5.044479, 5.000314, 4.956141, 4.912849, 4.871207, 4.831842, 
    4.795206, 4.763745, 4.751428, 4.727627, 4.710842, 4.700696, 4.696517, 
    4.701485, 4.710924, 4.725105, 4.742551, 4.762268, 4.782706, 4.802408, 
    4.81963, 4.83391, 4.843769, 4.853097, 4.858361, 4.860801, 4.86244, 
    4.865728, 4.873104, 4.886553, 4.907292, 4.935679, 4.971288, 5.01309, 
    5.059626, 5.109141, 5.159651, 5.208991, 5.254846, 5.29482, 5.326542, 
    5.347835,
  // totalHeight(11,9, 0-49)
    5.237248, 5.234728, 5.222235, 5.200835, 5.17199, 5.1373, 5.09833, 
    5.056515, 5.013119, 4.96924, 4.925823, 4.883679, 4.843467, 4.805668, 
    4.770514, 4.740153, 4.729591, 4.707032, 4.691422, 4.682123, 4.678374, 
    4.683771, 4.693341, 4.707723, 4.725875, 4.746894, 4.769297, 4.791569, 
    4.811847, 4.829095, 4.841227, 4.852277, 4.857747, 4.858494, 4.856425, 
    4.854231, 4.854913, 4.861206, 4.875076, 4.897473, 4.92833, 4.966763, 
    5.011302, 5.060114, 5.111127, 5.162135, 5.210836, 5.254894, 5.292007, 
    5.319999,
  // totalHeight(11,10, 0-49)
    5.226325, 5.219534, 5.203464, 5.179299, 5.148501, 5.112608, 5.073096, 
    5.031306, 4.988426, 4.94549, 4.903389, 4.862872, 4.824508, 4.788627, 
    4.755206, 4.725522, 4.715262, 4.694233, 4.679683, 4.670805, 4.666822, 
    4.671776, 4.680524, 4.694141, 4.712152, 4.733792, 4.757727, 4.782455, 
    4.806074, 4.826941, 4.84233, 4.856339, 4.863483, 4.86403, 4.859515, 
    4.852623, 4.846785, 4.845483, 4.851567, 4.866756, 4.891508, 4.925184, 
    4.966353, 5.013109, 5.063296, 5.114656, 5.164914, 5.211822, 5.253187, 
    5.286903,
  // totalHeight(11,11, 0-49)
    5.215777, 5.205538, 5.186835, 5.160881, 5.129076, 5.092853, 5.05357, 
    5.01247, 4.970669, 4.929159, 4.888799, 4.850304, 4.814176, 4.780593, 
    4.749253, 4.719546, 4.70758, 4.688578, 4.67502, 4.666077, 4.661113, 
    4.664628, 4.671499, 4.683293, 4.700191, 4.72163, 4.746493, 4.773363, 
    4.800385, 4.825321, 4.844834, 4.86298, 4.873383, 4.875564, 4.870417, 
    4.860304, 4.848796, 4.840018, 4.837758, 4.844696, 4.862033, 4.889554, 
    4.925972, 4.969349, 5.01745, 5.067966, 5.118637, 5.167293, 5.211854, 
    5.250307,
  // totalHeight(11,12, 0-49)
    5.206971, 5.194101, 5.173579, 5.146593, 5.114454, 5.078471, 5.039887, 
    4.99986, 4.959449, 4.919629, 4.88126, 4.845059, 4.811492, 4.78062, 
    4.751868, 4.72114, 4.705098, 4.688858, 4.676319, 4.666856, 4.660173, 
    4.661228, 4.665177, 4.674097, 4.688881, 4.709216, 4.734272, 4.762765, 
    4.792983, 4.822137, 4.846368, 4.869545, 4.884646, 4.890373, 4.886761, 
    4.875495, 4.859918, 4.844513, 4.833935, 4.83196, 4.84078, 4.860842, 
    4.891177, 4.929914, 4.974764, 5.023362, 5.073436, 5.12287, 5.169671, 
    5.211904,
  // totalHeight(11,13, 0-49)
    5.200899, 5.186135, 5.164429, 5.136922, 5.104827, 5.069341, 5.031617, 
    4.992749, 4.953773, 4.915673, 4.879345, 4.845548, 4.814764, 4.787011, 
    4.761545, 4.728561, 4.7061, 4.693552, 4.682205, 4.671872, 4.662838, 
    4.660499, 4.66059, 4.665687, 4.677411, 4.695735, 4.72017, 4.749611, 
    4.782543, 4.815727, 4.844905, 4.873561, 4.8944, 4.905334, 4.90543, 
    4.895422, 4.878002, 4.857599, 4.839486, 4.828537, 4.828136, 4.839681, 
    4.862757, 4.895705, 4.936254, 4.981984, 5.030586, 5.079952, 5.128131, 
    5.173246,
  // totalHeight(11,14, 0-49)
    5.198095, 5.182048, 5.159592, 5.13182, 5.099866, 5.064854, 5.027873, 
    4.989992, 4.952253, 4.915678, 4.881233, 4.849756, 4.82182, 4.797526, 
    4.776157, 4.739671, 4.70902, 4.701211, 4.69137, 4.679989, 4.668147, 
    4.661624, 4.657088, 4.65757, 4.665394, 4.680862, 4.703853, 4.733477, 
    4.768441, 4.805169, 4.839162, 4.873245, 4.9003, 4.917571, 4.923186, 
    4.916782, 4.900061, 4.876922, 4.852844, 4.83361, 4.823883, 4.826264, 
    4.841175, 4.867381, 4.902731, 4.944778, 4.991159, 5.039723, 5.088521, 
    5.135692,
  // totalHeight(11,15, 0-49)
    5.198611, 5.181742, 5.158781, 5.130789, 5.098861, 5.064082, 5.027527, 
    4.990268, 4.953382, 4.917949, 4.885024, 4.855564, 4.83031, 4.809587, 
    4.793001, 4.752295, 4.712822, 4.710817, 4.702914, 4.690477, 4.67556, 
    4.664219, 4.654443, 4.649671, 4.652883, 4.664748, 4.685534, 4.714571, 
    4.750784, 4.790377, 4.82878, 4.867803, 4.900972, 4.92504, 4.93734, 
    4.936428, 4.922827, 4.899501, 4.871641, 4.845568, 4.827119, 4.820251, 
    4.826494, 4.845283, 4.874737, 4.912448, 4.955987, 5.003134, 5.051886, 
    5.100367,
  // totalHeight(11,16, 0-49)
    5.202085, 5.184723, 5.161361, 5.133057, 5.10091, 5.066013, 5.029459, 
    4.99235, 4.955808, 4.920977, 4.889006, 4.860992, 4.837896, 4.820388, 
    4.808672, 4.76449, 4.717262, 4.722044, 4.716553, 4.703173, 4.685042, 
    4.668344, 4.652804, 4.642239, 4.640246, 4.647893, 4.665833, 4.693597, 
    4.730288, 4.771996, 4.814262, 4.857442, 4.896148, 4.926826, 4.946223, 
    4.951967, 4.943392, 4.922285, 4.893093, 4.862197, 4.836313, 4.820743, 
    4.818316, 4.829373, 4.852494, 4.885402, 4.925627, 4.970856, 5.019004, 
    5.068143,
  // totalHeight(11,17, 0-49)
    5.207882, 5.190274, 5.166554, 5.137811, 5.105181, 5.069798, 5.032796, 
    4.995312, 4.95851, 4.923584, 4.891758, 4.864257, 4.842258, 4.826826, 
    4.818871, 4.77463, 4.723094, 4.735348, 4.732672, 4.718445, 4.696949, 
    4.674356, 4.652512, 4.635655, 4.627968, 4.630945, 4.645575, 4.671546, 
    4.708066, 4.751193, 4.796754, 4.843171, 4.886521, 4.923114, 4.949328, 
    4.962093, 4.959697, 4.942693, 4.914481, 4.881027, 4.849508, 4.826371, 
    4.815795, 4.819218, 4.835872, 4.863728, 4.900331, 4.943276, 4.990375, 
    5.039623,
  // totalHeight(11,18, 0-49)
    5.215275, 5.197681, 5.173691, 5.144443, 5.111129, 5.074939, 5.037043, 
    4.998607, 4.960812, 4.924872, 4.892043, 4.863613, 4.840909, 4.825321, 
    4.818491, 4.781203, 4.73237, 4.751977, 4.752251, 4.737044, 4.711777, 
    4.682581, 4.653769, 4.630121, 4.616386, 4.614459, 4.625572, 4.649482, 
    4.685395, 4.729392, 4.777759, 4.826488, 4.873441, 4.914927, 4.947153, 
    4.966595, 4.970727, 4.958978, 4.933579, 4.899727, 4.8646, 4.835458, 
    4.817726, 4.814026, 4.824396, 4.847192, 4.880045, 4.920485, 4.966215, 
    5.015142,
  // totalHeight(11,19, 0-49)
    5.223647, 5.206471, 5.182448, 5.152765, 5.118663, 5.081373, 5.042089, 
    5.001988, 4.962242, 4.924037, 4.888577, 4.857102, 4.830956, 4.811839, 
    4.802468, 4.782428, 4.748799, 4.774101, 4.776849, 4.759989, 4.72988, 
    4.692934, 4.656215, 4.62528, 4.605374, 4.598666, 4.606437, 4.628368, 
    4.663541, 4.708077, 4.758886, 4.809097, 4.858589, 4.903782, 4.940869, 
    4.966106, 4.976411, 4.9703, 4.948884, 4.916395, 4.87963, 4.846251, 
    4.822695, 4.812732, 4.817303, 4.835267, 4.864427, 4.902291, 4.94647, 
    4.994776,
  // totalHeight(11,20, 0-49)
    5.228605, 5.209377, 5.183713, 5.153066, 5.118945, 5.08285, 5.046243, 
    5.010551, 4.977164, 4.947405, 4.922451, 4.903156, 4.889757, 4.881487, 
    4.876232, 30, 4.74619, 4.746288, 4.737542, 4.720608, 4.697607, 4.668127, 
    4.638677, 4.612827, 4.595506, 4.58938, 4.596458, 4.617135, 4.651025, 
    4.694868, 4.746641, 4.79661, 4.846766, 4.893705, 4.933717, 4.963015, 
    4.978206, 4.977147, 4.959987, 4.929938, 4.893122, 4.857208, 4.829299, 
    4.814166, 4.813659, 4.827224, 4.852918, 4.888282, 4.930861, 4.978384,
  // totalHeight(11,21, 0-49)
    5.2353, 5.216488, 5.190962, 5.160259, 5.125952, 5.089577, 5.052596, 
    5.016393, 4.982272, 4.951435, 4.92492, 4.903454, 4.887238, 4.875626, 
    4.866798, 30, 4.797721, 4.792305, 4.77688, 4.75208, 4.720561, 4.678942, 
    4.639472, 4.605354, 4.581752, 4.571404, 4.576097, 4.595869, 4.629888, 
    4.674782, 4.72919, 4.780305, 4.832267, 4.881819, 4.925358, 4.959108, 
    4.979494, 4.983882, 4.97161, 4.944922, 4.909168, 4.871809, 4.840419, 
    4.820678, 4.815356, 4.824558, 4.846657, 4.879263, 4.919861, 4.966089,
  // totalHeight(11,22, 0-49)
    5.239971, 5.221348, 5.19583, 5.165015, 5.130526, 5.093925, 5.056665, 
    5.020096, 4.985459, 4.95387, 4.926275, 4.903344, 4.885296, 4.871654, 
    4.860947, 30, 4.835303, 4.825794, 4.806291, 4.777096, 4.740961, 4.690882, 
    4.644479, 4.604306, 4.575753, 4.561767, 4.564087, 4.582548, 4.615982, 
    4.660958, 4.716836, 4.767711, 4.819979, 4.870557, 4.915993, 4.952604, 
    4.976768, 4.985557, 4.977713, 4.954643, 4.920895, 4.883494, 4.850173, 
    4.82724, 4.818252, 4.823944, 4.84304, 4.873272, 4.912107, 4.957114,
  // totalHeight(11,23, 0-49)
    5.242476, 5.223934, 5.198411, 5.167542, 5.132972, 5.096276, 5.058898, 
    5.022161, 4.987256, 4.95525, 4.927035, 4.903254, 4.884159, 4.869406, 
    4.857812, 30, 4.860757, 4.848539, 4.826694, 4.795172, 4.756673, 4.700799, 
    4.649669, 4.605175, 4.572934, 4.556139, 4.556563, 4.573909, 4.606749, 
    4.651597, 4.708432, 4.75862, 4.810601, 4.861441, 4.90783, 4.9462, 
    4.97295, 4.984998, 4.980686, 4.960799, 4.929197, 4.892447, 4.858245, 
    4.833289, 4.82172, 4.824795, 4.841565, 4.869889, 4.907241, 4.951149,
  // totalHeight(11,24, 0-49)
    5.242755, 5.224256, 5.198783, 5.167976, 5.133484, 5.096869, 5.059566, 
    5.022881, 4.987978, 4.955898, 4.927505, 4.903431, 4.883943, 4.868771, 
    4.856884, 30, 4.873823, 4.860311, 4.837456, 4.80504, 4.765738, 4.706779, 
    4.653216, 4.606438, 4.572193, 4.55386, 4.553253, 4.570012, 4.602548, 
    4.647337, 4.704798, 4.75439, 4.805976, 4.856723, 4.903411, 4.942552, 
    4.970578, 4.984347, 4.981996, 4.963964, 4.933707, 4.897477, 4.862895, 
    4.836847, 4.823806, 4.825346, 4.840734, 4.867923, 4.904401, 4.947665,
  // totalHeight(11,25, 0-49)
    5.240794, 5.22232, 5.196975, 5.166369, 5.132127, 5.095788, 5.058773, 
    5.022375, 4.987755, 4.955944, 4.927806, 4.903964, 4.884675, 4.869664, 
    4.8579, 30, 4.873703, 4.860322, 4.837665, 4.805562, 4.766716, 4.707583, 
    4.654046, 4.607269, 4.572984, 4.554605, 4.553962, 4.570693, 4.603181, 
    4.647916, 4.705504, 4.754699, 4.80592, 4.856369, 4.902862, 4.941946, 
    4.970081, 4.984127, 4.982181, 4.964595, 4.934705, 4.898656, 4.864019, 
    4.837709, 4.824278, 4.825392, 4.84038, 4.86723, 4.903439, 4.946502,
  // totalHeight(11,26, 0-49)
    5.236609, 5.218122, 5.192966, 5.162689, 5.128861, 5.092988, 5.056469, 
    5.020595, 4.98654, 4.955349, 4.927902, 4.904818, 4.886321, 4.872047, 
    4.860817, 30, 4.860604, 4.848742, 4.827468, 4.796851, 4.759639, 4.703284, 
    4.652233, 4.607754, 4.575406, 4.558476, 4.558778, 4.576014, 4.608685, 
    4.653347, 4.710508, 4.75958, 4.810529, 4.860532, 4.90638, 4.944607, 
    4.971689, 4.984544, 4.981393, 4.962756, 4.932151, 4.895843, 4.8614, 
    4.835618, 4.82288, 4.824695, 4.8403, 4.867644, 4.904226, 4.947563,
  // totalHeight(11,27, 0-49)
    5.230247, 5.211652, 5.186687, 5.156816, 5.12353, 5.088286, 5.052456, 
    5.017334, 4.984122, 4.953905, 4.927598, 4.90583, 4.888774, 4.875917, 
    4.8658, 30, 4.835612, 4.826562, 4.807929, 4.780112, 4.745865, 4.695104, 
    4.648843, 4.608716, 4.580005, 4.565769, 4.567803, 4.585944, 4.618935, 
    4.663445, 4.719617, 4.768734, 4.819421, 4.868762, 4.913473, 4.950031, 
    4.97492, 4.985185, 4.979329, 4.958301, 4.926076, 4.889226, 4.855335, 
    4.83092, 4.819949, 4.823555, 4.84074, 4.869361, 4.906916, 4.950954,
  // totalHeight(11,28, 0-49)
    5.221816, 5.202913, 5.178044, 5.148566, 5.115879, 5.081367, 5.046379, 
    5.012208, 4.980105, 4.951216, 4.926524, 4.906692, 4.891847, 4.881296, 
    4.873246, 30, 4.800921, 4.795757, 4.781104, 4.757642, 4.728002, 4.685359, 
    4.64586, 4.611671, 4.58779, 4.577054, 4.5813, 4.600579, 4.633968, 
    4.678254, 4.733004, 4.782204, 4.832494, 4.880813, 4.923745, 4.957682, 
    4.979128, 4.985353, 4.975339, 4.950729, 4.91621, 4.878789, 4.846007, 
    4.823902, 4.815784, 4.822229, 4.841906, 4.872549, 4.91166, 4.956846,
  // totalHeight(11,29, 0-49)
    5.211528, 5.191969, 5.166947, 5.13771, 5.105555, 5.071788, 5.037718, 
    5.004653, 4.97389, 4.946674, 4.924098, 4.906909, 4.895241, 4.888247, 
    4.883862, 30, 4.758096, 4.757624, 4.74851, 4.73148, 4.7087, 4.676564, 
    4.645609, 4.618504, 4.600053, 4.593021, 4.59944, 4.61967, 4.653188, 
    4.696864, 4.749561, 4.798358, 4.847646, 4.894192, 4.934445, 4.964732, 
    4.981649, 4.982831, 4.967932, 4.939481, 4.902971, 4.865784, 4.835213, 
    4.816581, 4.812366, 4.8225, 4.845302, 4.8784, 4.919327, 4.965767,
  // totalHeight(11,30, 0-49)
    5.203184, 5.185256, 5.161644, 5.13331, 5.101258, 5.066503, 5.030076, 
    4.993026, 4.956442, 4.921446, 4.889181, 4.860801, 4.837526, 4.82086, 
    4.81322, 4.793564, 4.759291, 4.783369, 4.786592, 4.771524, 4.744068, 
    4.707412, 4.671654, 4.641252, 4.621176, 4.613644, 4.620066, 4.640306, 
    4.673593, 4.716428, 4.766704, 4.814546, 4.862028, 4.905797, 4.942236, 
    4.967708, 4.97907, 4.974526, 4.954614, 4.922864, 4.885518, 4.850087, 
    4.823308, 4.809544, 4.810329, 4.82495, 4.851427, 4.887334, 4.930273, 
    4.978027,
  // totalHeight(11,31, 0-49)
    5.191897, 5.173043, 5.149139, 5.121112, 5.08991, 5.056485, 5.021814, 
    4.986914, 4.952852, 4.920757, 4.891789, 4.867128, 4.847923, 4.835331, 
    4.830701, 4.793941, 4.74672, 4.765321, 4.765812, 4.751783, 4.728415, 
    4.699248, 4.671027, 4.647578, 4.633379, 4.630328, 4.639804, 4.661777, 
    4.695667, 4.737928, 4.785717, 4.832349, 4.877781, 4.918511, 4.950845, 
    4.971227, 4.976875, 4.966708, 4.942261, 4.908067, 4.87096, 4.838338, 
    4.81617, 4.807773, 4.813767, 4.832868, 4.862859, 4.901292, 4.945847, 
    4.994394,
  // totalHeight(11,32, 0-49)
    5.182117, 5.162619, 5.138494, 5.110645, 5.079966, 5.047355, 5.013735, 
    4.980078, 4.947419, 4.916849, 4.889486, 4.866421, 4.848642, 4.836962, 
    4.832007, 4.788759, 4.739945, 4.751895, 4.749567, 4.736239, 4.716129, 
    4.69341, 4.671788, 4.654728, 4.646223, 4.647764, 4.660519, 4.684406, 
    4.718903, 4.760376, 4.805366, 4.850052, 4.892422, 4.928905, 4.955868, 
    4.970041, 4.969263, 4.95342, 4.925176, 4.889977, 4.854934, 4.826926, 
    4.810857, 4.808888, 4.820767, 4.844739, 4.87844, 4.919459, 4.965571, 
    5.014742,
  // totalHeight(11,33, 0-49)
    5.174572, 5.154589, 5.13018, 5.102248, 5.071674, 5.039321, 5.00607, 
    4.972849, 4.940649, 4.910503, 4.883449, 4.860447, 4.842265, 4.829318, 
    4.82152, 4.779136, 4.735283, 4.740807, 4.736142, 4.723701, 4.706699, 
    4.689884, 4.674292, 4.663169, 4.660039, 4.665985, 4.681876, 4.707491, 
    4.742249, 4.782453, 4.824167, 4.866026, 4.904251, 4.935326, 4.955851, 
    4.96308, 4.955732, 4.934846, 4.90422, 4.869962, 4.83904, 4.817427, 
    4.808751, 4.814018, 4.832221, 4.861261, 4.898711, 4.942233, 4.989711, 
    5.039204,
  // totalHeight(11,34, 0-49)
    5.170084, 5.149796, 5.125022, 5.096713, 5.065773, 5.033074, 4.999493, 
    4.965929, 4.933328, 4.902668, 4.874899, 4.850855, 4.831088, 4.815667, 
    4.803902, 4.766072, 4.730641, 4.730635, 4.724333, 4.713195, 4.699438, 
    4.68818, 4.678235, 4.672667, 4.674529, 4.684519, 4.703167, 4.730061, 
    4.764484, 4.802741, 4.840598, 4.878656, 4.91169, 4.936383, 4.949773, 
    4.949892, 4.936552, 4.912015, 4.881037, 4.849986, 4.825233, 4.811538, 
    4.81119, 4.824152, 4.848831, 4.882911, 4.923972, 4.969772, 5.0183, 
    5.067683,
  // totalHeight(11,35, 0-49)
    5.16936, 5.149054, 5.123928, 5.095007, 5.063273, 5.029659, 4.99507, 
    4.960418, 4.926631, 4.894642, 4.865333, 4.839435, 4.817364, 4.798974, 
    4.783234, 4.750862, 4.725138, 4.7207, 4.713482, 4.704073, 4.693744, 
    4.687737, 4.683125, 4.682759, 4.689171, 4.702719, 4.723572, 4.751113, 
    4.784435, 4.819942, 4.853301, 4.886603, 4.913572, 4.931258, 4.937376, 
    4.930943, 4.912982, 4.886868, 4.857957, 4.832395, 4.815557, 4.810833, 
    4.819266, 4.839981, 4.870982, 4.909855, 4.954227, 5.001952, 5.051094, 
    5.099827,
  // totalHeight(11,36, 0-49)
    5.172808, 5.152929, 5.127627, 5.098027, 5.065219, 5.030244, 4.994094, 
    4.95773, 4.922098, 4.888113, 4.856624, 4.828312, 4.803537, 4.782102, 
    4.762949, 4.735329, 4.718907, 4.711125, 4.703607, 4.696209, 4.689353, 
    4.688214, 4.688584, 4.693012, 4.703455, 4.719961, 4.742342, 4.769779, 
    4.801148, 4.833087, 4.861357, 4.889116, 4.909484, 4.920085, 4.919499, 
    4.907862, 4.887349, 4.862151, 4.837749, 4.819602, 4.811847, 4.816537, 
    4.833683, 4.861814, 4.898704, 4.941922, 4.989157, 5.038332, 5.08755, 
    5.134997,
  // totalHeight(11,37, 0-49)
    5.180398, 5.161556, 5.136457, 5.106329, 5.072402, 5.035862, 4.997823, 
    4.959341, 4.921418, 4.884993, 4.850913, 4.819863, 4.792229, 4.767898, 
    4.746009, 4.72179, 4.713002, 4.702868, 4.695462, 4.6901, 4.686528, 
    4.689706, 4.694558, 4.703251, 4.717091, 4.735848, 4.758998, 4.785535, 
    4.814129, 4.841794, 4.864573, 4.886342, 4.900098, 4.904203, 4.898227, 
    4.883398, 4.862806, 4.841026, 4.823173, 4.813704, 4.815465, 4.829372, 
    4.854675, 4.889541, 4.931647, 4.978592, 5.028115, 5.07816, 5.126826, 
    5.172269,
  // totalHeight(11,38, 0-49)
    5.191592, 5.174534, 5.150224, 5.119972, 5.085162, 5.047144, 5.007191, 
    4.966487, 4.926123, 4.887098, 4.850299, 4.816452, 4.786022, 4.759057, 
    4.735008, 4.712789, 4.70924, 4.697576, 4.690451, 4.686867, 4.686113, 
    4.692836, 4.701461, 4.713706, 4.730173, 4.750387, 4.773516, 4.798402, 
    4.82355, 4.846487, 4.86371, 4.879532, 4.88728, 4.886151, 4.876693, 
    4.861042, 4.842818, 4.826513, 4.816519, 4.816159, 4.827136, 4.849496, 
    4.882006, 4.922656, 4.969118, 5.019029, 5.070147, 5.120387, 5.167787, 
    5.210437,
  // totalHeight(11,39, 0-49)
    5.205347, 5.190912, 5.168145, 5.138416, 5.103247, 5.064161, 5.022605, 
    4.979915, 4.937297, 4.895839, 4.856494, 4.820059, 4.787104, 4.757856, 
    4.732081, 4.710703, 4.709868, 4.697269, 4.690359, 4.688056, 4.689408, 
    4.698699, 4.710176, 4.72507, 4.743271, 4.764093, 4.786444, 4.809061, 
    4.830353, 4.848471, 4.860497, 4.870972, 4.873897, 4.869296, 4.858545, 
    4.844366, 4.830497, 4.82097, 4.819266, 4.827655, 4.846931, 4.876558, 
    4.915043, 4.960332, 5.010135, 5.06212, 5.114024, 5.163682, 5.209023, 
    5.248034,
  // totalHeight(11,40, 0-49)
    5.220186, 5.209238, 5.188896, 5.160541, 5.125803, 5.086365, 5.043848, 
    4.999744, 4.955394, 4.911988, 4.870568, 4.832009, 4.796983, 4.765884, 
    4.73874, 4.717393, 4.717087, 4.703911, 4.69698, 4.695314, 4.697904, 
    4.708665, 4.721914, 4.738419, 4.75739, 4.777978, 4.798889, 4.81882, 
    4.836173, 4.849782, 4.857394, 4.863602, 4.863284, 4.857172, 4.847208, 
    4.836345, 4.828079, 4.825771, 4.831997, 4.848148, 4.874382, 4.90982, 
    4.95287, 5.001508, 5.053501, 5.106535, 5.158285, 5.206468, 5.248866, 
    5.283354,
  // totalHeight(11,41, 0-49)
    5.23431, 5.227661, 5.210699, 5.184736, 5.151451, 5.112651, 5.070111, 
    5.025473, 4.980214, 4.935633, 4.892861, 4.852852, 4.816367, 4.783926, 
    4.755749, 4.733974, 4.732622, 4.719017, 4.711739, 4.710033, 4.712957, 
    4.724083, 4.737983, 4.755019, 4.773808, 4.793388, 4.812348, 4.829412, 
    4.84305, 4.852812, 4.85709, 4.860407, 4.858553, 4.852761, 4.845245, 
    4.838876, 4.836684, 4.841298, 4.854504, 4.87704, 4.908657, 4.948308, 
    4.994401, 5.044983, 5.097881, 5.150779, 5.201279, 5.246957, 5.285442, 
    5.314502,
  // totalHeight(11,42, 0-49)
    5.245757, 5.244094, 5.231469, 5.209024, 5.178406, 5.141475, 5.100114, 
    5.056091, 5.011003, 4.966255, 4.923054, 4.882427, 4.845201, 4.811985, 
    4.783129, 4.76075, 4.75743, 4.7434, 4.735441, 4.733069, 4.735492, 
    4.745985, 4.759491, 4.776057, 4.793811, 4.811748, 4.828418, 4.84264, 
    4.853035, 4.859815, 4.861965, 4.863824, 4.861996, 4.857988, 4.854019, 
    4.852657, 4.856369, 4.867102, 4.886012, 4.913383, 4.948726, 4.99094, 
    5.038484, 5.089493, 5.141856, 5.193256, 5.241224, 5.283213, 5.316723, 
    5.33947,
  // totalHeight(11,43, 0-49)
    5.252583, 5.256382, 5.248981, 5.231237, 5.20464, 5.171007, 5.132254, 
    5.090226, 5.046606, 5.002879, 4.96032, 4.92001, 4.882821, 4.849424, 
    4.820261, 4.797302, 4.791629, 4.777101, 4.768164, 4.764614, 4.765842, 
    4.774894, 4.787142, 4.802403, 4.818435, 4.834261, 4.848473, 4.860041, 
    4.867776, 4.872492, 4.873652, 4.875337, 4.87478, 4.873552, 4.873688, 
    4.877326, 4.886364, 4.902164, 4.925396, 4.95604, 4.993475, 5.036603, 
    5.083958, 5.133768, 5.18399, 5.232327, 5.276277, 5.313229, 5.340635, 
    5.356261,
  // totalHeight(11,44, 0-49)
    5.253074, 5.262515, 5.261069, 5.249179, 5.228035, 5.199276, 5.164745, 
    5.12628, 5.085594, 5.044218, 5.003467, 4.964456, 4.928098, 4.895112, 
    4.866016, 4.842618, 4.834599, 4.819472, 4.809327, 4.804217, 4.803734, 
    4.810767, 4.821117, 4.834463, 4.848287, 4.861711, 4.873432, 4.882618, 
    4.888287, 4.891765, 4.892875, 4.89539, 4.896967, 4.89908, 4.90345, 
    4.911751, 4.925344, 4.945101, 4.971322, 5.003768, 5.041742, 5.084168, 
    5.129661, 5.176544, 5.222858, 5.266371, 5.304625, 5.335056, 5.355216, 
    5.363077,
  // totalHeight(11,45, 0-49)
    5.245976, 5.260865, 5.26584, 5.260825, 5.246549, 5.224311, 5.19573, 
    5.162527, 5.126361, 5.08875, 5.05102, 5.014307, 4.97956, 4.947553, 
    4.918889, 4.895254, 4.885153, 4.869344, 4.85784, 4.850928, 4.848397, 
    4.853063, 4.861111, 4.872155, 4.883486, 4.894375, 4.903677, 4.910774, 
    4.914892, 4.917789, 4.919525, 4.923557, 4.927764, 4.933413, 4.941857, 
    4.954303, 4.971632, 4.994293, 5.02229, 5.055206, 5.092278, 5.13245, 
    5.174401, 5.216556, 5.257073, 5.293852, 5.324604, 5.34698, 5.358833, 
    5.358551,
  // totalHeight(11,46, 0-49)
    5.230698, 5.250425, 5.261923, 5.264531, 5.258378, 5.244246, 5.223355, 
    5.197155, 5.167138, 5.134735, 5.101245, 5.067813, 5.035434, 5.004955, 
    4.977088, 4.953472, 4.941727, 4.925207, 4.912287, 4.903466, 4.898721, 
    4.900876, 4.90643, 4.914997, 4.923724, 4.932077, 4.939089, 4.944373, 
    4.94734, 4.950113, 4.952881, 4.958815, 4.965834, 4.974938, 4.987098, 
    5.003079, 5.023328, 5.047932, 5.076622, 5.108816, 5.143669, 5.180115, 
    5.216885, 5.252507, 5.285301, 5.313405, 5.334856, 5.347742, 5.35046, 
    5.342037,
  // totalHeight(11,47, 0-49)
    5.207477, 5.23103, 5.248695, 5.259253, 5.262141, 5.257459, 5.24584, 
    5.228285, 5.205985, 5.18019, 5.152124, 5.122934, 5.093671, 5.065282, 
    5.03861, 5.015327, 5.00253, 4.985361, 4.971079, 4.96038, 4.953408, 
    4.953086, 4.956131, 4.962209, 4.968366, 4.974279, 4.979176, 4.982888, 
    4.984988, 4.987902, 4.991867, 4.999817, 5.009564, 5.021826, 5.037194, 
    5.056029, 5.07839, 5.104032, 5.132427, 5.162814, 5.194239, 5.225595, 
    5.255641, 5.283024, 5.306286, 5.323929, 5.334507, 5.336784, 5.329955, 
    5.313877,
  // totalHeight(11,48, 0-49)
    5.177426, 5.203481, 5.226476, 5.244749, 5.257052, 5.262691, 5.261548, 
    5.253999, 5.240782, 5.222868, 5.201346, 5.177341, 5.151967, 5.126286, 
    5.101289, 5.078762, 5.06565, 5.04801, 5.03255, 5.020142, 5.011084, 
    5.008462, 5.009127, 5.012832, 5.016562, 5.020209, 5.023188, 5.025537, 
    5.026949, 5.030105, 5.035226, 5.045074, 5.057245, 5.072175, 5.090107, 
    5.111032, 5.134658, 5.16043, 5.187572, 5.215123, 5.242, 5.267024, 
    5.288981, 5.30666, 5.318905, 5.324718, 5.323361, 5.314494, 5.298303, 
    5.275572,
  // totalHeight(11,49, 0-49)
    5.130487, 5.157133, 5.184359, 5.21029, 5.233043, 5.250996, 5.26301, 
    5.268517, 5.267499, 5.260395, 5.247995, 5.231311, 5.211483, 5.189702, 
    5.167173, 5.146682, 5.140685, 5.122538, 5.104847, 5.089356, 5.0769, 
    5.074059, 5.074942, 5.079597, 5.082418, 5.084044, 5.083921, 5.082497, 
    5.079126, 5.079224, 5.082874, 5.095003, 5.110043, 5.128022, 5.148745, 
    5.171737, 5.196276, 5.221437, 5.24613, 5.269165, 5.289305, 5.305318, 
    5.316079, 5.32065, 5.318389, 5.309089, 5.293078, 5.271255, 5.245065, 
    5.216325,
  // totalHeight(12,0, 0-49)
    5.283156, 5.303393, 5.315825, 5.319623, 5.31465, 5.301387, 5.280786, 
    5.254111, 5.222781, 5.188264, 5.151982, 5.115261, 5.079288, 5.045088, 
    5.013504, 4.985375, 4.962522, 4.942296, 4.926528, 4.915215, 4.908121, 
    4.905272, 4.90585, 4.909438, 4.915286, 4.922814, 4.93137, 4.940413, 
    4.949502, 4.958674, 4.967987, 4.978175, 4.989471, 5.002637, 5.018452, 
    5.037585, 5.060488, 5.087313, 5.117883, 5.15169, 5.18792, 5.225489, 
    5.263074, 5.299156, 5.332043, 5.359944, 5.381062, 5.393738, 5.396669, 
    5.389134,
  // totalHeight(12,1, 0-49)
    5.289672, 5.306209, 5.313846, 5.31217, 5.301459, 5.28255, 5.256652, 
    5.225194, 5.189679, 5.15159, 5.112332, 5.073187, 5.035285, 4.999592, 
    4.966884, 4.938138, 4.916506, 4.896032, 4.880301, 4.86932, 4.862805, 
    4.861174, 4.863127, 4.868292, 4.875661, 4.884639, 4.894459, 4.904496, 
    4.91414, 4.923573, 4.932739, 4.942745, 4.953437, 4.965678, 4.980408, 
    4.998491, 5.020582, 5.047031, 5.077825, 5.112586, 5.150586, 5.19079, 
    5.231888, 5.272332, 5.310356, 5.344034, 5.371366, 5.390417, 5.399523, 
    5.397548,
  // totalHeight(12,2, 0-49)
    5.289351, 5.301156, 5.303457, 5.296273, 5.280246, 5.256473, 5.226311, 
    5.191248, 5.152781, 5.112347, 5.071281, 5.030792, 4.991937, 4.955608, 
    4.922512, 4.893762, 4.873818, 4.853418, 4.837952, 4.827422, 4.821506, 
    4.821013, 4.824201, 4.830774, 4.839534, 4.849892, 4.860994, 4.872135, 
    4.882534, 4.892459, 4.901697, 4.911676, 4.921791, 4.932947, 4.946202, 
    4.962606, 4.983036, 5.008065, 5.037891, 5.072294, 5.110664, 5.152039, 
    5.195147, 5.238437, 5.280128, 5.318251, 5.350725, 5.375486, 5.390674, 
    5.394858,
  // totalHeight(12,3, 0-49)
    5.282612, 5.289087, 5.285932, 5.273549, 5.252862, 5.225129, 5.191766, 
    5.154241, 5.113979, 5.072326, 5.030522, 4.989674, 4.950751, 4.914566, 
    4.881744, 4.85353, 4.835714, 4.815639, 4.800602, 4.790585, 4.785224, 
    4.785729, 4.789946, 4.797691, 4.807655, 4.819279, 4.831649, 4.843991, 
    4.855368, 4.866057, 4.875648, 4.885847, 4.895519, 4.905539, 4.917031, 
    4.931207, 4.949178, 4.971781, 4.999463, 5.032219, 5.069589, 5.110712, 
    5.154368, 5.199042, 5.24297, 5.2842, 5.320669, 5.350304, 5.37118, 5.381702,
  // totalHeight(12,4, 0-49)
    5.270433, 5.271401, 5.263016, 5.245987, 5.221428, 5.190666, 5.15511, 
    5.116154, 5.07512, 5.033241, 4.991632, 4.951296, 4.9131, 4.877757, 
    4.845793, 4.818586, 4.803279, 4.783717, 4.769216, 4.759707, 4.754789, 
    4.756079, 4.761035, 4.769634, 4.780541, 4.793252, 4.806829, 4.820447, 
    4.833023, 4.844786, 4.855074, 4.865842, 4.87534, 4.884321, 4.893908, 
    4.905432, 4.92024, 4.93947, 4.963875, 4.993721, 5.02876, 5.068261, 
    5.111091, 5.155785, 5.200624, 5.243716, 5.283067, 5.316677, 5.342657, 
    5.359342,
  // totalHeight(12,5, 0-49)
    5.254186, 5.249829, 5.236703, 5.215734, 5.188132, 5.155237, 5.118395, 
    5.078903, 5.037965, 4.996687, 4.956069, 4.916993, 4.880211, 4.84632, 
    4.815726, 4.789899, 4.777379, 4.758461, 4.744543, 4.735467, 4.730793, 
    4.732566, 4.737878, 4.74691, 4.758401, 4.771935, 4.786589, 4.801508, 
    4.815494, 4.828657, 4.840042, 4.851838, 4.861586, 4.869823, 4.877574, 
    4.886226, 4.897335, 4.912361, 4.932431, 4.958163, 4.989584, 5.026161, 
    5.066878, 5.110339, 5.154894, 5.19872, 5.239929, 5.276628, 5.30701, 
    5.329417,
  // totalHeight(12,6, 0-49)
    5.235466, 5.226234, 5.209022, 5.184886, 5.155065, 5.120851, 5.083508, 
    5.044224, 5.004089, 4.964089, 4.925107, 4.88791, 4.853123, 4.821205, 
    4.792401, 4.768209, 4.758565, 4.740386, 4.727033, 4.718237, 4.713521, 
    4.715374, 4.720548, 4.729478, 4.741088, 4.755076, 4.770578, 4.786751, 
    4.802309, 4.817187, 4.830103, 4.84348, 4.854072, 4.862099, 4.868368, 
    4.874223, 4.881364, 4.891574, 4.906406, 4.926915, 4.953505, 4.985915, 
    5.023302, 5.064378, 5.107562, 5.151116, 5.193247, 5.232182, 5.266211, 
    5.293715,
  // totalHeight(12,7, 0-49)
    5.215919, 5.202434, 5.181869, 5.155337, 5.124051, 5.089231, 5.052039, 
    5.013558, 4.974773, 4.936571, 4.899731, 4.864904, 4.832586, 4.803066, 
    4.776391, 4.753929, 4.746964, 4.729606, 4.716753, 4.708011, 4.702882, 
    4.704314, 4.708754, 4.716944, 4.728096, 4.742053, 4.758061, 4.775326, 
    4.792534, 4.809388, 4.824256, 4.839813, 4.851985, 4.860579, 4.86606, 
    4.869582, 4.872879, 4.878002, 4.88695, 4.901301, 4.921952, 4.949025, 
    4.981931, 5.019534, 5.060344, 5.102702, 5.144898, 5.185256, 5.222154, 
    5.254018,
  // totalHeight(12,8, 0-49)
    5.197084, 5.180053, 5.15687, 5.128651, 5.096552, 5.0617, 5.02516, 
    4.987918, 4.950877, 4.914841, 4.880503, 4.848413, 4.818925, 4.792144, 
    4.76786, 4.747036, 4.742175, 4.725766, 4.713326, 4.70436, 4.698389, 
    4.698829, 4.701871, 4.708604, 4.71863, 4.731961, 4.748012, 4.766073, 
    4.784878, 4.803852, 4.82102, 4.839316, 4.853869, 4.863999, 4.869711, 
    4.871802, 4.871869, 4.872107, 4.874922, 4.882471, 4.896258, 4.916928, 
    4.944264, 4.977354, 5.014838, 5.055129, 5.096582, 5.137584, 5.17657, 
    5.212003,
  // totalHeight(12,9, 0-49)
    5.180264, 5.160401, 5.13527, 5.105958, 5.07355, 5.03908, 5.003524, 
    4.967793, 4.932725, 4.899067, 4.86745, 4.838332, 4.811933, 4.788154, 
    4.766489, 4.747004, 4.743248, 4.728023, 4.715933, 4.706465, 4.699218, 
    4.698076, 4.699035, 4.70357, 4.711748, 4.723778, 4.739289, 4.757714, 
    4.777895, 4.798965, 4.818629, 4.840088, 4.857762, 4.870472, 4.877666, 
    4.879622, 4.877593, 4.873718, 4.870685, 4.871213, 4.877508, 4.890886, 
    4.911653, 4.939244, 4.972483, 5.00987, 5.049802, 5.090693, 5.131, 5.169196,
  // totalHeight(12,10, 0-49)
    5.166411, 5.144372, 5.117849, 5.087887, 5.0555, 5.021643, 4.987225, 
    4.9531, 4.920068, 4.888845, 4.86002, 4.833982, 4.810833, 4.790262, 
    4.771456, 4.752806, 4.748785, 4.735146, 4.723433, 4.713244, 4.704352, 
    4.701074, 4.699321, 4.700947, 4.706553, 4.716559, 4.730864, 4.749084, 
    4.770245, 4.79319, 4.815342, 4.840149, 4.861498, 4.877731, 4.887707, 
    4.891069, 4.888515, 4.881875, 4.873897, 4.867746, 4.866354, 4.871841, 
    4.885215, 4.906405, 4.934523, 4.968196, 5.005853, 5.045899, 5.086775, 
    5.126939,
  // totalHeight(12,11, 0-49)
    5.156057, 5.132392, 5.104886, 5.074547, 5.042329, 5.009131, 4.975822, 
    4.943227, 4.912133, 4.883249, 4.85715, 4.83418, 4.814344, 4.797164, 
    4.781535, 4.763055, 4.757185, 4.745727, 4.734569, 4.723561, 4.712773, 
    4.706907, 4.701915, 4.700012, 4.70236, 4.709619, 4.721997, 4.739341, 
    4.760933, 4.785336, 4.809756, 4.837816, 4.863089, 4.883525, 4.89742, 
    4.90373, 4.902445, 4.894832, 4.883407, 4.871558, 4.862848, 4.860272, 
    4.865705, 4.879758, 4.901966, 4.931159, 4.965813, 5.004309, 5.045033, 
    5.086396,
  // totalHeight(12,12, 0-49)
    5.149285, 5.12441, 5.096178, 5.065566, 5.033495, 5.000843, 4.968459, 
    4.937173, 4.907782, 4.881011, 4.857444, 4.837414, 4.820879, 4.807252, 
    4.795251, 4.776213, 4.766981, 4.758471, 4.748212, 4.73646, 4.723689, 
    4.714914, 4.706287, 4.700346, 4.698822, 4.702633, 4.712355, 4.728104, 
    4.74946, 4.774756, 4.801041, 4.831972, 4.861088, 4.886032, 4.904624, 
    4.915174, 4.916892, 4.910286, 4.897347, 4.881368, 4.866335, 4.856068, 
    4.853416, 4.859857, 4.875521, 4.899554, 4.930533, 4.966812, 5.006703, 
    5.048541,
  // totalHeight(12,13, 0-49)
    5.145769, 5.119963, 5.09112, 5.060205, 5.028135, 4.995795, 4.964047, 
    4.933748, 4.905724, 4.880737, 4.859405, 4.842088, 4.828754, 4.818828, 
    4.811018, 4.790828, 4.777141, 4.772433, 4.763588, 4.751352, 4.736684, 
    4.724803, 4.712266, 4.701881, 4.695943, 4.695662, 4.70202, 4.715442, 
    4.735847, 4.761384, 4.789021, 4.822229, 4.854795, 4.884152, 4.90777, 
    4.923401, 4.929517, 4.925776, 4.913407, 4.895278, 4.875484, 4.858485, 
    4.848105, 4.846823, 4.855548, 4.87389, 4.900612, 4.934071, 4.9725, 5.01414,
  // totalHeight(12,14, 0-49)
    5.144871, 5.118295, 5.088853, 5.057521, 5.02524, 4.992924, 4.961475, 
    4.931789, 4.904742, 4.881144, 4.861664, 4.846729, 4.836396, 4.830227, 
    4.827164, 4.805708, 4.787249, 4.787188, 4.780379, 4.768078, 4.751752, 
    4.736667, 4.720029, 4.704872, 4.694035, 4.689069, 4.691406, 4.701812, 
    4.720558, 4.745669, 4.774117, 4.808887, 4.844282, 4.877623, 4.906136, 
    4.927167, 4.938556, 4.939137, 4.929252, 4.911079, 4.888462, 4.866208, 
    4.848984, 4.840306, 4.842016, 4.854346, 4.876366, 4.906497, 4.942909, 
    4.983748,
  // totalHeight(12,15, 0-49)
    5.145796, 5.118527, 5.088447, 5.056561, 5.023852, 4.991281, 4.959796, 
    4.930346, 4.903856, 4.881192, 4.863095, 4.850088, 4.842387, 4.839818, 
    4.841783, 4.819959, 4.797536, 4.802824, 4.798692, 4.786848, 4.769209, 
    4.750873, 4.72998, 4.709755, 4.693579, 4.683396, 4.681126, 4.687901, 
    4.70434, 4.728413, 4.75718, 4.792764, 4.83025, 4.866904, 4.899821, 
    4.926082, 4.943048, 4.948842, 4.942933, 4.92663, 4.903234, 4.877543, 
    4.854808, 4.839509, 4.834488, 4.840753, 4.857808, 4.884229, 4.918171, 
    4.957691,
  // totalHeight(12,16, 0-49)
    5.14775, 5.119838, 5.089086, 5.056542, 5.023234, 4.99017, 4.958349, 
    4.928762, 4.902383, 4.88013, 4.862822, 4.851107, 4.845402, 4.84588, 
    4.852536, 4.832886, 4.808788, 4.819836, 4.818934, 4.808081, 4.789505, 
    4.767872, 4.742556, 4.716972, 4.695046, 4.67918, 4.671813, 4.674458, 
    4.688052, 4.710579, 4.739286, 4.774993, 4.813807, 4.852983, 4.889573, 
    4.920512, 4.942851, 4.954165, 4.953143, 4.940207, 4.917892, 4.890668, 
    4.864047, 4.843275, 4.83217, 4.832603, 4.844646, 4.867138, 4.898277, 
    4.936063,
  // totalHeight(12,17, 0-49)
    5.150093, 5.121617, 5.090219, 5.056981, 5.022968, 4.989228, 4.956792, 
    4.926682, 4.899899, 4.877413, 4.860113, 4.84878, 4.844049, 4.846456, 
    4.856596, 4.843801, 4.822259, 4.838977, 4.841652, 4.832212, 4.813004, 
    4.787975, 4.758004, 4.726743, 4.698685, 4.676764, 4.663949, 4.662121, 
    4.672501, 4.693131, 4.72155, 4.756793, 4.796225, 4.837117, 4.876529, 
    4.911358, 4.938486, 4.955118, 4.959318, 4.950685, 4.930918, 4.903908, 
    4.875101, 4.850234, 4.833983, 4.829096, 4.836311, 4.854834, 4.882985, 
    4.918743,
  // totalHeight(12,18, 0-49)
    5.152446, 5.123583, 5.091654, 5.057766, 5.023003, 4.988423, 4.955067, 
    4.923962, 4.896122, 4.872548, 4.854192, 4.841951, 4.836679, 4.839291, 
    4.851016, 4.851833, 4.839601, 4.861182, 4.867465, 4.859635, 4.839867, 
    4.81117, 4.776155, 4.738822, 4.704293, 4.676091, 4.657684, 4.651282, 
    4.65831, 4.676892, 4.704975, 4.739322, 4.778765, 4.820615, 4.861983, 
    4.8998, 4.930897, 4.952261, 4.961515, 4.957573, 4.941316, 4.915917, 
    4.886491, 4.85898, 4.838706, 4.829237, 4.832021, 4.846715, 4.871841, 
    4.905409,
  // totalHeight(12,19, 0-49)
    5.154763, 5.125841, 5.093623, 5.059199, 5.023643, 4.987998, 4.95329, 
    4.920535, 4.890742, 4.864912, 4.844035, 4.829114, 4.82127, 4.821993, 
    4.833523, 4.855882, 4.862566, 4.887558, 4.897141, 4.890828, 4.870145, 
    4.837114, 4.796288, 4.752288, 4.710979, 4.67649, 4.652683, 4.64197, 
    4.645842, 4.66249, 4.690382, 4.723572, 4.762553, 4.804698, 4.847201, 
    4.887078, 4.921197, 4.946469, 4.960234, 4.960886, 4.948586, 4.925761, 
    4.897009, 4.868209, 4.845094, 4.831927, 4.83085, 4.842024, 4.864239, 
    4.895589,
  // totalHeight(12,20, 0-49)
    5.154693, 5.1242, 5.09093, 5.056166, 5.021146, 4.987069, 4.955105, 
    4.926386, 4.901967, 4.88274, 4.869288, 4.861674, 4.859224, 4.860402, 
    4.862944, 30, 4.887241, 4.889175, 4.884861, 4.87331, 4.854144, 4.824542, 
    4.78899, 4.749675, 4.711314, 4.677715, 4.653001, 4.640221, 4.641569, 
    4.655976, 4.682993, 4.71405, 4.751464, 4.792706, 4.835068, 4.875674, 
    4.911485, 4.939419, 4.956679, 4.961297, 4.952844, 4.933036, 4.905849, 
    4.876883, 4.852042, 4.836103, 4.831837, 4.839926, 4.859478, 4.888717,
  // totalHeight(12,21, 0-49)
    5.155864, 5.125593, 5.092457, 5.057732, 5.02263, 4.988307, 4.955864, 
    4.926349, 4.90071, 4.879722, 4.863865, 4.853156, 4.846985, 4.843976, 
    4.841977, 30, 4.928431, 4.928067, 4.921334, 4.906662, 4.883474, 4.84574, 
    4.802858, 4.756638, 4.712227, 4.67375, 4.64543, 4.630235, 4.630127, 
    4.64397, 4.671875, 4.702372, 4.7396, 4.78107, 4.82414, 4.866025, 
    4.903787, 4.934397, 4.954999, 4.963388, 4.958678, 4.941965, 4.916625, 
    4.887901, 4.861739, 4.843331, 4.83602, 4.841007, 4.857741, 4.884601,
  // totalHeight(12,22, 0-49)
    5.156168, 5.126009, 5.092949, 5.05825, 5.023098, 4.988604, 4.955816, 
    4.925714, 4.899168, 4.876884, 4.859283, 4.846379, 4.837635, 4.831826, 
    4.826962, 30, 4.95737, 4.955109, 4.947015, 4.931, 4.906226, 4.863213, 
    4.81588, 4.765259, 4.716686, 4.674536, 4.643195, 4.62569, 4.623909, 
    4.63674, 4.664946, 4.694184, 4.7305, 4.771442, 4.814431, 4.856776, 
    4.895633, 4.928053, 4.951179, 4.962662, 4.96128, 4.947614, 4.924472, 
    4.896675, 4.870069, 4.850082, 4.840516, 4.843034, 4.857418, 4.882221,
  // totalHeight(12,23, 0-49)
    5.155862, 5.125789, 5.092804, 5.058161, 5.023019, 4.988459, 4.955489, 
    4.925042, 4.897942, 4.874845, 4.856148, 4.84187, 4.831531, 4.824033, 
    4.817537, 30, 4.976377, 4.972693, 4.963794, 4.947212, 4.921901, 4.875348, 
    4.825215, 4.771749, 4.720391, 4.675718, 4.642266, 4.623123, 4.620123, 
    4.632184, 4.660638, 4.688662, 4.724012, 4.764284, 4.806946, 4.849384, 
    4.888843, 4.92245, 4.947373, 4.961187, 4.962439, 4.951327, 4.930201, 
    4.903494, 4.876895, 4.855958, 4.8448, 4.845447, 4.857971, 4.881085,
  // totalHeight(12,24, 0-49)
    5.155117, 5.125144, 5.092268, 5.057733, 5.022682, 4.988179, 4.955212, 
    4.924688, 4.897405, 4.873996, 4.85484, 4.839958, 4.828905, 4.820646, 
    4.81344, 30, 4.985891, 4.981441, 4.972165, 4.95543, 4.930089, 4.881607, 
    4.830071, 4.775189, 4.722447, 4.676545, 4.642097, 4.622215, 4.618693, 
    4.630451, 4.65923, 4.686486, 4.721179, 4.760937, 4.803261, 4.84558, 
    4.885197, 4.919293, 4.945075, 4.960088, 4.962771, 4.953119, 4.93321, 
    4.907235, 4.880754, 4.85936, 4.84734, 4.846935, 4.858387, 4.880515,
  // totalHeight(12,25, 0-49)
    5.154003, 5.124162, 5.091442, 5.057076, 5.022206, 4.987893, 4.955125, 
    4.924804, 4.897723, 4.874507, 4.855525, 4.840787, 4.829843, 4.821658, 
    4.814504, 30, 4.985445, 4.981015, 4.971813, 4.955236, 4.930161, 4.881445, 
    4.829905, 4.775073, 4.722418, 4.676649, 4.642362, 4.622644, 4.61925, 
    4.63111, 4.66012, 4.687131, 4.721565, 4.761066, 4.803155, 4.84528, 
    4.884767, 4.918823, 4.94467, 4.959867, 4.962834, 4.953512, 4.933909, 
    4.908139, 4.88171, 4.860214, 4.847972, 4.847279, 4.858426, 4.880264,
  // totalHeight(12,26, 0-49)
    5.152479, 5.122794, 5.090271, 5.056139, 5.021544, 4.98756, 4.955191, 
    4.925356, 4.898864, 4.876347, 4.858164, 4.84431, 4.834285, 4.826993, 
    4.820641, 30, 4.975043, 4.971416, 4.962752, 4.946657, 4.92212, 4.874942, 
    4.824836, 4.771557, 4.72049, 4.676219, 4.64323, 4.624537, 4.621883, 
    4.634203, 4.663285, 4.690606, 4.725205, 4.764738, 4.80672, 4.848597, 
    4.887678, 4.921165, 4.946287, 4.960632, 4.962692, 4.952519, 4.932245, 
    4.906088, 4.879598, 4.858325, 4.846496, 4.846295, 4.857932, 4.880213,
  // totalHeight(12,27, 0-49)
    5.150397, 5.120863, 5.088561, 5.054716, 5.020484, 4.986965, 4.955193, 
    4.926123, 4.900596, 4.879271, 4.862515, 4.85029, 4.842027, 4.836516, 
    4.831839, 30, 4.955084, 4.952917, 4.945256, 4.930057, 4.906505, 4.862667, 
    4.815493, 4.76527, 4.717227, 4.67572, 4.645051, 4.628139, 4.626747, 
    4.639816, 4.668792, 4.696878, 4.731983, 4.77176, 4.813708, 4.855239, 
    4.893616, 4.925999, 4.949613, 4.96211, 4.962144, 4.950032, 4.928223, 
    4.901196, 4.874612, 4.853933, 4.843158, 4.844211, 4.857095, 4.880501,
  // totalHeight(12,28, 0-49)
    5.147523, 5.118073, 5.085974, 5.052443, 5.018648, 4.985715, 4.954721, 
    4.926675, 4.902474, 4.882824, 4.868122, 4.858309, 4.85273, 4.850033, 
    4.848179, 30, 4.926608, 4.926298, 4.920071, 4.906347, 4.884541, 4.845834, 
    4.803155, 4.757463, 4.713751, 4.676086, 4.648576, 4.634062, 4.63437, 
    4.648452, 4.677229, 4.706404, 4.742229, 4.782332, 4.82418, 4.865112, 
    4.902321, 4.932904, 4.95409, 4.963649, 4.960521, 4.945456, 4.921401, 
    4.893226, 4.866715, 4.847156, 4.838172, 4.84128, 4.85618, 4.881395,
  // totalHeight(12,29, 0-49)
    5.143562, 5.11403, 5.082041, 5.048799, 5.015478, 4.983227, 4.953168, 
    4.926374, 4.903827, 4.886317, 4.874309, 4.867758, 4.86593, 4.867328, 
    4.869853, 30, 4.889934, 4.891613, 4.88732, 4.875996, 4.857266, 4.825638, 
    4.789297, 4.749714, 4.711526, 4.678509, 4.654641, 4.642774, 4.644877, 
    4.659924, 4.688231, 4.718379, 4.754757, 4.794957, 4.836395, 4.876332, 
    4.911868, 4.940042, 4.958111, 4.964036, 4.957141, 4.938742, 4.912372, 
    4.883308, 4.857393, 4.839608, 4.833077, 4.838827, 4.856208, 4.883573,
  // totalHeight(12,30, 0-49)
    5.140514, 5.112536, 5.081708, 5.049011, 5.015432, 4.981946, 4.949521, 
    4.919111, 4.891653, 4.868042, 4.849143, 4.835805, 4.82899, 4.830027, 
    4.841019, 4.861464, 4.864655, 4.888956, 4.899061, 4.894265, 4.875897, 
    4.843383, 4.804152, 4.761779, 4.721758, 4.68805, 4.664435, 4.653369, 
    4.656442, 4.672151, 4.699848, 4.730855, 4.767568, 4.807538, 4.848127, 
    4.886528, 4.91977, 4.944874, 4.959198, 4.960996, 4.950107, 4.928501, 
    4.900321, 4.871173, 4.846792, 4.831698, 4.828403, 4.837403, 4.857709, 
    4.887527,
  // totalHeight(12,31, 0-49)
    5.134956, 5.106979, 5.076535, 5.044599, 5.012144, 4.980138, 4.949538, 
    4.921287, 4.896299, 4.875444, 4.859525, 4.84926, 4.845331, 4.848502, 
    4.859925, 4.859009, 4.845135, 4.865917, 4.872577, 4.866015, 4.848228, 
    4.820029, 4.786397, 4.750472, 4.717049, 4.68944, 4.671017, 4.664021, 
    4.67, 4.687367, 4.714871, 4.746837, 4.783939, 4.823677, 4.863338, 
    4.900009, 4.93064, 4.952261, 4.962398, 4.959703, 4.944641, 4.919906, 
    4.890231, 4.861438, 4.83902, 4.826921, 4.826994, 4.839206, 4.862264, 
    4.894248,
  // totalHeight(12,32, 0-49)
    5.129212, 5.101433, 5.071481, 5.040294, 5.008811, 4.97796, 4.948673, 
    4.921868, 4.898431, 4.87919, 4.864866, 4.856045, 4.853179, 4.856658, 
    4.867016, 4.852871, 4.831022, 4.847097, 4.850173, 4.841893, 4.824452, 
    4.79999, 4.771226, 4.741108, 4.713883, 4.692271, 4.679163, 4.676469, 
    4.685562, 4.704714, 4.732142, 4.764843, 4.801892, 4.840762, 4.878683, 
    4.912685, 4.939712, 4.956912, 4.96214, 4.954616, 4.93555, 4.908378, 
    4.878297, 4.851113, 4.831837, 4.823677, 4.827783, 4.84363, 4.869668, 
    4.90391,
  // totalHeight(12,33, 0-49)
    5.12343, 5.095872, 5.066374, 5.035829, 5.005118, 4.975122, 4.946723, 
    4.920801, 4.898202, 4.879708, 4.865957, 4.8574, 4.854257, 4.856545, 
    4.864198, 4.843874, 4.820434, 4.831309, 4.831038, 4.821383, 4.804472, 
    4.783561, 4.75934, 4.73466, 4.713286, 4.697415, 4.689446, 4.690929, 
    4.70299, 4.723768, 4.751048, 4.784074, 4.82048, 4.857722, 4.89301, 
    4.92337, 4.945841, 4.957834, 4.957703, 4.945395, 4.922944, 4.894461, 
    4.865391, 4.841245, 4.82632, 4.822978, 4.831672, 4.851446, 4.880571, 
    4.91704,
  // totalHeight(12,34, 0-49)
    5.118104, 5.090694, 5.0615, 5.031375, 5.001149, 4.971647, 4.943697, 
    4.918133, 4.895763, 4.877318, 4.863366, 4.854235, 4.849931, 4.850104, 
    4.854072, 4.83257, 4.811661, 4.817543, 4.81448, 4.804032, 4.788081, 
    4.770701, 4.75087, 4.731368, 4.715502, 4.705021, 4.701844, 4.707161, 
    4.721816, 4.74386, 4.770767, 4.803555, 4.838606, 4.873378, 4.905098, 
    4.930877, 4.947974, 4.954234, 4.948682, 4.932118, 4.907397, 4.87913, 
    4.852721, 4.83309, 4.823634, 4.825835, 4.8395, 4.863335, 4.895511, 
    4.934046,
  // totalHeight(12,35, 0-49)
    5.113986, 5.086621, 5.057515, 5.027502, 4.997377, 4.967923, 4.939924, 
    4.914174, 4.891447, 4.872436, 4.85766, 4.847354, 4.841359, 4.839027, 
    4.839162, 4.81933, 4.803371, 4.80494, 4.799863, 4.789345, 4.774886, 
    4.761084, 4.745565, 4.731028, 4.720322, 4.714813, 4.715966, 4.724633, 
    4.74135, 4.764152, 4.790324, 4.822191, 4.855091, 4.886513, 4.913769, 
    4.934159, 4.945316, 4.945704, 4.935174, 4.915422, 4.890007, 4.863766, 
    4.841733, 4.827977, 4.824899, 4.833127, 4.851935, 4.879796, 4.914845, 
    4.955168,
  // totalHeight(12,36, 0-49)
    5.111942, 5.084561, 5.055326, 5.025081, 4.994619, 4.964703, 4.936105, 
    4.909595, 4.885931, 4.865786, 4.849653, 4.83772, 4.829732, 4.824864, 
    4.821609, 4.804615, 4.794687, 4.792881, 4.786672, 4.776821, 4.764374, 
    4.754197, 4.742932, 4.733154, 4.727239, 4.726232, 4.731174, 4.742603, 
    4.760743, 4.7837, 4.808667, 4.838854, 4.868789, 4.896034, 4.918074, 
    4.932533, 4.937595, 4.932491, 4.91799, 4.896621, 4.872406, 4.850078, 
    4.833977, 4.827167, 4.831044, 4.845499, 4.8694, 4.901079, 4.938695, 
    4.980416,
  // totalHeight(12,37, 0-49)
    5.112801, 5.08544, 5.055923, 5.025138, 4.993912, 4.963036, 4.933292, 
    4.905466, 4.880316, 4.858521, 4.840577, 4.826664, 4.81651, 4.809246, 
    4.803285, 4.789212, 4.785302, 4.781154, 4.774646, 4.766088, 4.756061, 
    4.7495, 4.742392, 4.737138, 4.735608, 4.738574, 4.746701, 4.76024, 
    4.779102, 4.801551, 4.82479, 4.852537, 4.878767, 4.901183, 4.917546, 
    4.92596, 4.9253, 4.915676, 4.898742, 4.877671, 4.856634, 4.839904, 
    4.830922, 4.831695, 4.84272, 4.863298, 4.892019, 4.927155, 4.966915, 
    5.009552,
  // totalHeight(12,38, 0-49)
    5.117163, 5.089993, 5.060169, 5.028653, 4.996345, 4.964101, 4.932761, 
    4.903154, 4.876072, 4.852218, 4.83211, 4.815961, 4.803544, 4.794055, 
    4.786015, 4.774364, 4.77559, 4.770068, 4.763923, 4.757067, 4.749672, 
    4.746599, 4.743455, 4.742412, 4.744793, 4.75115, 4.761802, 4.776754, 
    4.795622, 4.81691, 4.837911, 4.862556, 4.884535, 4.90178, 4.912446, 
    4.915242, 4.909836, 4.897208, 4.879747, 4.860974, 4.844863, 4.834976, 
    4.833762, 4.842255, 4.86022, 4.886531, 4.919603, 4.957696, 4.999078, 
    5.042069,
  // totalHeight(12,39, 0-49)
    5.125264, 5.098615, 5.068628, 5.036368, 5.002841, 4.969013, 4.935816, 
    4.904154, 4.874874, 4.84872, 4.826249, 4.807725, 4.793006, 4.781432, 
    4.771742, 4.761746, 4.766644, 4.760505, 4.755105, 4.750071, 4.74527, 
    4.745384, 4.745862, 4.74859, 4.754327, 4.763429, 4.775914, 4.791576, 
    4.809772, 4.829317, 4.847673, 4.868758, 4.88626, 4.898421, 4.903902, 
    4.902092, 4.893451, 4.879701, 4.863706, 4.849003, 4.839085, 4.836678, 
    4.843287, 4.859147, 4.883482, 4.914883, 4.951668, 4.992102, 5.034494, 
    5.077206,
  // totalHeight(12,40, 0-49)
    5.136877, 5.111238, 5.081432, 5.048639, 5.014005, 4.978633, 4.943581, 
    4.909848, 4.878351, 4.849883, 4.825041, 4.804149, 4.787166, 4.773599, 
    4.76246, 4.753274, 4.760116, 4.753808, 4.749212, 4.745819, 4.743309, 
    4.746111, 4.749687, 4.755607, 4.764044, 4.775191, 4.788807, 4.804513, 
    4.821455, 4.83882, 4.854307, 4.871682, 4.884876, 4.892533, 4.893868, 
    4.888951, 4.878927, 4.866021, 4.853262, 4.843918, 4.840827, 4.845891, 
    4.859829, 4.882285, 4.912125, 4.94777, 4.987484, 5.029533, 5.072239, 
    5.113965,
  // totalHeight(12,41, 0-49)
    5.151308, 5.127309, 5.098226, 5.065358, 5.030005, 4.993429, 4.956825, 
    4.921301, 4.887843, 4.857288, 4.830274, 4.807172, 4.78804, 4.772555, 
    4.759991, 4.750806, 4.757907, 4.751545, 4.747518, 4.745323, 4.744565, 
    4.749381, 4.755365, 4.763759, 4.774164, 4.786629, 4.800695, 4.81586, 
    4.83112, 4.846073, 4.858711, 4.872571, 4.882043, 4.886209, 4.884839, 
    4.878588, 4.869079, 4.858769, 4.850559, 4.847245, 4.850982, 4.862956, 
    4.883301, 4.911276, 4.945533, 4.98441, 5.026139, 5.068966, 5.111191, 
    5.151146,
  // totalHeight(12,42, 0-49)
    5.167433, 5.145825, 5.118198, 5.085958, 5.05056, 5.013422, 4.975871, 
    4.939118, 4.904213, 4.872023, 4.84321, 4.818187, 4.797098, 4.779766, 
    4.765706, 4.755823, 4.761775, 4.755195, 4.751298, 4.749695, 4.749995, 
    4.756035, 4.763631, 4.773695, 4.7853, 4.798368, 4.81227, 4.826428, 
    4.839757, 4.852291, 4.862344, 4.873213, 4.879873, 4.881848, 4.879389, 
    4.873567, 4.866244, 4.859843, 4.856923, 4.859726, 4.86978, 4.887712, 
    4.91327, 4.945491, 4.982934, 5.023899, 5.066599, 5.109246, 5.150087, 
    5.187401,
  // totalHeight(12,43, 0-49)
    5.183809, 5.165433, 5.140165, 5.109489, 5.074985, 5.038198, 5.000572, 
    4.963393, 4.927755, 4.894545, 4.864434, 4.837869, 4.815063, 4.795979, 
    4.780333, 4.769211, 4.773004, 4.765872, 4.76158, 4.759906, 4.760523, 
    4.766987, 4.77537, 4.786294, 4.798351, 4.811367, 4.824594, 4.837421, 
    4.848752, 4.859057, 4.866989, 4.875616, 4.880549, 4.881706, 4.879692, 
    4.875801, 4.871909, 4.870196, 4.872773, 4.881325, 4.896852, 4.919589, 
    4.94904, 4.984147, 5.023449, 5.065253, 5.107759, 5.149135, 5.187568, 
    5.22127,
  // totalHeight(12,44, 0-49)
    5.198803, 5.184547, 5.162685, 5.134711, 5.102264, 5.066974, 5.03035, 
    4.993721, 4.9582, 4.924677, 4.893834, 4.866149, 4.841905, 4.821187, 
    4.803893, 4.791168, 4.792223, 4.784158, 4.778965, 4.776611, 4.77686, 
    4.783025, 4.79144, 4.802482, 4.814332, 4.826746, 4.838907, 4.85022, 
    4.859634, 4.868042, 4.874416, 4.881635, 4.88592, 4.887495, 4.887174, 
    4.886299, 4.886583, 4.889843, 4.897708, 4.911355, 4.931366, 4.957692, 
    4.989709, 5.026331, 5.066129, 5.10744, 5.148468, 5.187353, 5.222224, 
    5.251262,
  // totalHeight(12,45, 0-49)
    5.210752, 5.201502, 5.184183, 5.160196, 5.131147, 5.098663, 5.064255, 
    5.029252, 4.994759, 4.961669, 4.930681, 4.902313, 4.876929, 4.854733, 
    4.835791, 4.821271, 4.819385, 4.810057, 4.803559, 4.800041, 4.799366, 
    4.804659, 4.81249, 4.82304, 4.834153, 4.845552, 4.856387, 4.866125, 
    4.873801, 4.880695, 4.886077, 4.892675, 4.897229, 4.900172, 4.9024, 
    4.905163, 4.909904, 4.918032, 4.9307, 4.948648, 4.972125, 5.000875, 
    5.034193, 5.071006, 5.109934, 5.149368, 5.187541, 5.222595, 5.252655, 
    5.275915,
  // totalHeight(12,46, 0-49)
    5.218122, 5.214686, 5.20306, 5.184418, 5.160201, 5.131918, 5.101005, 
    5.068739, 5.036206, 5.004301, 4.973755, 4.945153, 4.91895, 4.895483, 
    4.874975, 4.858628, 4.853901, 4.843082, 4.835012, 4.830008, 4.828019, 
    4.832044, 4.838839, 4.848449, 4.858446, 4.868553, 4.87793, 4.886125, 
    4.892288, 4.898044, 4.902914, 4.909524, 4.915015, 4.919935, 4.925162, 
    4.93177, 4.940877, 4.953484, 4.970314, 4.991725, 5.017685, 5.047775, 
    5.081226, 5.116975, 5.153697, 5.189855, 5.223742, 5.253561, 5.277506, 
    5.293887,
  // totalHeight(12,47, 0-49)
    5.21968, 5.222688, 5.21781, 5.205827, 5.18786, 5.16517, 5.139026, 
    5.110605, 5.080956, 5.050987, 5.021486, 4.993125, 4.966475, 4.942011, 
    4.920112, 4.902047, 4.89479, 4.88238, 4.87262, 4.865965, 4.86244, 
    4.86497, 4.870446, 4.87882, 4.88747, 4.896142, 4.904027, 4.910778, 
    4.91566, 4.9206, 4.925312, 4.932374, 4.939193, 4.946368, 4.954691, 
    4.965012, 4.978126, 4.994638, 5.014892, 5.038917, 5.066428, 5.09685, 
    5.129348, 5.162853, 5.19609, 5.227598, 5.255783, 5.278975, 5.295548, 
    5.304067,
  // totalHeight(12,48, 0-49)
    5.214645, 5.224436, 5.227116, 5.222918, 5.212476, 5.196669, 5.176497, 
    5.152991, 5.127141, 5.099882, 5.07207, 5.044486, 5.017835, 4.992734, 
    4.969724, 4.950169, 4.940837, 4.926858, 4.91543, 4.907111, 4.90198, 
    4.902931, 4.906935, 4.913908, 4.921101, 4.9283, 4.934745, 4.940191, 
    4.944019, 4.94839, 4.953168, 4.960919, 4.969209, 4.978634, 4.989865, 
    5.003521, 5.020082, 5.039804, 5.062685, 5.088459, 5.11661, 5.146403, 
    5.176918, 5.207063, 5.235599, 5.261165, 5.28232, 5.297623, 5.305756, 
    5.305692,
  // totalHeight(12,49, 0-49)
    5.192284, 5.210041, 5.222421, 5.228807, 5.229014, 5.22324, 5.211989, 
    5.195982, 5.176065, 5.153151, 5.128168, 5.102034, 5.075628, 5.049784, 
    5.025281, 5.004552, 5.000236, 4.983833, 4.969202, 4.957649, 4.949624, 
    4.951151, 4.956371, 4.96534, 4.972784, 4.978915, 4.982822, 4.984548, 
    4.983208, 4.98358, 4.985592, 4.994268, 5.004465, 5.016714, 5.031483, 
    5.049073, 5.069549, 5.092734, 5.118204, 5.145324, 5.173291, 5.201159, 
    5.227886, 5.252362, 5.273417, 5.289875, 5.300619, 5.304664, 5.301308, 
    5.290269,
  // totalHeight(13,0, 0-49)
    5.302906, 5.297866, 5.283644, 5.261401, 5.232627, 5.198957, 5.162014, 
    5.123312, 5.084203, 5.045848, 5.009209, 4.975058, 4.943973, 4.916348, 
    4.892391, 4.872317, 4.857236, 4.844203, 4.834624, 4.828238, 4.824745, 
    4.82422, 4.826094, 4.830255, 4.836333, 4.844073, 4.853085, 4.862946, 
    4.873157, 4.88348, 4.893552, 4.903595, 4.913329, 4.923114, 4.933573, 
    4.945522, 4.959881, 4.977537, 4.999209, 5.025342, 5.056015, 5.090916, 
    5.129323, 5.170135, 5.211916, 5.252959, 5.291361, 5.325141, 5.352355, 
    5.371239,
  // totalHeight(13,1, 0-49)
    5.28951, 5.280722, 5.263025, 5.237669, 5.206186, 5.170209, 5.131349, 
    5.091095, 5.05077, 5.011506, 4.974237, 4.939699, 4.908432, 4.880779, 
    4.856899, 4.837128, 4.823848, 4.810921, 4.801519, 4.795393, 4.792206, 
    4.792432, 4.795098, 4.800194, 4.807179, 4.81584, 4.825731, 4.836394, 
    4.847203, 4.858047, 4.868423, 4.878859, 4.888578, 4.897897, 4.907441, 
    4.918092, 4.930884, 4.946864, 4.966928, 4.991677, 5.021327, 5.055649, 
    5.093979, 5.135242, 5.178015, 5.220617, 5.26118, 5.297764, 5.328457, 
    5.351484,
  // totalHeight(13,2, 0-49)
    5.270072, 5.257787, 5.237234, 5.209664, 5.176543, 5.139416, 5.099804, 
    5.059119, 5.018622, 4.979402, 4.942351, 4.90817, 4.877359, 4.850216, 
    4.826835, 4.807679, 4.796417, 4.78367, 4.774438, 4.768469, 4.765407, 
    4.766132, 4.769279, 4.774964, 4.782534, 4.791835, 4.802403, 4.813765, 
    4.825194, 4.836684, 4.847581, 4.858711, 4.868759, 4.877928, 4.886779, 
    4.896184, 4.907245, 4.921134, 4.938916, 4.961381, 4.988906, 5.021394, 
    5.058273, 5.098534, 5.14082, 5.18352, 5.224868, 5.263035, 5.29622, 
    5.322726,
  // totalHeight(13,3, 0-49)
    5.246368, 5.230927, 5.208125, 5.179145, 5.145323, 5.108055, 5.068716, 
    5.028602, 4.988883, 4.950584, 4.914549, 4.881436, 4.851695, 4.825564, 
    4.803069, 4.78479, 4.775711, 4.763161, 4.754032, 4.748058, 4.744871, 
    4.745768, 4.749006, 4.754856, 4.762612, 4.77221, 4.783199, 4.795122, 
    4.807179, 4.819442, 4.831099, 4.843277, 4.85408, 4.863536, 4.872057, 
    4.880424, 4.889727, 4.901223, 4.916138, 4.935462, 4.959786, 4.989203, 
    5.023292, 5.061168, 5.10159, 5.143067, 5.183972, 5.222636, 5.257412, 
    5.286727,
  // totalHeight(13,4, 0-49)
    5.220337, 5.202127, 5.177616, 5.147886, 5.114111, 5.077507, 5.039276, 
    5.000571, 4.962453, 4.925858, 4.89157, 4.860184, 4.83209, 4.80745, 
    4.786195, 4.768989, 4.762178, 4.749801, 4.740659, 4.734465, 4.730842, 
    4.731516, 4.734381, 4.73989, 4.747362, 4.756843, 4.767935, 4.780223, 
    4.792881, 4.806018, 4.818665, 4.832267, 4.844315, 4.854602, 4.863307, 
    4.871026, 4.878742, 4.887725, 4.899331, 4.91477, 4.934896, 4.960064, 
    4.990092, 5.024294, 5.061602, 5.100693, 5.140108, 5.178351, 5.21394, 
    5.245433,
  // totalHeight(13,5, 0-49)
    5.193888, 5.173308, 5.147536, 5.117548, 5.084359, 5.048999, 5.012493, 
    4.975842, 4.939978, 4.905743, 4.873834, 4.84477, 4.818851, 4.796136, 
    4.776439, 4.760425, 4.755842, 4.743599, 4.734304, 4.72764, 4.723233, 
    4.723243, 4.725216, 4.729818, 4.736472, 4.745353, 4.756155, 4.768545, 
    4.781706, 4.795761, 4.809578, 4.824949, 4.838744, 4.850475, 4.860016, 
    4.867673, 4.874217, 4.880829, 4.88893, 4.899941, 4.915029, 4.9349, 
    4.959711, 4.989072, 5.022166, 5.057874, 5.094924, 5.131988, 5.167728, 
    5.200819,
  // totalHeight(13,6, 0-49)
    5.168723, 5.146162, 5.119484, 5.089571, 5.057295, 5.023526, 4.989129, 
    4.954954, 4.92181, 4.890425, 4.861399, 4.835148, 4.811861, 4.791458, 
    4.773588, 4.758794, 4.756223, 4.744107, 4.734529, 4.727149, 4.721606, 
    4.720503, 4.721052, 4.724154, 4.729415, 4.737158, 4.74721, 4.759347, 
    4.772826, 4.78774, 4.802809, 4.820201, 4.836185, 4.849976, 4.861088, 
    4.869447, 4.875493, 4.880192, 4.884932, 4.891296, 4.900784, 4.914537, 
    4.933163, 4.956684, 4.984612, 5.016095, 5.050054, 5.085308, 5.12063, 
    5.154777,
  // totalHeight(13,7, 0-49)
    5.146191, 5.122014, 5.094694, 5.065038, 5.033816, 5.001769, 4.969636, 
    4.938137, 4.907962, 4.879731, 4.853929, 4.830854, 4.810551, 4.792776, 
    4.776973, 4.763321, 4.762328, 4.750426, 4.740496, 4.732202, 4.72523, 
    4.722604, 4.721231, 4.72226, 4.725554, 4.73159, 4.740366, 4.751813, 
    4.765307, 4.780891, 4.797148, 4.816651, 4.835127, 4.851506, 4.864916, 
    4.874842, 4.881288, 4.884869, 4.886801, 4.888733, 4.892467, 4.899627, 
    4.911375, 4.928267, 4.950256, 4.976807, 5.007057, 5.039953, 5.074344, 
    5.109021,
  // totalHeight(13,8, 0-49)
    5.12719, 5.101721, 5.073936, 5.044599, 5.01441, 4.984032, 4.95411, 
    4.92527, 4.898105, 4.873127, 4.850711, 4.831019, 4.81394, 4.799034, 
    4.785518, 4.77283, 4.772757, 4.761313, 4.751078, 4.74178, 4.733187, 
    4.728723, 4.725017, 4.723469, 4.724253, 4.728013, 4.734952, 4.745189, 
    4.758284, 4.7742, 4.791411, 4.812908, 4.833974, 4.853284, 4.869596, 
    4.881938, 4.889804, 4.893339, 4.893427, 4.891637, 4.889973, 4.890526, 
    4.895082, 4.90484, 4.920309, 4.941354, 4.96736, 4.997399, 5.030363, 
    5.06504,
  // totalHeight(13,9, 0-49)
    5.112118, 5.085622, 5.057474, 5.028415, 4.999117, 4.970207, 4.94228, 
    4.915903, 4.891597, 4.869787, 4.850737, 4.834479, 4.820738, 4.808884, 
    4.7979, 4.785911, 4.785915, 4.775369, 4.765037, 4.754792, 4.744537, 
    4.73805, 4.731728, 4.727205, 4.725008, 4.725948, 4.730473, 4.738923, 
    4.7511, 4.766879, 4.784646, 4.8078, 4.831308, 4.853636, 4.873232, 
    4.888683, 4.898961, 4.903659, 4.903191, 4.898856, 4.892699, 4.88718, 
    4.884699, 4.887177, 4.895783, 4.910887, 4.932183, 4.958889, 4.989927, 
    5.024058,
  // totalHeight(13,10, 0-49)
    5.100892, 5.073568, 5.045088, 5.016195, 4.987566, 4.959826, 4.933566, 
    4.909325, 4.887583, 4.868696, 4.852839, 4.839923, 4.829534, 4.820874, 
    4.812728, 4.801129, 4.800285, 4.791276, 4.781237, 4.770275, 4.758482, 
    4.749933, 4.740851, 4.733079, 4.727515, 4.725141, 4.726683, 4.732738, 
    4.743409, 4.758473, 4.776271, 4.800553, 4.826117, 4.851284, 4.874251, 
    4.893243, 4.906741, 4.913769, 4.914171, 4.908805, 4.899549, 4.88904, 
    4.880201, 4.875673, 4.877369, 4.886271, 4.902476, 4.925397, 4.954008, 
    4.987036,
  // totalHeight(13,11, 0-49)
    5.093023, 5.064999, 5.036164, 5.007285, 4.979065, 4.952162, 4.927186, 
    4.904684, 4.885119, 4.868808, 4.855855, 4.846086, 4.838981, 4.833637, 
    4.828726, 4.817231, 4.814683, 4.807994, 4.798809, 4.787527, 4.774482, 
    4.76396, 4.75211, 4.74093, 4.731703, 4.725581, 4.723604, 4.726661, 
    4.7352, 4.748919, 4.766147, 4.790886, 4.817931, 4.845511, 4.87165, 
    4.894293, 4.911518, 4.921821, 4.924446, 4.919686, 4.909037, 4.895079, 
    4.881061, 4.870255, 4.86534, 4.868004, 4.878853, 4.897589, 4.923282, 
    4.954648,
  // totalHeight(13,12, 0-49)
    5.087749, 5.05909, 5.029847, 5.00082, 4.972756, 4.946362, 4.92229, 
    4.901118, 4.883312, 4.869174, 4.858771, 4.851879, 4.847934, 4.846014, 
    4.844818, 4.833281, 4.828422, 4.824882, 4.817225, 4.80616, 4.792282, 
    4.779981, 4.765455, 4.75081, 4.737704, 4.727466, 4.721484, 4.720968, 
    4.72675, 4.738482, 4.754528, 4.778989, 4.806825, 4.836215, 4.865081, 
    4.891179, 4.912287, 4.926467, 4.932404, 4.92977, 4.919513, 4.903913, 
    4.886283, 4.870348, 4.859491, 4.856153, 4.861555, 4.875796, 4.898129, 
    4.927302,
  // totalHeight(13,13, 0-49)
    5.084192, 5.054919, 5.025204, 4.995886, 4.967764, 4.941601, 4.918097, 
    4.897873, 4.881418, 4.86904, 4.860798, 4.856464, 4.8555, 4.857069, 
    4.860056, 4.848661, 4.84133, 4.84169, 4.836272, 4.826051, 4.811856, 
    4.798031, 4.780994, 4.762904, 4.745772, 4.731121, 4.720706, 4.716094, 
    4.718533, 4.727675, 4.741975, 4.765423, 4.793318, 4.823824, 4.854806, 
    4.883918, 4.908742, 4.927023, 4.936974, 4.937667, 4.929421, 4.914011, 
    4.894545, 4.874947, 4.859157, 4.850342, 4.850424, 4.860008, 4.878631, 
    4.905142,
  // totalHeight(13,14, 0-49)
    5.081517, 5.05163, 5.021392, 4.991681, 4.963344, 4.937195, 4.913986, 
    4.89438, 4.878895, 4.867865, 4.861372, 4.85923, 4.860987, 4.865987, 
    4.87346, 4.863003, 4.853669, 4.858477, 4.855946, 4.847213, 4.833271, 
    4.818205, 4.798866, 4.777408, 4.756172, 4.736881, 4.721683, 4.712525, 
    4.7111, 4.717124, 4.729209, 4.750969, 4.778223, 4.809133, 4.841548, 
    4.873077, 4.901201, 4.923458, 4.937708, 4.942506, 4.937534, 4.923936, 
    4.904391, 4.882751, 4.863289, 4.849806, 4.844934, 4.849881, 4.864576, 
    4.888054,
  // totalHeight(13,15, 0-49)
    5.079049, 5.048556, 5.017774, 4.987615, 4.958967, 4.932677, 4.909543, 
    4.890262, 4.875388, 4.865291, 4.8601, 4.859703, 4.863788, 4.871943, 
    4.883821, 4.876032, 4.865983, 4.875477, 4.876322, 4.869667, 4.856545, 
    4.840522, 4.819111, 4.794412, 4.769051, 4.744977, 4.724737, 4.710681, 
    4.704965, 4.707441, 4.716984, 4.73648, 4.762472, 4.793127, 4.826293, 
    4.859575, 4.890423, 4.916268, 4.934734, 4.94397, 4.943079, 4.932546, 
    4.914461, 4.892363, 4.870615, 4.853478, 4.844249, 4.844784, 4.855497, 
    4.875701,
  // totalHeight(13,16, 0-49)
    5.076357, 5.04529, 5.013985, 4.983371, 4.954356, 4.927814, 4.90456, 
    4.885322, 4.870687, 4.861065, 4.85665, 4.857431, 4.863256, 4.873969, 
    4.889624, 4.887436, 4.878976, 4.892997, 4.897475, 4.893355, 4.881554, 
    4.864819, 4.841561, 4.813771, 4.784333, 4.755423, 4.729992, 4.710805, 
    4.700493, 4.699131, 4.705956, 4.722753, 4.746984, 4.776818, 4.810111, 
    4.844488, 4.877415, 4.906292, 4.928608, 4.942223, 4.945766, 4.939097, 
    4.923651, 4.902481, 4.879802, 4.860133, 4.84732, 4.843862, 4.850718, 
    4.867552,
  // totalHeight(13,17, 0-49)
    5.073276, 5.041718, 5.00995, 4.978906, 4.949494, 4.922585, 4.899002, 
    4.879483, 4.864644, 4.854941, 4.850645, 4.851858, 4.858593, 4.870928, 
    4.889231, 4.896774, 4.893412, 4.911368, 4.919476, 4.918165, 4.908042, 
    4.890761, 4.865815, 4.835064, 4.801618, 4.767901, 4.737255, 4.712861, 
    4.697815, 4.692492, 4.696613, 4.710435, 4.732548, 4.761121, 4.794013, 
    4.828882, 4.86324, 4.894509, 4.920127, 4.937771, 4.94571, 4.943258, 
    4.931211, 4.912036, 4.889621, 4.86853, 4.853006, 4.846128, 4.849413, 
    4.862942,
  // totalHeight(13,18, 0-49)
    5.069894, 5.037993, 5.005871, 4.974439, 4.94458, 4.917144, 4.89294, 
    4.872707, 4.857082, 4.846572, 4.841537, 4.842215, 4.848804, 4.861626, 
    4.881323, 4.903514, 4.910012, 4.930978, 4.94249, 4.944072, 4.935783, 
    4.917948, 4.891298, 4.857579, 4.820136, 4.781682, 4.745924, 4.716439, 
    4.696753, 4.687572, 4.689219, 4.699979, 4.719781, 4.746784, 4.778859, 
    4.813701, 4.848888, 4.881894, 4.910168, 4.931293, 4.943286, 4.945026, 
    4.936729, 4.920257, 4.899048, 4.877536, 4.860189, 4.850558, 4.850698, 
    4.861127,
  // totalHeight(13,19, 0-49)
    5.066533, 5.034526, 5.002198, 4.970406, 4.939985, 4.911748, 4.886477, 
    4.864903, 4.847689, 4.835394, 4.828495, 4.827422, 4.832679, 4.845, 
    4.865422, 4.907155, 4.92915, 4.952248, 4.966908, 4.971374, 4.964861, 
    4.946195, 4.917465, 4.88041, 4.838736, 4.795547, 4.754904, 4.720706, 
    4.696789, 4.684154, 4.683802, 4.691631, 4.709097, 4.734366, 4.765323, 
    4.799715, 4.83519, 4.869302, 4.899551, 4.923498, 4.939002, 4.944619, 
    4.940077, 4.926665, 4.907319, 4.886206, 4.86786, 4.856178, 4.853689, 
    4.861349,
  // totalHeight(13,20, 0-49)
    5.062326, 5.029428, 4.996673, 4.965066, 4.935573, 4.909109, 4.88653, 
    4.868585, 4.85582, 4.848474, 4.846332, 4.848631, 4.854045, 4.860835, 
    4.867209, 30, 4.960554, 4.96489, 4.966611, 4.9642, 4.956264, 4.938369, 
    4.913416, 4.881072, 4.843659, 4.803276, 4.763498, 4.72832, 4.70213, 
    4.68676, 4.684481, 4.689006, 4.70359, 4.72649, 4.755638, 4.788839, 
    4.823808, 4.858182, 4.88953, 4.915427, 4.93366, 4.942553, 4.941444, 
    4.931111, 4.913975, 4.893856, 4.875212, 4.86215, 4.857589, 4.862891,
  // totalHeight(13,21, 0-49)
    5.05939, 5.026729, 4.99416, 4.962648, 4.9331, 4.906367, 4.883225, 
    4.864333, 4.850152, 4.840854, 4.836205, 4.83551, 4.837572, 4.840788, 
    4.843318, 30, 4.988412, 4.991874, 4.992982, 4.989769, 4.980573, 4.958037, 
    4.92908, 4.892868, 4.851937, 4.808477, 4.766072, 4.728681, 4.700647, 
    4.683903, 4.681386, 4.684261, 4.697501, 4.719358, 4.747776, 4.780595, 
    4.815596, 4.850495, 4.882943, 4.910565, 4.93112, 4.942796, 4.944633, 
    4.936992, 4.921839, 4.902638, 4.883723, 4.869337, 4.862715, 4.865593,
  // totalHeight(13,22, 0-49)
    5.056715, 5.024198, 4.991746, 4.960288, 4.930684, 4.903732, 4.880151, 
    4.860536, 4.845291, 4.834549, 4.828082, 4.825235, 4.824912, 4.825584, 
    4.825378, 30, 5.007531, 5.01016, 5.010991, 5.007695, 4.998391, 4.972798, 
    4.941637, 4.903322, 4.860387, 4.814988, 4.770687, 4.731456, 4.701693, 
    4.683507, 4.680566, 4.681566, 4.693231, 4.713815, 4.741263, 4.773442, 
    4.808179, 4.843255, 4.876388, 4.905256, 4.92762, 4.941576, 4.94595, 
    4.940767, 4.927596, 4.90955, 4.890788, 4.875599, 4.867455, 4.868394,
  // totalHeight(13,23, 0-49)
    5.054629, 5.022224, 4.989868, 4.958463, 4.928839, 4.901758, 4.877898, 
    4.857814, 4.841877, 4.830197, 4.822548, 4.818313, 4.816451, 4.815497, 
    4.813565, 30, 5.020011, 5.021922, 5.022535, 5.019291, 5.010156, 4.982364, 
    4.949795, 4.910171, 4.86599, 4.819386, 4.773896, 4.733502, 4.702621, 
    4.683495, 4.680393, 4.679896, 4.690282, 4.709814, 4.73644, 4.768047, 
    4.802501, 4.837631, 4.871211, 4.900962, 4.924655, 4.940331, 4.946666, 
    4.94344, 4.931912, 4.914906, 4.89641, 4.880715, 4.871446, 4.870869,
  // totalHeight(13,24, 0-49)
    5.053342, 5.021052, 4.988799, 4.957475, 4.927895, 4.900801, 4.876853, 
    4.856582, 4.840339, 4.828224, 4.820012, 4.8151, 4.812484, 4.810732, 
    4.807968, 30, 5.026357, 5.027834, 5.028316, 5.025136, 5.016194, 4.987086, 
    4.953739, 4.913423, 4.868618, 4.821458, 4.775474, 4.734633, 4.703346, 
    4.683897, 4.680958, 4.67964, 4.689296, 4.708194, 4.734291, 4.765488, 
    4.799673, 4.834713, 4.868412, 4.898533, 4.92286, 4.939422, 4.946823, 
    4.944707, 4.934157, 4.91782, 4.899562, 4.883654, 4.873792, 4.872372,
  // totalHeight(13,25, 0-49)
    5.052937, 5.020776, 4.988652, 4.957452, 4.927993, 4.901019, 4.877185, 
    4.857019, 4.840869, 4.828824, 4.820656, 4.815761, 4.813137, 4.811367, 
    4.80859, 30, 5.026131, 5.027595, 5.028104, 5.025001, 5.016189, 4.986772, 
    4.953303, 4.912925, 4.868127, 4.821061, 4.775249, 4.73463, 4.703572, 
    4.684343, 4.681725, 4.680303, 4.68982, 4.708557, 4.734481, 4.76551, 
    4.799545, 4.834464, 4.868091, 4.898201, 4.922594, 4.939297, 4.946908, 
    4.945036, 4.934718, 4.918549, 4.900354, 4.884392, 4.874371, 4.872713,
  // totalHeight(13,26, 0-49)
    5.053365, 5.021352, 4.989378, 4.958348, 4.92909, 4.902367, 4.878851, 
    4.859085, 4.843421, 4.831948, 4.824425, 4.82023, 4.81834, 4.817324, 
    4.815344, 30, 5.019228, 5.021117, 5.02184, 5.018843, 5.010098, 4.981457, 
    4.948575, 4.908823, 4.864714, 4.818419, 4.773448, 4.7337, 4.703471, 
    4.684952, 4.682744, 4.681938, 4.691911, 4.710961, 4.737072, 4.768174, 
    4.802174, 4.836944, 4.870301, 4.900016, 4.923895, 4.939982, 4.946925, 
    4.944401, 4.933534, 4.917, 4.89867, 4.8828, 4.873055, 4.871789,
  // totalHeight(13,27, 0-49)
    5.054453, 5.022583, 4.990769, 4.959939, 4.930949, 4.904599, 4.881593, 
    4.862506, 4.847711, 4.837303, 4.831028, 4.82823, 4.827834, 4.828379, 
    4.828067, 30, 5.005809, 5.008458, 5.00954, 5.006703, 4.998044, 4.971261, 
    4.939735, 4.901355, 4.858659, 4.813832, 4.770372, 4.732119, 4.703287, 
    4.685929, 4.684206, 4.684655, 4.695604, 4.715379, 4.741986, 4.773363, 
    4.807406, 4.841971, 4.874848, 4.903781, 4.926571, 4.941309, 4.946741, 
    4.942723, 4.93059, 4.913219, 4.894607, 4.879008, 4.86998, 4.869713,
  // totalHeight(13,28, 0-49)
    5.055897, 5.024127, 4.992451, 4.961824, 4.933147, 4.907266, 4.884938, 
    4.866787, 4.853227, 4.844376, 4.839968, 4.839299, 4.841219, 4.844214, 
    4.846556, 30, 4.986444, 4.989986, 4.991482, 4.988878, 4.980467, 4.956567, 
    4.927253, 4.891089, 4.850602, 4.80798, 4.766706, 4.730566, 4.703684, 
    4.687934, 4.686851, 4.689076, 4.701419, 4.722225, 4.749526, 4.781257, 
    4.815298, 4.849463, 4.8815, 4.909118, 4.930127, 4.942695, 4.945752, 
    4.939439, 4.925432, 4.906913, 4.88804, 4.873039, 4.865275, 4.866679,
  // totalHeight(13,29, 0-49)
    5.057277, 5.025501, 4.993886, 4.963425, 4.935068, 4.909718, 4.888201, 
    4.871215, 4.859243, 4.852449, 4.850572, 4.852848, 4.858019, 4.864477, 
    4.870577, 30, 4.960837, 4.965211, 4.967146, 4.96498, 4.957272, 4.937307, 
    4.911318, 4.878489, 4.841214, 4.801627, 4.763185, 4.72964, 4.705064, 
    4.691149, 4.690714, 4.694875, 4.708726, 4.730634, 4.758652, 4.790708, 
    4.824646, 4.858231, 4.889145, 4.915062, 4.933808, 4.943669, 4.943821, 
    4.934777, 4.918635, 4.898928, 4.87997, 4.865904, 4.859822, 4.863319,
  // totalHeight(13,30, 0-49)
    5.059418, 5.028654, 4.997622, 4.96715, 4.938057, 4.911136, 4.887138, 
    4.866747, 4.850553, 4.839038, 4.832601, 4.831628, 4.836618, 4.848354, 
    4.867994, 4.90837, 4.928143, 4.951606, 4.967244, 4.973113, 4.968354, 
    4.949694, 4.92203, 4.886323, 4.846043, 4.804104, 4.764419, 4.730797, 
    4.707057, 4.694342, 4.694369, 4.700532, 4.715995, 4.739077, 4.76782, 
    4.800131, 4.833815, 4.866575, 4.896039, 4.919852, 4.935893, 4.942627, 
    4.93956, 4.927652, 4.909478, 4.888913, 4.870369, 4.857808, 4.853965, 
    4.860042,
  // totalHeight(13,31, 0-49)
    5.060282, 5.029759, 4.999126, 4.96925, 4.940992, 4.915175, 4.892564, 
    4.873836, 4.859542, 4.850095, 4.845772, 4.846765, 4.85328, 4.865714, 
    4.884841, 4.905748, 4.911053, 4.932447, 4.945031, 4.948086, 4.941575, 
    4.923994, 4.898461, 4.866093, 4.830063, 4.792876, 4.758057, 4.729052, 
    4.709362, 4.699802, 4.701348, 4.710032, 4.727447, 4.751931, 4.781534, 
    4.814127, 4.847456, 4.879147, 4.906764, 4.927947, 4.940672, 4.94366, 
    4.936833, 4.921684, 4.90129, 4.879853, 4.861801, 4.850834, 4.849262, 
    4.857854,
  // totalHeight(13,32, 0-49)
    5.060558, 5.030423, 5.000259, 4.970952, 4.943376, 4.918372, 4.896713, 
    4.879066, 4.865955, 4.857725, 4.854555, 4.856493, 4.863556, 4.875896, 
    4.894008, 4.900531, 4.896977, 4.915523, 4.924882, 4.9252, 4.916963, 
    4.900275, 4.876549, 4.847143, 4.815058, 4.782508, 4.752657, 4.728541, 
    4.713242, 4.707185, 4.710644, 4.721965, 4.741295, 4.766997, 4.797129, 
    4.829546, 4.861939, 4.891879, 4.916902, 4.9347, 4.943443, 4.94221, 
    4.931443, 4.913217, 4.891095, 4.869491, 4.85271, 4.844056, 4.845331, 
    4.856855,
  // totalHeight(13,33, 0-49)
    5.059862, 5.03015, 5.000467, 4.971692, 4.944696, 4.920317, 4.899325, 
    4.882373, 4.869952, 4.862354, 4.859664, 4.861796, 4.868586, 4.879933, 
    4.896007, 4.893321, 4.885574, 4.900522, 4.906545, 4.904282, 4.894521, 
    4.878765, 4.856861, 4.8304, 4.802221, 4.774295, 4.749418, 4.730218, 
    4.719326, 4.716811, 4.722351, 4.736221, 4.757266, 4.783872, 4.814105, 
    4.845798, 4.876605, 4.904065, 4.925737, 4.939448, 4.943662, 4.93793, 
    4.923305, 4.902457, 4.879358, 4.858486, 4.843853, 4.838239, 4.842885, 
    4.857669,
  // totalHeight(13,34, 0-49)
    5.058055, 5.028715, 4.999457, 4.971143, 4.944623, 4.920722, 4.900189, 
    4.883659, 4.871587, 4.864218, 4.861553, 4.863379, 4.869329, 4.879015, 
    4.892175, 4.88469, 4.876192, 4.887134, 4.889908, 4.885369, 4.874451, 
    4.859777, 4.839851, 4.816452, 4.79222, 4.768898, 4.748909, 4.734482, 
    4.727811, 4.728682, 4.736307, 4.752478, 4.774912, 4.802001, 4.831811, 
    4.862161, 4.890678, 4.914915, 4.93252, 4.941554, 4.94089, 4.930667, 
    4.912594, 4.889904, 4.866834, 4.847734, 4.836153, 4.834247, 4.842685, 
    4.860934,
  // totalHeight(13,35, 0-49)
    5.055274, 5.02619, 4.997241, 4.969266, 4.943089, 4.919506, 4.899241, 
    4.882901, 4.870915, 4.863482, 4.860535, 4.861737, 4.866537, 4.874239, 
    4.884109, 4.875016, 4.868087, 4.875023, 4.874868, 4.868522, 4.85693, 
    4.843543, 4.825792, 4.805592, 4.785332, 4.766533, 4.751252, 4.741336, 
    4.738557, 4.742521, 4.752098, 4.770198, 4.793586, 4.820644, 4.849438, 
    4.87777, 4.90328, 4.923584, 4.936518, 4.940488, 4.934902, 4.920564, 
    4.899837, 4.876399, 4.854555, 4.838321, 4.830633, 4.832978, 4.845473, 
    4.86724,
  // totalHeight(13,36, 0-49)
    5.051935, 5.022963, 4.994163, 4.966357, 4.940342, 4.916883, 4.896673, 
    4.880292, 4.868145, 4.860397, 4.856926, 4.857306, 4.860819, 4.866513, 
    4.873233, 4.864482, 4.860516, 4.863798, 4.861239, 4.853672, 4.841947, 
    4.830064, 4.814686, 4.797793, 4.781472, 4.767046, 4.756203, 4.750443, 
    4.751133, 4.757798, 4.76908, 4.788637, 4.812456, 4.838905, 4.86604, 
    4.891673, 4.9135, 4.929286, 4.937158, 4.935996, 4.925839, 4.908185, 
    4.885969, 4.863123, 4.843789, 4.831448, 4.828336, 4.835277, 4.851907, 
    4.87708,
  // totalHeight(13,37, 0-49)
    5.048712, 5.019714, 4.990895, 4.963061, 4.936992, 4.91342, 4.893018, 
    4.876333, 4.863755, 4.855429, 4.851202, 4.850588, 4.852764, 4.856591, 
    4.860627, 4.853176, 4.852786, 4.853034, 4.848742, 4.840593, 4.829271, 
    4.819106, 4.806266, 4.79274, 4.780269, 4.769989, 4.763242, 4.761208, 
    4.764874, 4.773776, 4.78642, 4.806883, 4.830554, 4.855775, 4.880613, 
    4.902925, 4.920528, 4.931437, 4.934191, 4.928248, 4.914334, 4.894584, 
    4.87234, 4.851547, 4.83594, 4.828331, 4.830231, 4.841869, 4.862504, 
    4.890805,
  // totalHeight(13,38, 0-49)
    5.046463, 5.017363, 4.988382, 4.960333, 4.933984, 4.910048, 4.889175, 
    4.871894, 4.858581, 4.849375, 4.84412, 4.842312, 4.843084, 4.84521, 
    4.847122, 4.841239, 4.84439, 4.842373, 4.837064, 4.828948, 4.818515, 
    4.810253, 4.800081, 4.789934, 4.781161, 4.774736, 4.771679, 4.772884, 
    4.778982, 4.789603, 4.803183, 4.82395, 4.846866, 4.87026, 4.892232, 
    4.910744, 4.923823, 4.92984, 4.927855, 4.917969, 4.901567, 4.881282, 
    4.860622, 4.843279, 4.832405, 4.830073, 4.83712, 4.853296, 4.877594, 
    4.908586,
  // totalHeight(13,39, 0-49)
    5.046107, 5.016935, 4.987735, 4.959342, 4.932527, 4.907993, 4.886375, 
    4.86819, 4.853814, 4.843393, 4.836789, 4.833525, 4.832754, 4.833261, 
    4.833495, 4.82901, 4.835154, 4.83167, 4.826, 4.818432, 4.809279, 
    4.803062, 4.795628, 4.788808, 4.783522, 4.780604, 4.780778, 4.78469, 
    4.79264, 4.804419, 4.818454, 4.838909, 4.860484, 4.881526, 4.900217, 
    4.914691, 4.92329, 4.924838, 4.918981, 4.90646, 4.889201, 4.870115, 
    4.852602, 4.839882, 4.834409, 4.837548, 4.849568, 4.869874, 4.897309, 
    4.930414,
  // totalHeight(13,40, 0-49)
    5.048494, 5.019421, 4.990073, 4.961317, 4.933938, 4.90864, 4.886052, 
    4.866689, 4.850931, 4.838945, 4.830641, 4.8256, 4.823055, 4.82189, 
    4.82068, 4.817156, 4.825377, 4.821116, 4.815586, 4.808927, 4.801313, 
    4.797197, 4.792489, 4.788867, 4.786796, 4.786984, 4.789888, 4.795939, 
    4.805148, 4.817516, 4.831503, 4.85106, 4.870792, 4.889106, 4.904329, 
    4.914861, 4.919432, 4.917396, 4.908987, 4.895493, 4.879183, 4.862983, 
    4.84994, 4.842655, 4.842869, 4.851325, 4.86787, 4.891695, 4.921583, 
    4.956109,
  // totalHeight(13,41, 0-49)
    5.05427, 5.025635, 4.996369, 4.967378, 4.939467, 4.913352, 4.889659, 
    4.868913, 4.851506, 4.837645, 4.827295, 4.820136, 4.815523, 4.812502, 
    4.809849, 4.806692, 4.81588, 4.811314, 4.806209, 4.800623, 4.794641, 
    4.79257, 4.790468, 4.789821, 4.790624, 4.793467, 4.798572, 4.806185, 
    4.816072, 4.828482, 4.841944, 4.860108, 4.877642, 4.893072, 4.90494, 
    4.911988, 4.913404, 4.909066, 4.899735, 4.887073, 4.87345, 4.861562, 
    4.85393, 4.852476, 4.858293, 4.871628, 4.892047, 4.918634, 4.950186, 
    4.985343,
  // totalHeight(13,42, 0-49)
    5.063781, 5.036088, 5.007306, 4.978371, 4.950112, 4.923259, 4.898448, 
    4.876221, 4.856994, 4.841022, 4.828345, 4.818758, 4.811777, 4.806639, 
    4.802362, 4.798909, 4.80793, 4.803259, 4.798624, 4.794068, 4.789628, 
    4.789413, 4.789672, 4.791672, 4.794939, 4.799946, 4.806708, 4.815324, 
    4.825358, 4.837329, 4.84987, 4.866296, 4.881484, 4.894133, 4.903078, 
    4.907446, 4.906895, 4.90178, 4.893241, 4.883102, 4.873612, 4.867048, 
    4.865321, 4.869707, 4.880752, 4.898339, 4.921859, 4.950371, 4.982732, 
    5.017666,
  // totalHeight(13,43, 0-49)
    5.077024, 5.050926, 5.02318, 4.994742, 4.966463, 4.939089, 4.913278, 
    4.889596, 4.868496, 4.850291, 4.835114, 4.822883, 4.813281, 4.80576, 
    4.799586, 4.79519, 4.80303, 4.798201, 4.793865, 4.790109, 4.786953, 
    4.788271, 4.790523, 4.794739, 4.799999, 4.80666, 4.814556, 4.823662, 
    4.8334, 4.84456, 4.855913, 4.87045, 4.883365, 4.893603, 4.900323, 
    4.903059, 4.901888, 4.897532, 4.891333, 4.885078, 4.880715, 4.880008, 
    4.884263, 4.894188, 4.909894, 4.931011, 4.956826, 4.986413, 5.018707, 
    5.052526,
  // totalHeight(13,44, 0-49)
    5.09363, 5.069897, 5.04386, 5.016483, 4.988629, 4.96107, 4.934496, 
    4.909508, 4.886611, 4.866188, 4.848468, 4.833498, 4.82113, 4.811025, 
    4.802682, 4.796786, 4.802666, 4.797429, 4.793074, 4.789756, 4.787496, 
    4.789924, 4.7937, 4.79963, 4.806377, 4.814182, 4.822727, 4.831895, 
    4.841009, 4.85113, 4.861181, 4.873878, 4.884815, 4.893214, 4.898576, 
    4.900804, 4.900312, 4.898042, 4.895368, 4.893885, 4.895139, 4.900371, 
    4.910341, 4.925292, 4.945001, 4.968908, 4.996238, 5.026088, 5.057459, 
    5.089253,
  // totalHeight(13,45, 0-49)
    5.112896, 5.092362, 5.068785, 5.043111, 5.016217, 4.988903, 4.961903, 
    4.935873, 4.911382, 4.88889, 4.868727, 4.851068, 4.835922, 4.823139, 
    4.812431, 4.804618, 4.808037, 4.802051, 4.79729, 4.793986, 4.792167, 
    4.79523, 4.800014, 4.807119, 4.814841, 4.823317, 4.832101, 4.841004, 
    4.8493, 4.858297, 4.867085, 4.878168, 4.887572, 4.894811, 4.899705, 
    4.902462, 4.903721, 4.904501, 4.906074, 4.909746, 4.916643, 4.927522, 
    4.942692, 4.962025, 4.985044, 5.011038, 5.039169, 5.068532, 5.098169, 
    5.127051,
  // totalHeight(13,46, 0-49)
    5.133814, 5.117327, 5.096988, 5.073705, 5.048361, 5.021798, 4.994802, 
    4.968101, 4.942336, 4.918055, 4.895684, 4.87552, 4.857718, 4.842292, 
    4.829139, 4.81916, 4.819887, 4.812812, 4.807271, 4.803571, 4.801742, 
    4.80497, 4.81025, 4.818002, 4.826226, 4.834962, 4.843659, 4.852087, 
    4.859497, 4.867418, 4.875102, 4.884908, 4.893291, 4.900041, 4.905254, 
    4.909355, 4.913095, 4.917461, 4.923537, 4.932306, 4.944498, 4.960462, 
    4.980148, 5.003146, 5.028774, 5.056185, 5.084462, 5.112659, 5.139817, 
    5.164942,
  // totalHeight(13,47, 0-49)
    5.155118, 5.143477, 5.127144, 5.10696, 5.083807, 5.058568, 5.032099, 
    5.005201, 4.978597, 4.952922, 4.928703, 4.906341, 4.886123, 4.868207, 
    4.85265, 4.840416, 4.838448, 4.830011, 4.823393, 4.818952, 4.816723, 
    4.819705, 4.825018, 4.832941, 4.841257, 4.849924, 4.85831, 4.866159, 
    4.872729, 4.879717, 4.886525, 4.895436, 4.903288, 4.910117, 4.91623, 
    4.922192, 4.928778, 4.936869, 4.947312, 4.960783, 4.977658, 4.997964, 
    5.021375, 5.047264, 5.074781, 5.102951, 5.130748, 5.157147, 5.181139, 
    5.201734,
  // totalHeight(13,48, 0-49)
    5.17534, 5.169244, 5.157641, 5.141272, 5.120998, 5.09774, 5.072417, 
    5.045903, 5.019007, 4.992444, 4.966833, 4.942678, 4.920383, 4.900235, 
    4.882427, 4.867987, 4.863477, 4.85351, 4.845624, 4.840209, 4.837288, 
    4.839696, 4.844657, 4.852349, 4.860429, 4.868786, 4.876736, 4.884, 
    4.889857, 4.896114, 4.9023, 4.910675, 4.918396, 4.925701, 4.933056, 
    4.941097, 4.950563, 4.962187, 4.976577, 4.994122, 5.014909, 5.038708, 
    5.064978, 5.092928, 5.121566, 5.149796, 5.176466, 5.200438, 5.22062, 5.236,
  // totalHeight(13,49, 0-49)
    5.18919, 5.190837, 5.186273, 5.175988, 5.160712, 5.141308, 5.11869, 
    5.09377, 5.067405, 5.04039, 5.013444, 4.987204, 4.962228, 4.938995, 
    4.917903, 4.901022, 4.900822, 4.888001, 4.877112, 4.869137, 4.864331, 
    4.86836, 4.875689, 4.886596, 4.896372, 4.905116, 4.911828, 4.916348, 
    4.917615, 4.919777, 4.922395, 4.930235, 4.938002, 4.946137, 4.955254, 
    4.966011, 4.979034, 4.994824, 5.013668, 5.035591, 5.060346, 5.087408, 
    5.116018, 5.145223, 5.173903, 5.200845, 5.22479, 5.244488, 5.258783, 
    5.266685,
  // totalHeight(14,0, 0-49)
    5.229131, 5.206501, 5.178502, 5.14638, 5.111412, 5.074858, 5.037918, 
    5.001689, 4.967128, 4.935019, 4.905952, 4.880305, 4.858244, 4.839743, 
    4.824595, 4.812624, 4.804584, 4.797328, 4.792109, 4.788625, 4.78663, 
    4.786323, 4.787329, 4.789779, 4.793612, 4.798909, 4.805624, 4.813658, 
    4.822749, 4.832749, 4.84324, 4.854219, 4.865003, 4.875406, 4.885445, 
    4.89538, 4.905724, 4.917185, 4.930576, 4.94668, 4.966119, 4.989237, 
    5.016041, 5.046188, 5.079033, 5.113686, 5.149096, 5.184103, 5.21749, 
    5.247988,
  // totalHeight(14,1, 0-49)
    5.207026, 5.182279, 5.152763, 5.119683, 5.084245, 5.047626, 5.010942, 
    4.975212, 4.941328, 4.910021, 4.881835, 4.857101, 4.835941, 4.818269, 
    4.80382, 4.79253, 4.786399, 4.779195, 4.773937, 4.770339, 4.768142, 
    4.767947, 4.769014, 4.771609, 4.775563, 4.781028, 4.787959, 4.796264, 
    4.805616, 4.816019, 4.826934, 4.838686, 4.850087, 4.860837, 4.870841, 
    4.880264, 4.889561, 4.899436, 4.910755, 4.924414, 4.941188, 4.961601, 
    4.985838, 5.013726, 5.044766, 5.078192, 5.113054, 5.148269, 5.182673, 
    5.215027,
  // totalHeight(14,2, 0-49)
    5.183304, 5.15703, 5.12666, 5.093325, 5.058139, 5.022183, 4.986475, 
    4.951942, 4.919401, 4.889516, 4.862769, 4.839439, 4.819584, 4.803053, 
    4.789515, 4.779003, 4.774808, 4.767579, 4.762142, 4.758224, 4.755566, 
    4.755175, 4.755948, 4.758294, 4.761974, 4.767229, 4.774033, 4.782334, 
    4.791769, 4.802477, 4.813826, 4.826488, 4.838775, 4.850249, 4.860665, 
    4.870028, 4.878657, 4.887173, 4.896429, 4.907394, 4.921, 4.937978, 
    4.958755, 4.983394, 5.011603, 5.042788, 5.076122, 5.110613, 5.14515, 
    5.178529,
  // totalHeight(14,3, 0-49)
    5.159269, 5.132011, 5.101366, 5.068372, 5.034046, 4.999361, 4.965226, 
    4.932481, 4.901851, 4.873924, 4.849108, 4.82761, 4.809415, 4.794293, 
    4.781828, 4.772121, 4.769814, 4.762452, 4.756672, 4.752212, 4.748813, 
    4.747893, 4.747982, 4.749643, 4.752614, 4.757233, 4.763523, 4.771494, 
    4.780782, 4.791656, 4.803401, 4.817072, 4.830497, 4.84309, 4.854418, 
    4.864275, 4.872768, 4.880341, 4.887757, 4.896002, 4.906137, 4.919126, 
    4.935688, 4.956191, 4.980619, 5.008601, 5.039472, 5.072342, 5.106161, 
    5.139763,
  // totalHeight(14,4, 0-49)
    5.136073, 5.108289, 5.077836, 5.045656, 5.012658, 4.979708, 4.947617, 
    4.91712, 4.888855, 4.863318, 4.840836, 4.821526, 4.805284, 4.791785, 
    4.780509, 4.771574, 4.771007, 4.763416, 4.75714, 4.751925, 4.747519, 
    4.745743, 4.744758, 4.745288, 4.747094, 4.75062, 4.755964, 4.763226, 
    4.772083, 4.782914, 4.794947, 4.809652, 4.824399, 4.838461, 4.851204, 
    4.862165, 4.871171, 4.878408, 4.884452, 4.890225, 4.896865, 4.905565, 
    4.917366, 4.933001, 4.952807, 4.976699, 5.004219, 5.034612, 5.066907, 
    5.099984,
  // totalHeight(14,5, 0-49)
    5.114647, 5.08669, 5.056768, 5.025724, 4.994371, 4.96347, 4.933736, 
    4.905807, 4.880225, 4.857395, 4.837543, 4.82069, 4.806624, 4.794909, 
    4.784913, 4.776653, 4.77757, 4.769712, 4.76284, 4.756712, 4.751087, 
    4.748175, 4.745767, 4.744746, 4.744943, 4.746911, 4.750852, 4.756979, 
    4.765056, 4.775557, 4.787667, 4.803314, 4.819453, 4.835233, 4.849818, 
    4.862471, 4.872696, 4.88035, 4.885726, 4.889578, 4.893041, 4.89748, 
    4.90426, 4.914527, 4.929033, 4.948059, 4.97142, 4.998543, 5.028562, 
    5.060421,
  // totalHeight(14,6, 0-49)
    5.095639, 5.06775, 5.038558, 5.008825, 4.979269, 4.950567, 4.923344, 
    4.898149, 4.875429, 4.855488, 4.838451, 4.824225, 4.812485, 4.802677, 
    4.79404, 4.786319, 4.788359, 4.780312, 4.772842, 4.76574, 4.758781, 
    4.754543, 4.750437, 4.747506, 4.745694, 4.74566, 4.747729, 4.752261, 
    4.759154, 4.768952, 4.780826, 4.797183, 4.814626, 4.832209, 4.848913, 
    4.86374, 4.875854, 4.884737, 4.890322, 4.893084, 4.894041, 4.894635, 
    4.896505, 4.901212, 4.909982, 4.923539, 4.942053, 4.9652, 4.992265, 
    5.022275,
  // totalHeight(14,7, 0-49)
    5.079382, 5.051685, 5.023293, 4.994893, 4.967136, 4.940629, 4.915915, 
    4.893468, 4.873641, 4.856643, 4.842487, 4.830967, 4.821641, 4.813837, 
    4.806674, 4.799337, 4.802044, 4.794051, 4.786124, 4.778114, 4.769837, 
    4.764191, 4.758224, 4.753119, 4.748968, 4.746531, 4.746279, 4.748741, 
    4.754, 4.762649, 4.773867, 4.790557, 4.809045, 4.82832, 4.847221, 
    4.864514, 4.879047, 4.889917, 4.896648, 4.899345, 4.898779, 4.896335, 
    4.893821, 4.893167, 4.896089, 4.903821, 4.916978, 4.935566, 4.959084, 
    4.986681,
  // totalHeight(14,8, 0-49)
    5.065872, 5.038401, 5.01076, 4.983597, 4.95751, 4.933054, 4.910717, 
    4.890898, 4.87387, 4.859747, 4.848433, 4.839616, 4.832747, 4.827052, 
    4.821545, 4.814451, 4.817304, 4.809798, 4.801712, 4.793008, 4.783563, 
    4.776557, 4.76869, 4.761254, 4.754529, 4.749352, 4.746367, 4.746292, 
    4.749443, 4.756443, 4.766504, 4.783024, 4.80213, 4.822789, 4.843732, 
    4.863547, 4.880808, 4.894256, 4.903001, 4.906718, 4.905815, 4.901471, 
    4.895508, 4.890118, 4.887469, 4.889338, 4.896865, 4.91048, 4.92997, 
    4.954655,
  // totalHeight(14,9, 0-49)
    5.054821, 5.027532, 5.000518, 4.974404, 4.949765, 4.927123, 4.906926, 
    4.889516, 4.875094, 4.863682, 4.855093, 4.848915, 4.84452, 4.841063, 
    4.837492, 4.83054, 4.83301, 4.826586, 4.818791, 4.809748, 4.799422, 
    4.791223, 4.781535, 4.77173, 4.762289, 4.754117, 4.748044, 4.744996, 
    4.74556, 4.750387, 4.75874, 4.774489, 4.79366, 4.815218, 4.837843, 
    4.859991, 4.880027, 4.896397, 4.907828, 4.913559, 4.913555, 4.908646, 
    4.9005, 4.891405, 4.883876, 4.880214, 4.88213, 4.890561, 4.905677, 
    4.927028,
  // totalHeight(14,10, 0-49)
    5.04573, 5.018534, 4.991975, 4.96668, 4.943219, 4.922101, 4.903752, 
    4.888469, 4.876389, 4.867462, 4.861423, 4.857787, 4.855875, 4.854819, 
    4.85357, 4.846726, 4.848333, 4.843694, 4.836761, 4.827849, 4.817042, 
    4.807907, 4.796583, 4.784479, 4.772281, 4.760951, 4.751504, 4.745098, 
    4.742626, 4.744754, 4.750842, 4.765165, 4.783755, 4.805612, 4.829389, 
    4.853467, 4.876074, 4.895433, 4.909956, 4.918473, 4.920488, 4.916383, 
    4.907503, 4.896041, 4.8847, 4.876213, 4.872857, 4.876142, 4.886695, 
    4.904379,
  // totalHeight(14,11, 0-49)
    5.038, 5.010782, 4.984499, 4.959789, 4.937232, 4.917344, 4.900531, 
    4.887064, 4.877037, 4.870335, 4.866637, 4.86542, 4.865989, 4.867517, 
    4.869044, 4.862404, 4.862796, 4.860651, 4.855209, 4.846973, 4.836166, 
    4.826419, 4.813724, 4.799486, 4.784587, 4.770025, 4.757013, 4.746933, 
    4.741017, 4.73996, 4.74325, 4.755486, 4.772819, 4.794303, 4.818602, 
    4.844064, 4.868836, 4.890996, 4.908724, 4.92051, 4.925418, 4.923341, 
    4.915177, 4.902844, 4.889031, 4.87675, 4.86878, 4.867208, 4.873197, 
    4.886992,
  // totalHeight(14,12, 0-49)
    5.031034, 5.003688, 4.977518, 4.953181, 4.931284, 4.912348, 4.896778, 
    4.884824, 4.876548, 4.871799, 4.870219, 4.871272, 4.8743, 4.878574, 
    4.883319, 4.877185, 4.876233, 4.87719, 4.873849, 4.866863, 4.856576, 
    4.846573, 4.832829, 4.816703, 4.799254, 4.781491, 4.764815, 4.750834, 
    4.741136, 4.736468, 4.736497, 4.746009, 4.761425, 4.781863, 4.806017, 
    4.832239, 4.858638, 4.883218, 4.904005, 4.919235, 4.927595, 4.928498, 
    4.922335, 4.910599, 4.895769, 4.880947, 4.869279, 4.863392, 4.865007, 
    4.874826,
  // totalHeight(14,13, 0-49)
    5.024333, 4.99677, 4.970584, 4.946457, 4.925018, 4.906796, 4.892203, 
    4.881479, 4.874665, 4.87159, 4.871881, 4.875025, 4.880433, 4.887527, 
    4.895803, 4.890821, 4.888721, 4.893181, 4.89245, 4.887251, 4.878012, 
    4.868104, 4.853672, 4.835969, 4.816206, 4.795377, 4.775051, 4.757049, 
    4.743318, 4.734697, 4.731096, 4.73732, 4.750211, 4.768974, 4.792344, 
    4.818688, 4.846123, 4.872623, 4.896131, 4.91471, 4.926751, 4.931248, 
    4.928075, 4.918214, 4.903775, 4.887743, 4.873465, 4.864006, 4.861628, 
    4.867535,
  // totalHeight(14,14, 0-49)
    5.017553, 4.989715, 4.963422, 4.939384, 4.918242, 4.90054, 4.88669, 
    4.876932, 4.871295, 4.869604, 4.871495, 4.876493, 4.884107, 4.893934, 
    4.905785, 4.903114, 4.900491, 4.908577, 4.910793, 4.907833, 4.900127, 
    4.890634, 4.875879, 4.856959, 4.835193, 4.811535, 4.787686, 4.765656, 
    4.747746, 4.734937, 4.727468, 4.729933, 4.739788, 4.756329, 4.778342, 
    4.804221, 4.832108, 4.85998, 4.88575, 4.90738, 4.923053, 4.931413, 
    4.931864, 4.92485, 4.912005, 4.896032, 4.880286, 4.868128, 4.8623, 
    4.864512,
  // totalHeight(14,15, 0-49)
    5.010522, 4.982379, 4.955929, 4.931895, 4.910927, 4.893575, 4.880256, 
    4.871205, 4.866455, 4.865833, 4.869004, 4.875539, 4.885052, 4.897312, 
    4.912402, 4.913854, 4.911866, 4.923392, 4.928685, 4.928277, 4.922505, 
    4.913686, 4.898948, 4.879184, 4.855774, 4.829604, 4.802463, 4.776515, 
    4.754398, 4.737293, 4.725864, 4.724226, 4.730651, 4.744537, 4.764725, 
    4.789639, 4.817448, 4.846156, 4.873679, 4.897934, 4.916968, 4.929162, 
    4.933515, 4.929967, 4.919626, 4.90479, 4.888655, 4.874717, 4.866093, 
    4.864969,
  // totalHeight(14,16, 0-49)
    5.003232, 4.974789, 4.948159, 4.924067, 4.903166, 4.886005, 4.872997, 
    4.864381, 4.860195, 4.860283, 4.864339, 4.872, 4.882958, 4.897115, 
    4.91473, 4.922801, 4.923217, 4.937708, 4.946001, 4.948301, 4.94475, 
    4.936777, 4.92233, 4.902053, 4.877351, 4.849022, 4.818892, 4.789238, 
    4.76301, 4.74164, 4.726334, 4.720396, 4.723143, 4.734078, 4.752094, 
    4.775647, 4.802935, 4.831992, 4.860762, 4.887154, 4.909132, 4.924897, 
    4.93313, 4.933318, 4.926054, 4.91317, 4.897569, 4.882729, 4.872013, 
    4.868022,
  // totalHeight(14,17, 0-49)
    4.995819, 4.967114, 4.940305, 4.916105, 4.895159, 4.878008, 4.865059, 
    4.856553, 4.85254, 4.852895, 4.857356, 4.865614, 4.877438, 4.892803, 
    4.912023, 4.929695, 4.934912, 4.951701, 4.962767, 4.967796, 4.966612, 
    4.959546, 4.945543, 4.924974, 4.899243, 4.869065, 4.836262, 4.803187, 
    4.773059, 4.747612, 4.728692, 4.718437, 4.717418, 4.725255, 4.740889, 
    4.762807, 4.789228, 4.818224, 4.84777, 4.875792, 4.900223, 4.919144, 
    4.930996, 4.934896, 4.930968, 4.920557, 4.906198, 4.891222, 4.879112, 
    4.872787,
  // totalHeight(14,18, 0-49)
    4.988537, 4.959641, 4.932666, 4.9083, 4.887167, 4.869789, 4.856569, 
    4.847752, 4.843416, 4.843479, 4.847744, 4.855983, 4.868048, 4.88397, 
    4.904027, 4.934335, 4.947203, 4.965634, 4.979208, 4.98692, 4.988139, 
    4.981914, 4.968329, 4.947478, 4.920774, 4.888891, 4.85365, 4.81746, 
    4.783762, 4.754593, 4.73253, 4.71814, 4.713455, 4.718208, 4.731387, 
    4.75151, 4.776821, 4.805424, 4.835332, 4.864502, 4.890868, 4.912439, 
    4.927494, 4.934857, 4.934252, 4.926565, 4.913923, 4.899424, 4.88655, 
    4.878451,
  // totalHeight(14,19, 0-49)
    4.981731, 4.952747, 4.925626, 4.901007, 4.879478, 4.86154, 4.847589, 
    4.837891, 4.832567, 4.831611, 4.834948, 4.842501, 4.854297, 4.870481, 
    4.891221, 4.936656, 4.959976, 4.979749, 4.995747, 5.00617, 5.009804, 
    5.004245, 4.990828, 4.969369, 4.941361, 4.907585, 4.869937, 4.830897, 
    4.794071, 4.761743, 4.73723, 4.719127, 4.711077, 4.712924, 4.723711, 
    4.741991, 4.766041, 4.793996, 4.823914, 4.853789, 4.881576, 4.90526, 
    4.923007, 4.933437, 4.93594, 4.930997, 4.920331, 4.906754, 4.893658, 
    4.88432,
  // totalHeight(14,20, 0-49)
    4.975356, 4.946013, 4.918895, 4.894783, 4.874384, 4.858284, 4.846906, 
    4.840438, 4.838765, 4.841401, 4.847481, 4.8558, 4.864954, 4.87357, 
    4.880587, 30, 4.989855, 4.995119, 5.000073, 5.003455, 5.004048, 4.997201, 
    4.985688, 4.96794, 4.944427, 4.914887, 4.880343, 4.842763, 4.805717, 
    4.771926, 4.745841, 4.724278, 4.712812, 4.711535, 4.719627, 4.735713, 
    4.758105, 4.784973, 4.814407, 4.844437, 4.873043, 4.898208, 4.918039, 
    4.931002, 4.936229, 4.933856, 4.92523, 4.912845, 4.899946, 4.889857,
  // totalHeight(14,21, 0-49)
    4.970289, 4.941153, 4.914182, 4.890114, 4.869606, 4.853193, 4.841239, 
    4.833877, 4.830952, 4.831978, 4.836136, 4.842323, 4.849247, 4.85558, 
    4.860119, 30, 5.006929, 5.011988, 5.017016, 5.020457, 5.020889, 5.011185, 
    4.997466, 4.977767, 4.952747, 4.922137, 4.886837, 4.848618, 4.81087, 
    4.776311, 4.749987, 4.726534, 4.71325, 4.710298, 4.716912, 4.731764, 
    4.753213, 4.779468, 4.808661, 4.838869, 4.868112, 4.894393, 4.915797, 
    4.930689, 4.938019, 4.937646, 4.930596, 4.919082, 4.906178, 4.895215,
  // totalHeight(14,22, 0-49)
    4.96617, 4.937153, 4.910255, 4.886184, 4.865558, 4.848874, 4.83646, 
    4.828418, 4.824572, 4.824438, 4.827231, 4.831902, 4.837212, 4.841824, 
    4.844385, 30, 5.018405, 5.023205, 5.02841, 5.032224, 5.033048, 5.021325, 
    5.00638, 4.985718, 4.960042, 4.928993, 4.893322, 4.85464, 4.816243, 
    4.780902, 4.754295, 4.728978, 4.713942, 4.709406, 4.71464, 4.728346, 
    4.748909, 4.774562, 4.803468, 4.833735, 4.863416, 4.890533, 4.913163, 
    4.929612, 4.938688, 4.940041, 4.934431, 4.923813, 4.911096, 4.899575,
  // totalHeight(14,23, 0-49)
    4.96328, 4.934348, 4.907502, 4.883425, 4.862714, 4.845841, 4.833112, 
    4.824607, 4.820145, 4.819244, 4.821142, 4.824821, 4.829068, 4.832527, 
    4.833734, 30, 5.025937, 5.030453, 5.035746, 5.039857, 5.041064, 5.027761, 
    5.011934, 4.990608, 4.964503, 4.9332, 4.897349, 4.85845, 4.819719, 
    4.783957, 4.757343, 4.730652, 4.714336, 4.708647, 4.712873, 4.725742, 
    4.745659, 4.770877, 4.799579, 4.829896, 4.859901, 4.887634, 4.911168, 
    4.928766, 4.939146, 4.941798, 4.937283, 4.927362, 4.914799, 4.902847,
  // totalHeight(14,24, 0-49)
    4.961791, 4.932945, 4.906162, 4.882113, 4.861383, 4.844429, 4.831546, 
    4.822805, 4.81802, 4.816717, 4.818145, 4.821302, 4.824994, 4.827858, 
    4.828371, 30, 5.029955, 5.034287, 5.039621, 5.043921, 5.045398, 5.031094, 
    5.014718, 4.992973, 4.966591, 4.935138, 4.899226, 4.8603, 4.821521, 
    4.785698, 4.759323, 4.731932, 4.714949, 4.708636, 4.712295, 4.724666, 
    4.744171, 4.76908, 4.797589, 4.827847, 4.857946, 4.88594, 4.909908, 
    4.928101, 4.939186, 4.942573, 4.93871, 4.929234, 4.916815, 4.904671,
  // totalHeight(14,25, 0-49)
    4.961771, 4.933026, 4.906334, 4.882361, 4.86169, 4.844777, 4.831912, 
    4.823165, 4.818351, 4.816997, 4.818359, 4.821449, 4.825079, 4.827899, 
    4.828384, 30, 5.03003, 5.034381, 5.039783, 5.044186, 5.045787, 5.031203, 
    5.014672, 4.992793, 4.966319, 4.934835, 4.89897, 4.860161, 4.821557, 
    4.785944, 4.759897, 4.732482, 4.715449, 4.709057, 4.712609, 4.724858, 
    4.744236, 4.769025, 4.797433, 4.827615, 4.857674, 4.88567, 4.909687, 
    4.927975, 4.939195, 4.942734, 4.939016, 4.929639, 4.917246, 4.905041,
  // totalHeight(14,26, 0-49)
    4.963167, 4.93454, 4.907962, 4.884112, 4.863579, 4.846827, 4.834151, 
    4.825628, 4.821076, 4.820027, 4.821736, 4.825215, 4.829287, 4.832619, 
    4.833757, 30, 5.026039, 5.030636, 5.036156, 5.040594, 5.042174, 5.028095, 
    5.011848, 4.990179, 4.963848, 4.932496, 4.896807, 4.858271, 4.820046, 
    4.784883, 4.759194, 4.73243, 4.715955, 4.710011, 4.713904, 4.726387, 
    4.745905, 4.770749, 4.799131, 4.829207, 4.85908, 4.886809, 4.91048, 
    4.928358, 4.939132, 4.942234, 4.938139, 4.928508, 4.91602, 4.903892,
  // totalHeight(14,27, 0-49)
    4.965813, 4.937301, 4.910845, 4.887145, 4.866809, 4.850321, 4.837995, 
    4.829924, 4.825934, 4.825562, 4.828056, 4.832419, 4.837465, 4.841897, 
    4.844372, 30, 5.018102, 5.023104, 5.028753, 5.033145, 5.034584, 5.021748, 
    5.006234, 4.985136, 4.959219, 4.928194, 4.892848, 4.854764, 4.817146, 
    4.782689, 4.757411, 4.731923, 4.71657, 4.711563, 4.716202, 4.729245, 
    4.749143, 4.774192, 4.802603, 4.832528, 4.862057, 4.88924, 4.912171, 
    4.929139, 4.938899, 4.940991, 4.93603, 4.925817, 4.913135, 4.901226,
  // totalHeight(14,28, 0-49)
    4.969423, 4.940984, 4.914621, 4.891065, 4.870954, 4.854809, 4.842978, 
    4.835584, 4.832475, 4.833191, 4.836968, 4.842775, 4.849395, 4.855551, 
    4.860049, 30, 5.006672, 5.0121, 5.017801, 5.022041, 5.023263, 5.01228, 
    4.997938, 4.977812, 4.952632, 4.922198, 4.887433, 4.850056, 4.81334, 
    4.779905, 4.755203, 4.731562, 4.717834, 4.714186, 4.719908, 4.733754, 
    4.754178, 4.779477, 4.80786, 4.837467, 4.866374, 4.892624, 4.914323, 
    4.929817, 4.937974, 4.938513, 4.932271, 4.921261, 4.908408, 4.896985,
  // totalHeight(14,29, 0-49)
    4.973598, 4.945132, 4.91878, 4.895313, 4.875417, 4.859663, 4.848455, 
    4.841969, 4.840096, 4.842386, 4.848045, 4.855969, 4.864852, 4.873392, 
    4.88053, 30, 4.991336, 4.997087, 5.002714, 5.006726, 5.007765, 4.999115, 
    4.986455, 4.96784, 4.943899, 4.91449, 4.880672, 4.844324, 4.808808, 
    4.776659, 4.752664, 4.731198, 4.719398, 4.717382, 4.724414, 4.739241, 
    4.760315, 4.785926, 4.81427, 4.84347, 4.871576, 4.896624, 4.916734, 
    4.930334, 4.936449, 4.935032, 4.927205, 4.915243, 4.902236, 4.891462,
  // totalHeight(14,30, 0-49)
    4.978459, 4.950448, 4.924171, 4.90026, 4.879285, 4.861737, 4.848003, 
    4.838342, 4.832888, 4.831677, 4.83469, 4.841944, 4.853562, 4.869802, 
    4.890952, 4.937116, 4.960141, 4.981357, 4.999086, 5.011297, 5.016665, 
    5.010939, 4.99806, 4.977265, 4.949973, 4.916874, 4.879813, 4.841241, 
    4.804756, 4.772696, 4.748902, 4.729621, 4.719982, 4.719895, 4.728523, 
    4.744562, 4.766439, 4.792431, 4.820715, 4.84939, 4.876489, 4.900041, 
    4.918213, 4.929551, 4.93329, 4.929682, 4.920183, 4.907356, 4.894434, 
    4.88467,
  // totalHeight(14,31, 0-49)
    4.983125, 4.955338, 4.929348, 4.905835, 4.885411, 4.868597, 4.85578, 
    4.847207, 4.842966, 4.843014, 4.847225, 4.855464, 4.867691, 4.884041, 
    4.904872, 4.935839, 4.949141, 4.969279, 4.984799, 4.994443, 4.997485, 
    4.991339, 4.978379, 4.958244, 4.932343, 4.901263, 4.86675, 4.83112, 
    4.797772, 4.768725, 4.747015, 4.731064, 4.72435, 4.726704, 4.737257, 
    4.754694, 4.777433, 4.803735, 4.831755, 4.85956, 4.885167, 4.906618, 
    4.922161, 4.930507, 4.931175, 4.92478, 4.913159, 4.899173, 4.886178, 
    4.877337,
  // totalHeight(14,32, 0-49)
    4.987358, 4.959856, 4.934148, 4.91095, 4.890905, 4.874556, 4.862307, 
    4.854393, 4.850876, 4.851655, 4.85653, 4.865274, 4.877754, 4.894031, 
    4.914469, 4.932961, 4.939357, 4.958105, 4.971329, 4.978452, 4.979202, 
    4.972534, 4.959299, 4.939528, 4.914677, 4.885373, 4.853353, 4.820845, 
    4.790998, 4.765457, 4.746442, 4.73423, 4.730731, 4.735687, 4.748199, 
    4.766947, 4.790341, 4.816634, 4.843962, 4.870373, 4.893885, 4.912594, 
    4.924883, 4.929708, 4.926944, 4.917631, 4.904008, 4.889196, 4.876601, 
    4.869208,
  // totalHeight(14,33, 0-49)
    4.99063, 4.963439, 4.938015, 4.915095, 4.895347, 4.879332, 4.867464, 
    4.859974, 4.856893, 4.858074, 4.863241, 4.872085, 4.88437, 4.900063, 
    4.919447, 4.928698, 4.931004, 4.947732, 4.958413, 4.962972, 4.961474, 
    4.954248, 4.940749, 4.921361, 4.897592, 4.870147, 4.840767, 4.811585, 
    4.785475, 4.763719, 4.747799, 4.739508, 4.739332, 4.746913, 4.761318, 
    4.78121, 4.804995, 4.83091, 4.85707, 4.88152, 4.902306, 4.917626, 
    4.926063, 4.926908, 4.920468, 4.908258, 4.892908, 4.877741, 4.866107, 
    4.860717,
  // totalHeight(14,34, 0-49)
    4.992525, 4.96564, 4.940499, 4.917854, 4.898386, 4.882666, 4.871113, 
    4.863943, 4.86116, 4.862561, 4.867793, 4.876443, 4.888147, 4.902713, 
    4.920231, 4.923387, 4.923928, 4.937998, 4.945892, 4.947875, 4.944241, 
    4.936496, 4.92287, 4.90407, 4.881607, 4.856267, 4.829761, 4.804101, 
    4.781861, 4.764022, 4.751439, 4.747082, 4.750193, 4.760307, 4.776446, 
    4.797251, 4.821106, 4.846224, 4.870707, 4.892605, 4.910032, 4.921345, 
    4.92542, 4.921961, 4.911783, 4.896895, 4.880278, 4.865354, 4.855299, 
    4.852454,
  // totalHeight(14,35, 0-49)
    4.99278, 4.96617, 4.941314, 4.91896, 4.899793, 4.884388, 4.873153, 
    4.866287, 4.863753, 4.865289, 4.87046, 4.87873, 4.889587, 4.902627, 
    4.917654, 4.917314, 4.917788, 4.928729, 4.933709, 4.933207, 4.927653, 
    4.919489, 4.905965, 4.888046, 4.867195, 4.844253, 4.820849, 4.798853, 
    4.780519, 4.766601, 4.757459, 4.756906, 4.763144, 4.775598, 4.793231, 
    4.814648, 4.838199, 4.862067, 4.884343, 4.903111, 4.916597, 4.923395, 
    4.922756, 4.914888, 4.901155, 4.884047, 4.866805, 4.85282, 4.844973, 
    4.84515,
  // totalHeight(14,36, 0-49)
    4.991346, 4.964972, 4.940395, 4.918357, 4.899533, 4.884483, 4.873598, 
    4.867045, 4.864746, 4.866374, 4.871405, 4.879189, 4.889049, 4.900362, 
    4.912611, 4.910634, 4.912133, 4.919724, 4.921842, 4.919075, 4.911914, 
    4.903495, 4.890347, 4.873635, 4.854704, 4.834425, 4.814302, 4.79603, 
    4.781533, 4.77143, 4.765703, 4.768709, 4.777803, 4.792308, 4.811116, 
    4.832782, 4.855612, 4.877761, 4.897319, 4.912441, 4.921529, 4.923491, 
    4.918043, 4.905955, 4.889152, 4.870528, 4.853456, 4.841154, 4.836089, 
    4.839647,
  // totalHeight(14,37, 0-49)
    4.988453, 4.962273, 4.937971, 4.916267, 4.897817, 4.883152, 4.872628, 
    4.866377, 4.864271, 4.865924, 4.870734, 4.877946, 4.88674, 4.896296, 
    4.905811, 4.903345, 4.906444, 4.910737, 4.910229, 4.90555, 4.897175, 
    4.888714, 4.876239, 4.86105, 4.844311, 4.826896, 4.810146, 4.795563, 
    4.784745, 4.778251, 4.77579, 4.782004, 4.793592, 4.809768, 4.829356, 
    4.850853, 4.87252, 4.892492, 4.908888, 4.919978, 4.924416, 4.921508, 
    4.911499, 4.895743, 4.87667, 4.857455, 4.841446, 4.831538, 4.829711, 
    4.836845,
  // totalHeight(14,38, 0-49)
    4.984639, 4.958626, 4.934591, 4.913228, 4.895154, 4.880854, 4.870646, 
    4.86461, 4.862578, 4.864117, 4.868563, 4.875087, 4.882763, 4.890626, 
    4.897676, 4.89531, 4.900163, 4.901466, 4.898746, 4.892606, 4.88346, 
    4.875215, 4.863713, 4.850336, 4.836003, 4.821574, 4.808197, 4.797181, 
    4.789793, 4.786611, 4.787156, 4.796136, 4.809761, 4.82715, 4.84706, 
    4.867931, 4.887993, 4.905383, 4.918293, 4.92518, 4.925019, 4.917578, 
    4.903661, 4.885168, 4.864916, 4.846192, 4.832146, 4.825239, 4.826932, 
    4.837641,
  // totalHeight(14,39, 0-49)
    4.980752, 4.95491, 4.931138, 4.910096, 4.892348, 4.878327, 4.868291, 
    4.862281, 4.86009, 4.861258, 4.865097, 4.870739, 4.877207, 4.88346, 
    4.888396, 4.886341, 4.892785, 4.891613, 4.887215, 4.88012, 4.87067, 
    4.862928, 4.852697, 4.841382, 4.829606, 4.818201, 4.808114, 4.800452, 
    4.796173, 4.795929, 4.799117, 4.810341, 4.825474, 4.843554, 4.863278, 
    4.883053, 4.901103, 4.915614, 4.924913, 4.927712, 4.92337, 4.912158, 
    4.895406, 4.875451, 4.855321, 4.838219, 4.826949, 4.82348, 4.828774, 
    4.842854,
  // totalHeight(14,40, 0-49)
    4.977879, 4.952263, 4.928766, 4.908001, 4.890475, 4.876557, 4.866449, 
    4.860152, 4.857441, 4.857857, 4.860724, 4.86519, 4.87028, 4.874952, 
    4.878095, 4.876329, 4.883979, 4.880965, 4.875467, 4.867936, 4.858642, 
    4.851704, 4.843017, 4.833961, 4.824832, 4.816414, 4.809454, 4.804865, 
    4.80331, 4.805566, 4.810947, 4.823834, 4.839893, 4.8581, 4.87712, 
    4.895356, 4.911077, 4.92258, 4.928399, 4.927567, 4.919873, 4.906066, 
    4.88791, 4.868001, 4.849374, 4.834966, 4.827127, 4.827327, 4.836097, 
    4.853168,
  // totalHeight(14,41, 0-49)
    4.977243, 4.951975, 4.928784, 4.908237, 4.890777, 4.876709, 4.866188, 
    4.859186, 4.855484, 4.854657, 4.856086, 4.858981, 4.862435, 4.865462, 
    4.867022, 4.865379, 4.873715, 4.869505, 4.863459, 4.855964, 4.84724, 
    4.841386, 4.834473, 4.827814, 4.821355, 4.81582, 4.811758, 4.8099, 
    4.810643, 4.814913, 4.82198, 4.835919, 4.852301, 4.870073, 4.8879, 
    4.904237, 4.91746, 4.92605, 4.928823, 4.925181, 4.915336, 4.900439, 
    4.882529, 4.864255, 4.848449, 4.837637, 4.833674, 4.837571, 4.849523, 
    4.869064,
  // totalHeight(14,42, 0-49)
    4.980048, 4.955317, 4.932497, 4.912102, 4.894521, 4.880002, 4.868662, 
    4.860474, 4.855247, 4.852629, 4.852093, 4.852965, 4.854447, 4.855668, 
    4.855711, 4.853931, 4.862373, 4.857519, 4.851374, 4.844295, 4.836475, 
    4.831925, 4.826941, 4.822737, 4.818897, 4.816074, 4.814629, 4.815122, 
    4.817711, 4.823489, 4.831711, 4.846095, 4.862226, 4.879052, 4.895293, 
    4.909513, 4.92027, 4.926304, 4.926771, 4.921447, 4.910919, 4.896608, 
    4.88063, 4.865476, 4.85361, 4.847065, 4.847208, 4.854662, 4.869378, 
    4.89079,
  // totalHeight(14,43, 0-49)
    4.987293, 4.963366, 4.941016, 4.920723, 4.902826, 4.887541, 4.874972, 
    4.865113, 4.857836, 4.852889, 4.849873, 4.848258, 4.847405, 4.846586, 
    4.845038, 4.842797, 4.850761, 4.845643, 4.839696, 4.833277, 4.826568, 
    4.82345, 4.820451, 4.818665, 4.817314, 4.816969, 4.817812, 4.820253, 
    4.824242, 4.831039, 4.839899, 4.854184, 4.869569, 4.885051, 4.89946, 
    4.911537, 4.920093, 4.924184, 4.923324, 4.917646, 4.908003, 4.895916, 
    4.88339, 4.872587, 4.865491, 4.863626, 4.867915, 4.878666, 4.895671, 
    4.918324,
  // totalHeight(14,44, 0-49)
    4.999643, 4.97684, 4.955107, 4.934894, 4.916515, 4.900183, 4.886018, 
    4.874065, 4.864291, 4.85656, 4.850628, 4.846134, 4.842605, 4.839487, 
    4.83618, 4.833108, 4.840065, 4.83484, 4.82921, 4.823539, 4.818005, 
    4.81632, 4.815243, 4.815725, 4.816647, 4.818492, 4.821272, 4.825261, 
    4.830235, 4.837609, 4.846658, 4.8604, 4.874674, 4.888574, 4.901094, 
    4.911215, 4.918052, 4.921008, 4.91994, 4.915264, 4.907966, 4.899511, 
    4.891633, 4.886055, 4.884239, 4.887223, 4.895544, 4.909267, 4.928077, 
    4.951357,
  // totalHeight(14,45, 0-49)
    5.017312, 4.996, 4.97507, 4.95496, 4.935992, 4.918405, 4.902376, 4.88803, 
    4.875444, 4.864624, 4.855481, 4.847826, 4.841365, 4.835716, 4.83044, 
    4.826169, 4.831665, 4.826299, 4.820926, 4.815934, 4.811489, 4.81111, 
    4.811764, 4.814254, 4.81716, 4.820862, 4.825219, 4.830384, 4.835991, 
    4.843586, 4.852475, 4.865373, 4.878339, 4.890605, 4.901376, 4.909918, 
    4.915675, 4.918389, 4.918215, 4.915745, 4.911979, 4.908191, 4.905741, 
    4.90587, 4.909535, 4.917328, 4.92946, 4.945801, 4.965949, 4.989285,
  // totalHeight(14,46, 0-49)
    5.040022, 5.0206, 5.000702, 4.98078, 4.9612, 4.942265, 4.924236, 
    4.907354, 4.891817, 4.877773, 4.865296, 4.854357, 4.84483, 4.83649, 
    4.829052, 4.823248, 4.82694, 4.821243, 4.81594, 4.811431, 4.807864, 
    4.808546, 4.810627, 4.814773, 4.819308, 4.82451, 4.8301, 4.836121, 
    4.842098, 4.849669, 4.858179, 4.870093, 4.881728, 4.892483, 4.901812, 
    4.909278, 4.914648, 4.917972, 4.919623, 4.920277, 4.920839, 4.922309, 
    4.92564, 4.931595, 4.94067, 4.953065, 4.968709, 4.987298, 5.008345, 
    5.031216,
  // totalHeight(14,47, 0-49)
    5.067022, 5.049904, 5.031317, 5.011751, 4.991643, 4.971396, 4.951393, 
    4.931998, 4.913552, 4.896341, 4.880581, 4.866395, 4.853802, 4.842718, 
    4.832986, 4.825392, 4.827056, 4.820758, 4.815261, 4.810961, 4.807976, 
    4.809393, 4.812525, 4.817905, 4.823682, 4.830026, 4.836539, 4.843167, 
    4.849349, 4.856772, 4.86482, 4.875768, 4.8862, 4.89571, 4.904, 4.910928, 
    4.916553, 4.921173, 4.925306, 4.929629, 4.934891, 4.941786, 4.950864, 
    4.962459, 4.976653, 4.993308, 5.012097, 5.032546, 5.05407, 5.075994,
  // totalHeight(14,48, 0-49)
    5.097138, 5.082759, 5.065822, 5.046871, 5.026447, 5.005077, 4.983285, 
    4.961578, 4.940433, 4.920274, 4.901444, 4.884194, 4.868665, 4.854891, 
    4.842824, 4.833281, 4.832807, 4.825633, 4.819666, 4.81528, 4.812549, 
    4.814342, 4.818109, 4.824279, 4.830903, 4.838052, 4.845232, 4.852296, 
    4.858621, 4.86589, 4.873518, 4.883643, 4.893113, 4.901714, 4.90939, 
    4.916262, 4.922637, 4.928999, 4.935947, 4.944109, 4.954046, 4.966163, 
    4.980648, 4.997454, 5.016309, 5.036768, 5.058268, 5.080154, 5.101726, 
    5.122242,
  // totalHeight(14,49, 0-49)
    5.131782, 5.121768, 5.107812, 5.090503, 5.070491, 5.048445, 5.025044, 
    5.000954, 4.976798, 4.953141, 4.93047, 4.909184, 4.889575, 4.87183, 
    4.856054, 4.844022, 4.848143, 4.838534, 4.83033, 4.824347, 4.820787, 
    4.825149, 4.832235, 4.842608, 4.852149, 4.861037, 4.868387, 4.874065, 
    4.877024, 4.881012, 4.885324, 4.894529, 4.902976, 4.910685, 4.917894, 
    4.925021, 4.93263, 4.941376, 4.951897, 4.964715, 4.980152, 4.99826, 
    5.018826, 5.04138, 5.065258, 5.08966, 5.113735, 5.1366, 5.15739, 5.175267,
  // totalHeight(15,0, 0-49)
    5.116331, 5.087602, 5.057508, 5.02688, 4.99647, 4.966957, 4.938937, 
    4.912934, 4.889373, 4.86856, 4.850661, 4.835689, 4.823497, 4.813806, 
    4.806232, 4.800476, 4.797285, 4.793497, 4.79044, 4.787902, 4.785748, 
    4.784293, 4.783263, 4.78291, 4.783345, 4.784853, 4.787655, 4.791958, 
    4.797826, 4.805394, 4.814459, 4.825126, 4.83667, 4.848646, 4.860583, 
    4.872067, 4.882796, 4.892663, 4.901782, 4.910505, 4.919398, 4.929152, 
    4.940503, 4.954107, 4.970463, 4.989839, 5.012252, 5.037459, 5.064975, 
    5.094105,
  // totalHeight(15,1, 0-49)
    5.096625, 5.067094, 5.036662, 5.006133, 4.976219, 4.94755, 4.920673, 
    4.896048, 4.874031, 4.854852, 4.838602, 4.825209, 4.81445, 4.805967, 
    4.799304, 4.794245, 4.792803, 4.788857, 4.785463, 4.782435, 4.779634, 
    4.777761, 4.776192, 4.775315, 4.77516, 4.776093, 4.778361, 4.782217, 
    4.787709, 4.795141, 4.804237, 4.815469, 4.827672, 4.840302, 4.852779, 
    4.864544, 4.87516, 4.884389, 4.892262, 4.899111, 4.905552, 4.912408, 
    4.920602, 4.931015, 4.944372, 4.961137, 4.981477, 5.005255, 5.032047, 
    5.061183,
  // totalHeight(15,2, 0-49)
    5.078791, 5.048922, 5.018562, 4.988491, 4.95939, 4.931859, 4.906399, 
    4.883417, 4.863198, 4.845896, 4.831511, 4.819883, 4.810696, 4.803508, 
    4.797784, 4.793371, 4.793595, 4.789402, 4.78556, 4.781904, 4.778296, 
    4.775818, 4.773477, 4.771796, 4.770742, 4.770769, 4.772155, 4.775218, 
    4.780015, 4.787013, 4.795884, 4.807501, 4.820284, 4.833621, 4.846819, 
    4.859183, 4.870113, 4.879212, 4.886373, 4.891838, 4.89621, 4.900389, 
    4.905457, 4.912516, 4.922533, 4.936205, 4.953891, 4.975585, 5.000948, 
    5.029352,
  // totalHeight(15,3, 0-49)
    5.06324, 5.033447, 5.003518, 4.974208, 4.946181, 4.920012, 4.896168, 
    4.875008, 4.856752, 4.841472, 4.829074, 4.819304, 4.811752, 4.805884, 
    4.801088, 4.797221, 4.798965, 4.794469, 4.790111, 4.78574, 4.781212, 
    4.777983, 4.774674, 4.771935, 4.769695, 4.768483, 4.768632, 4.770534, 
    4.774281, 4.780493, 4.788819, 4.800562, 4.81377, 4.827785, 4.841828, 
    4.855076, 4.866765, 4.876311, 4.883421, 4.888182, 4.891104, 4.893085, 
    4.895307, 4.899062, 4.905564, 4.915772, 4.93028, 4.949261, 4.972499, 
    4.999438,
  // totalHeight(15,4, 0-49)
    5.050073, 5.020701, 4.9915, 4.963202, 4.936454, 4.911811, 4.889717, 
    4.87048, 4.854262, 4.841056, 4.830678, 4.822776, 4.81685, 4.812282, 
    4.808378, 4.804924, 4.807982, 4.803201, 4.798327, 4.79323, 4.787751, 
    4.783697, 4.779289, 4.77529, 4.771614, 4.768863, 4.767426, 4.767785, 
    4.770104, 4.775139, 4.782532, 4.794057, 4.807438, 4.822003, 4.836916, 
    4.851248, 4.864085, 4.874649, 4.88243, 4.887299, 4.88959, 4.890103, 
    4.890029, 4.890785, 4.89381, 4.900341, 4.911246, 4.92694, 4.947388, 
    4.972149,
  // totalHeight(15,5, 0-49)
    5.039103, 5.010417, 4.982175, 4.95508, 4.929761, 4.906757, 4.886483, 
    4.869208, 4.855032, 4.843874, 4.835467, 4.829376, 4.825019, 4.821709, 
    4.818674, 4.815492, 4.819603, 4.814657, 4.809369, 4.803624, 4.797256, 
    4.792387, 4.786834, 4.781446, 4.776152, 4.771607, 4.768267, 4.766716, 
    4.767217, 4.770647, 4.77667, 4.787555, 4.800759, 4.81563, 4.831312, 
    4.846801, 4.861059, 4.873127, 4.882268, 4.888099, 4.8907, 4.89067, 
    4.889099, 4.887434, 4.887277, 4.890124, 4.89716, 4.909099, 4.926156, 
    4.948071,
  // totalHeight(15,6, 0-49)
    5.029912, 5.00209, 4.974963, 4.949202, 4.925413, 4.904112, 4.885684, 
    4.870354, 4.85817, 4.848981, 4.84245, 4.838074, 4.835212, 4.833121, 
    4.830979, 4.827941, 4.832795, 4.827935, 4.822438, 4.816226, 4.809129, 
    4.803551, 4.796894, 4.790074, 4.783056, 4.776528, 4.771018, 4.767218, 
    4.765527, 4.766914, 4.771096, 4.780854, 4.793445, 4.80827, 4.824483, 
    4.841054, 4.856845, 4.870752, 4.88182, 4.889394, 4.893252, 4.893704, 
    4.891622, 4.888361, 4.885583, 4.885003, 4.888118, 4.895999, 4.909183, 
    4.927671,
  // totalHeight(15,7, 0-49)
    5.021935, 4.99507, 4.96914, 4.944782, 4.922575, 4.902999, 4.886406, 
    4.872977, 4.862704, 4.855379, 4.850611, 4.847847, 4.846417, 4.845552, 
    4.844402, 4.841412, 4.846661, 4.84226, 4.836864, 4.83046, 4.822882, 
    4.816778, 4.809143, 4.800937, 4.792175, 4.783555, 4.775673, 4.769339, 
    4.765112, 4.764037, 4.765896, 4.774005, 4.785484, 4.799817, 4.816212, 
    4.833632, 4.850895, 4.866778, 4.880141, 4.89007, 4.896023, 4.897958, 
    4.896429, 4.892569, 4.887981, 4.884502, 4.88391, 4.887653, 4.896658, 
    4.911267,
  // totalHeight(15,8, 0-49)
    5.014567, 4.988669, 4.963949, 4.941008, 4.920386, 4.902526, 4.887734, 
    4.876143, 4.867693, 4.862128, 4.859016, 4.857789, 4.857767, 4.858192, 
    4.858227, 4.855232, 4.860509, 4.857036, 4.852131, 4.845875, 4.838133, 
    4.83175, 4.82334, 4.813871, 4.803432, 4.792694, 4.782328, 4.773249, 
    4.766201, 4.762278, 4.76136, 4.767284, 4.777114, 4.790453, 4.806582, 
    4.824496, 4.842996, 4.860787, 4.876583, 4.889243, 4.897914, 4.902189, 
    4.902226, 4.898835, 4.893422, 4.887823, 4.884019, 4.883815, 4.888562, 
    4.899018,
  // totalHeight(15,9, 0-49)
    5.007263, 4.982272, 4.958714, 4.937149, 4.918076, 4.901892, 4.888849, 
    4.879029, 4.872319, 4.868426, 4.866897, 4.867163, 4.868573, 4.870416, 
    4.871912, 4.868925, 4.873866, 4.87183, 4.867853, 4.862131, 4.854586, 
    4.848204, 4.83927, 4.828737, 4.816766, 4.803984, 4.791113, 4.779171, 
    4.76909, 4.762001, 4.7579, 4.761126, 4.768773, 4.780583, 4.795938, 
    4.813896, 4.833264, 4.85271, 4.870847, 4.886352, 4.898101, 4.905329, 
    4.907785, 4.905872, 4.900687, 4.893928, 4.887661, 4.883976, 4.884649, 
    4.890883,
  // totalHeight(15,10, 0-49)
    4.999604, 4.975416, 4.952922, 4.932649, 4.915052, 4.900475, 4.889113, 
    4.880991, 4.875949, 4.873662, 4.873672, 4.875424, 4.878328, 4.881759, 
    4.885052, 4.882169, 4.886457, 4.886337, 4.883721, 4.878932, 4.87196, 
    4.865866, 4.856699, 4.845355, 4.832079, 4.817416, 4.802129, 4.787311, 
    4.774088, 4.7636, 4.755988, 4.756044, 4.760993, 4.770745, 4.784802, 
    4.802295, 4.822069, 4.84278, 4.862974, 4.881195, 4.896103, 4.906617, 
    4.912094, 4.912504, 4.908549, 4.901665, 4.893864, 4.887411, 4.884446, 
    4.886625,
  // totalHeight(15,11, 0-49)
    4.991342, 4.967822, 4.946262, 4.927166, 4.910937, 4.897869, 4.8881, 
    4.881597, 4.878156, 4.877424, 4.878942, 4.882198, 4.886673, 4.891865, 
    4.897288, 4.89474, 4.898158, 4.900331, 4.899464, 4.895978, 4.889944, 
    4.88441, 4.875308, 4.863452, 4.849164, 4.832879, 4.815373, 4.797784, 
    4.781417, 4.767402, 4.756055, 4.752538, 4.754327, 4.761522, 4.773763, 
    4.790272, 4.809944, 4.831436, 4.853266, 4.873887, 4.891792, 4.905651, 
    4.914472, 4.917807, 4.915928, 4.909914, 4.901585, 4.893248, 4.8873, 
    4.885808,
  // totalHeight(15,12, 0-49)
    4.982402, 4.959404, 4.938636, 4.920569, 4.905574, 4.893891, 4.885602, 
    4.880623, 4.878705, 4.879471, 4.882472, 4.887239, 4.893341, 4.900425, 
    4.908225, 4.906451, 4.908953, 4.913633, 4.914804, 4.91294, 4.908176, 
    4.903432, 4.894686, 4.88264, 4.867683, 4.850114, 4.830691, 4.810552, 
    4.791155, 4.773605, 4.758424, 4.751015, 4.749251, 4.753448, 4.763399, 
    4.778428, 4.797483, 4.819242, 4.842208, 4.86478, 4.885344, 4.90237, 
    4.914593, 4.92119, 4.922007, 4.917713, 4.90983, 4.900563, 4.892437, 
    4.887838,
  // totalHeight(15,13, 0-49)
    4.972854, 4.950241, 4.930109, 4.912913, 4.898992, 4.888544, 4.881598, 
    4.87802, 4.877524, 4.879713, 4.884143, 4.890391, 4.89812, 4.907125, 
    4.917382, 4.917123, 4.918903, 4.926107, 4.929477, 4.929471, 4.926257, 
    4.922477, 4.914348, 4.90243, 4.887171, 4.868714, 4.847758, 4.825398, 
    4.803198, 4.782228, 4.763248, 4.751732, 4.746114, 4.746946, 4.7542, 
    4.767303, 4.785262, 4.806781, 4.830365, 4.854382, 4.877144, 4.897, 
    4.912463, 4.922406, 4.926286, 4.924352, 4.917756, 4.908478, 4.899033, 
    4.892014,
  // totalHeight(15,14, 0-49)
    4.96287, 4.940514, 4.920871, 4.904384, 4.891365, 4.881975, 4.876204, 
    4.873875, 4.874665, 4.878159, 4.883919, 4.89156, 4.900823, 4.911641, 
    4.924194, 4.926576, 4.928138, 4.937673, 4.943261, 4.945259, 4.943804, 
    4.941094, 4.933791, 4.922291, 4.907089, 4.888156, 4.866101, 4.841918, 
    4.817236, 4.793077, 4.770475, 4.754752, 4.745088, 4.742292, 4.746523, 
    4.757329, 4.773777, 4.7946, 4.818307, 4.843254, 4.867715, 4.889956, 
    4.908341, 4.921505, 4.928574, 4.929399, 4.924733, 4.916243, 4.906309, 
    4.897605,
  // totalHeight(15,15, 0-49)
    4.952686, 4.930484, 4.911194, 4.895252, 4.88295, 4.874424, 4.869629, 
    4.868354, 4.870248, 4.874878, 4.881808, 4.890677, 4.901279, 4.913642, 
    4.92807, 4.93463, 4.936832, 4.948342, 4.95604, 4.960089, 4.960528, 
    4.958922, 4.952585, 4.941731, 4.926888, 4.907864, 4.885134, 4.85956, 
    4.832775, 4.80575, 4.779841, 4.759933, 4.746149, 4.739574, 4.740567, 
    4.748801, 4.763408, 4.783151, 4.806544, 4.831944, 4.857608, 4.881755, 
    4.90265, 4.918758, 4.928937, 4.932689, 4.930367, 4.923283, 4.913586, 
    4.903914,
  // totalHeight(15,16, 0-49)
    4.942564, 4.920435, 4.90138, 4.885822, 4.874048, 4.866168, 4.862118, 
    4.86166, 4.864422, 4.869958, 4.877826, 4.887679, 4.899335, 4.912846, 
    4.92854, 4.941131, 4.945195, 4.958213, 4.967833, 4.973904, 4.976303, 
    4.975766, 4.970457, 4.960384, 4.946107, 4.927279, 4.904236, 4.877665, 
    4.849168, 4.819665, 4.790876, 4.766929, 4.749082, 4.738706, 4.736363, 
    4.741861, 4.7544, 4.77277, 4.795497, 4.820938, 4.847348, 4.872924, 
    4.89588, 4.91456, 4.92762, 4.934264, 4.934485, 4.929224, 4.920336, 
    4.910336,
  // totalHeight(15,17, 0-49)
    4.932777, 4.910663, 4.891735, 4.876411, 4.864961, 4.857486, 4.853906, 
    4.853971, 4.857299, 4.863437, 4.871946, 4.88248, 4.894852, 4.909085, 
    4.925418, 4.945959, 4.953385, 4.967457, 4.978798, 4.986842, 4.991218, 
    4.991667, 4.987359, 4.978087, 4.964433, 4.945938, 4.922795, 4.895525, 
    4.865663, 4.834091, 4.80294, 4.77522, 4.753508, 4.739446, 4.733802, 
    4.736515, 4.746866, 4.76367, 4.785466, 4.810616, 4.837379, 4.863954, 
    4.888523, 4.909357, 4.924963, 4.934315, 4.937086, 4.933866, 4.926193, 
    4.916392,
  // totalHeight(15,18, 0-49)
    4.923589, 4.901454, 4.882562, 4.867312, 4.855964, 4.848607, 4.845161, 
    4.845378, 4.848886, 4.855247, 4.864042, 4.874938, 4.887739, 4.902402, 
    4.918972, 4.949069, 4.961415, 4.976269, 4.989225, 4.999232, 5.005604, 
    5.006928, 5.003522, 4.994929, 4.981759, 4.963496, 4.940249, 4.9124, 
    4.881422, 4.848179, 4.815248, 4.784146, 4.758912, 4.741425, 4.732646, 
    4.732654, 4.740804, 4.755947, 4.776639, 4.801248, 4.828047, 4.855239, 
    4.881002, 4.903563, 4.921335, 4.933104, 4.938289, 4.93716, 4.930946, 
    4.921741,
  // totalHeight(15,19, 0-49)
    4.915263, 4.893085, 4.874133, 4.858778, 4.847258, 4.839663, 4.83592, 
    4.835809, 4.838999, 4.845114, 4.853805, 4.864809, 4.877959, 4.89312, 
    4.910018, 4.950513, 4.968981, 4.984726, 4.999439, 5.011564, 5.02004, 
    5.022157, 5.019508, 5.011316, 4.998226, 4.979774, 4.956087, 4.927523, 
    4.895533, 4.860983, 4.826902, 4.792949, 4.764691, 4.744195, 4.732588, 
    4.730083, 4.736119, 4.749599, 4.769093, 4.792991, 4.819576, 4.847066, 
    4.873648, 4.897533, 4.917068, 4.93091, 4.938273, 4.939157, 4.934505, 
    4.926172,
  // totalHeight(15,20, 0-49)
    4.908185, 4.886056, 4.867468, 4.852916, 4.84274, 4.837077, 4.835821, 
    4.838592, 4.844738, 4.853366, 4.863411, 4.873747, 4.883327, 4.89133, 
    4.897302, 30, 4.994577, 4.999668, 5.005548, 5.011305, 5.016126, 5.015633, 
    5.013115, 5.006968, 4.997258, 4.982792, 4.962961, 4.937488, 4.907465, 
    4.873701, 4.839848, 4.803802, 4.772908, 4.749545, 4.735105, 4.72999, 
    4.733762, 4.745383, 4.763453, 4.786373, 4.812434, 4.839869, 4.866875, 
    4.891658, 4.912527, 4.928051, 4.937283, 4.939999, 4.936891, 4.929584,
  // totalHeight(15,21, 0-49)
    4.90235, 4.880386, 4.861916, 4.847402, 4.837146, 4.831253, 4.829581, 
    4.831733, 4.837054, 4.844685, 4.853627, 4.862837, 4.871323, 4.878238, 
    4.882979, 30, 5.004196, 5.009486, 5.015777, 5.021951, 5.027033, 5.024549, 
    5.020569, 5.013208, 5.002763, 4.988084, 4.968498, 4.943565, 4.914167, 
    4.880956, 4.847917, 4.810899, 4.778774, 4.753971, 4.737977, 4.73131, 
    4.733636, 4.743992, 4.761029, 4.783178, 4.80876, 4.836029, 4.863201, 
    4.888492, 4.910194, 4.926821, 4.937312, 4.941274, 4.939192, 4.932497,
  // totalHeight(15,22, 0-49)
    4.897773, 4.875886, 4.857458, 4.842922, 4.832562, 4.826463, 4.824469, 
    4.826171, 4.830924, 4.837883, 4.846084, 4.854511, 4.862186, 4.868207, 
    4.871812, 30, 5.010537, 5.015932, 5.022656, 5.029411, 5.035066, 5.0311, 
    5.026239, 5.01824, 5.007516, 4.992895, 4.973616, 4.949099, 4.920087, 
    4.887161, 4.854692, 4.816629, 4.78334, 4.757275, 4.739974, 4.732033, 
    4.73318, 4.742507, 4.758702, 4.78022, 4.805398, 4.83251, 4.859784, 
    4.885447, 4.907785, 4.925273, 4.936773, 4.941762, 4.940569, 4.934464,
  // totalHeight(15,23, 0-49)
    4.894632, 4.872791, 4.854372, 4.839801, 4.829348, 4.823086, 4.820855, 
    4.822244, 4.826617, 4.833141, 4.840868, 4.848798, 4.855937, 4.861334, 
    4.864092, 30, 5.014832, 5.020237, 5.02725, 5.034447, 5.040577, 5.035399, 
    5.029847, 5.021343, 5.010375, 4.995757, 4.976672, 4.952449, 4.923741, 
    4.891075, 4.859142, 4.82031, 4.786209, 4.75929, 4.741114, 4.732311, 
    4.73266, 4.741292, 4.75692, 4.778018, 4.802937, 4.829955, 4.857316, 
    4.883248, 4.906034, 4.924124, 4.93632, 4.94202, 4.941433, 4.935718,
  // totalHeight(15,24, 0-49)
    4.89303, 4.871227, 4.852822, 4.83823, 4.827715, 4.821345, 4.818963, 
    4.820161, 4.824309, 4.830588, 4.838061, 4.845731, 4.8526, 4.857682, 4.86, 
    30, 5.017446, 5.022851, 5.03004, 5.037525, 5.043984, 5.038036, 5.032043, 
    5.023195, 5.012022, 4.997339, 4.978312, 4.954233, 4.925709, 4.893244, 
    4.861749, 4.822506, 4.787988, 4.760626, 4.741983, 4.732702, 4.732585, 
    4.740788, 4.756044, 4.776845, 4.801548, 4.828448, 4.855792, 4.881816, 
    4.904807, 4.9232, 4.935774, 4.941876, 4.941653, 4.936192,
  // totalHeight(15,25, 0-49)
    4.892978, 4.871228, 4.852853, 4.838268, 4.827735, 4.821324, 4.818879, 
    4.820003, 4.824073, 4.830282, 4.8377, 4.84534, 4.852205, 4.857303, 
    4.859646, 30, 5.017977, 5.023447, 5.030755, 5.038391, 5.045011, 5.03886, 
    5.032743, 5.023767, 5.012475, 4.997696, 4.978612, 4.954521, 4.926036, 
    4.893661, 4.862384, 4.823091, 4.788538, 4.761134, 4.742421, 4.733041, 
    4.732802, 4.74087, 4.755989, 4.776659, 4.801252, 4.828063, 4.855346, 
    4.881342, 4.904335, 4.922764, 4.935397, 4.941571, 4.941417, 4.935998,
  // totalHeight(15,26, 0-49)
    4.894406, 4.87272, 4.854392, 4.839842, 4.829338, 4.822953, 4.820543, 
    4.82172, 4.82587, 4.832198, 4.839781, 4.84764, 4.854785, 4.860251, 
    4.863098, 30, 5.016332, 5.021949, 5.029336, 5.036996, 5.043603, 5.037862, 
    5.031976, 5.023129, 5.011848, 4.996982, 4.977752, 4.953513, 4.924929, 
    4.892527, 4.861219, 4.822248, 4.78804, 4.760976, 4.742573, 4.733451, 
    4.733408, 4.741605, 4.756795, 4.777483, 4.802044, 4.828778, 4.855942, 
    4.881776, 4.904565, 4.922753, 4.935126, 4.941044, 4.940664, 4.935086,
  // totalHeight(15,27, 0-49)
    4.89715, 4.875522, 4.857244, 4.842745, 4.83231, 4.826026, 4.823761, 
    4.825141, 4.829566, 4.836245, 4.84426, 4.852632, 4.860379, 4.866575, 
    4.870389, 30, 5.012642, 5.018445, 5.025831, 5.033369, 5.039788, 5.035005, 
    5.029674, 5.021203, 5.01006, 4.995123, 4.97568, 4.951184, 4.922391, 
    4.889878, 4.858337, 4.820057, 4.786572, 4.760231, 4.74251, 4.733994, 
    4.734449, 4.743031, 4.758483, 4.779317, 4.80391, 4.830564, 4.857533, 
    4.883053, 4.905414, 4.923075, 4.934859, 4.940183, 4.939286, 4.933345,
  // totalHeight(15,28, 0-49)
    4.900956, 4.87935, 4.861095, 4.846647, 4.83631, 4.830202, 4.828211, 
    4.829986, 4.834939, 4.842281, 4.851081, 4.860333, 4.869051, 4.876345, 
    4.881514, 30, 5.007342, 5.013274, 5.020514, 5.02774, 5.033801, 5.030379, 
    5.02587, 5.017995, 5.00712, 4.992149, 4.972463, 4.947652, 4.918607, 
    4.885978, 4.854132, 4.816909, 4.784528, 4.759285, 4.742601, 4.735004, 
    4.736219, 4.745374, 4.761208, 4.782232, 4.806831, 4.833304, 4.85991, 
    4.884882, 4.906523, 4.923325, 4.934174, 4.938588, 4.936932, 4.93051,
  // totalHeight(15,29, 0-49)
    4.905488, 4.883822, 4.865526, 4.851095, 4.840873, 4.835017, 4.833459, 
    4.83588, 4.841707, 4.850139, 4.860193, 4.870795, 4.8809, 4.889626, 
    4.896388, 30, 5.000063, 5.005975, 5.012874, 5.019604, 5.025175, 5.023331, 
    5.019852, 5.012797, 5.002379, 4.987502, 4.967638, 4.942543, 4.913272, 
    4.880569, 4.848407, 4.812506, 4.781537, 4.757733, 4.742431, 4.736076, 
    4.738331, 4.748291, 4.764679, 4.786003, 4.810646, 4.836909, 4.86304, 
    4.887277, 4.907935, 4.923557, 4.933121, 4.936285, 4.933587, 4.926498,
  // totalHeight(15,30, 0-49)
    4.910488, 4.888827, 4.870213, 4.855021, 4.843503, 4.83578, 4.831827, 
    4.831496, 4.834548, 4.840704, 4.849711, 4.861379, 4.875586, 4.892223, 
    4.911034, 4.954827, 4.973868, 4.991736, 5.008694, 5.022947, 5.033298, 
    5.035358, 5.033057, 5.025144, 5.012241, 4.993824, 4.97003, 4.941264, 
    4.909084, 4.874454, 4.840883, 4.805935, 4.77645, 4.754404, 4.74091, 
    4.73623, 4.739908, 4.750978, 4.768137, 4.789886, 4.814612, 4.84061, 
    4.866129, 4.889415, 4.908816, 4.922949, 4.930926, 4.932596, 4.928713, 
    4.920949,
  // totalHeight(15,31, 0-49)
    4.915942, 4.89447, 4.876083, 4.861194, 4.850078, 4.842865, 4.83952, 
    4.839871, 4.843635, 4.850474, 4.860056, 4.872119, 4.886497, 4.903143, 
    4.922074, 4.95497, 4.968733, 4.986028, 5.00144, 5.013679, 5.021948, 
    5.023351, 5.020294, 5.011942, 4.998954, 4.980783, 4.957542, 4.929637, 
    4.898599, 4.865321, 4.832775, 4.800514, 4.773793, 4.754419, 4.743352, 
    4.740744, 4.746068, 4.758324, 4.776205, 4.798216, 4.822738, 4.848071, 
    4.872464, 4.894181, 4.911629, 4.923537, 4.929198, 4.928702, 4.923073, 
    4.914211,
  // totalHeight(15,32, 0-49)
    4.921215, 4.899942, 4.881758, 4.8671, 4.856259, 4.849372, 4.846404, 
    4.847165, 4.851349, 4.858582, 4.868499, 4.880802, 4.895323, 4.912056, 
    4.93118, 4.954336, 4.96384, 4.98057, 4.994486, 5.004793, 5.011045, 
    5.011725, 5.007792, 4.99875, 4.985291, 4.966941, 4.943911, 4.916705, 
    4.886889, 4.855299, 4.824359, 4.795338, 4.771907, 4.755643, 4.747331, 
    4.746997, 4.754054, 4.767476, 4.785954, 4.808, 4.832004, 4.856267, 
    4.879059, 4.898688, 4.913652, 4.922843, 4.925797, 4.9229, 4.91548, 
    4.905674,
  // totalHeight(15,33, 0-49)
    4.92593, 4.904881, 4.886914, 4.872478, 4.861875, 4.855245, 4.852547, 
    4.853583, 4.858017, 4.865453, 4.875493, 4.887812, 4.902227, 4.91875, 
    4.937635, 4.952839, 4.959489, 4.975294, 4.98753, 4.995835, 5.000043, 
    4.999904, 4.99502, 4.985198, 4.971148, 4.952522, 4.929667, 4.903242, 
    4.874849, 4.845289, 4.816482, 4.7911, 4.771321, 4.758461, 4.753111, 
    4.755168, 4.763979, 4.778497, 4.797407, 4.819228, 4.842355, 4.865105, 
    4.885779, 4.902761, 4.914688, 4.920676, 4.920567, 4.915102, 4.905936, 
    4.895429,
  // totalHeight(15,34, 0-49)
    4.929762, 4.908973, 4.891263, 4.877086, 4.866748, 4.860384, 4.857946, 
    4.859209, 4.863815, 4.871333, 4.881327, 4.893431, 4.907422, 4.923276, 
    4.941233, 4.950496, 4.955647, 4.969988, 4.980257, 4.986433, 4.988561, 
    4.987503, 4.981656, 4.971096, 4.956528, 4.937751, 4.915259, 4.889861, 
    4.86318, 4.836005, 4.809812, 4.788346, 4.772446, 4.763155, 4.760866, 
    4.765345, 4.775867, 4.791358, 4.810493, 4.831789, 4.853648, 4.874407, 
    4.892422, 4.906191, 4.914549, 4.916904, 4.913468, 4.905375, 4.89462, 
    4.883753,
  // totalHeight(15,35, 0-49)
    4.932462, 4.911976, 4.894581, 4.880731, 4.870724, 4.864684, 4.862538, 
    4.864038, 4.868792, 4.87632, 4.886137, 4.897826, 4.911088, 4.925822, 
    4.942156, 4.947344, 4.952077, 4.964399, 4.972419, 4.976362, 4.976421, 
    4.974379, 4.967628, 4.95648, 4.941605, 4.922957, 4.901151, 4.877123, 
    4.852477, 4.828023, 4.80485, 4.787461, 4.77554, 4.769867, 4.77063, 
    4.777473, 4.789596, 4.805881, 4.824989, 4.845424, 4.865595, 4.883875, 
    4.898703, 4.908737, 4.913075, 4.911485, 4.904602, 4.893983, 4.881938, 
    4.87114,
  // totalHeight(15,36, 0-49)
    4.933903, 4.91376, 4.896746, 4.883297, 4.873699, 4.86805, 4.866251, 
    4.868015, 4.872907, 4.880397, 4.889943, 4.901053, 4.91335, 4.926611, 
    4.940794, 4.943399, 4.948446, 4.958294, 4.963863, 4.965548, 4.963623, 
    4.960588, 4.953065, 4.941565, 4.926686, 4.908533, 4.887803, 4.865521, 
    4.843225, 4.821772, 4.801928, 4.788659, 4.780696, 4.778567, 4.782275, 
    4.791337, 4.804873, 4.821717, 4.840497, 4.85971, 4.87777, 4.893103, 
    4.904272, 4.910153, 4.91017, 4.904511, 4.894277, 4.881431, 4.868542, 
    4.858325,
  // totalHeight(15,37, 0-49)
    4.934103, 4.914344, 4.897767, 4.884783, 4.875652, 4.870442, 4.86902, 
    4.871055, 4.876065, 4.883467, 4.892656, 4.903069, 4.914239, 4.925816, 
    4.937567, 4.938635, 4.944391, 4.951484, 4.954533, 4.954038, 4.950295, 
    4.946325, 4.938226, 4.926672, 4.912144, 4.894886, 4.875633, 4.855452, 
    4.83577, 4.817514, 4.801187, 4.791965, 4.787823, 4.789057, 4.795502, 
    4.806548, 4.821237, 4.838345, 4.856464, 4.874076, 4.889618, 4.9016, 
    4.908755, 4.910237, 4.905857, 4.896271, 4.883037, 4.868485, 4.855347, 
    4.846265,
  // totalHeight(15,38, 0-49)
    4.933275, 4.913924, 4.897812, 4.885321, 4.876671, 4.871897, 4.870824, 
    4.873085, 4.878146, 4.88538, 4.894122, 4.903744, 4.913695, 4.923514, 
    4.932799, 4.932977, 4.93955, 4.943816, 4.944435, 4.941947, 4.936632, 
    4.93186, 4.923436, 4.912159, 4.898354, 4.882379, 4.864967, 4.847182, 
    4.8303, 4.815341, 4.802587, 4.797229, 4.79666, 4.800972, 4.809848, 
    4.822561, 4.83807, 4.855095, 4.872189, 4.887829, 4.900504, 4.908844, 
    4.911808, 4.908888, 4.900332, 4.88727, 4.871682, 4.85616, 4.843473, 
    4.836088,
  // totalHeight(15,39, 0-49)
    4.931844, 4.912904, 4.897245, 4.885211, 4.876986, 4.87256, 4.871725, 
    4.874079, 4.879056, 4.885987, 4.894164, 4.902904, 4.911595, 4.919686, 
    4.926654, 4.926291, 4.933585, 4.935168, 4.933599, 4.929408, 4.922832, 
    4.91746, 4.909001, 4.898345, 4.885618, 4.871275, 4.856004, 4.840826, 
    4.826837, 4.815162, 4.805911, 4.804132, 4.80679, 4.813807, 4.824722, 
    4.838705, 4.85464, 4.871191, 4.88689, 4.900232, 4.909787, 4.914362, 
    4.913201, 4.906186, 4.894016, 4.878262, 4.861233, 4.845648, 4.834178, 
    4.828999,
  // totalHeight(15,40, 0-49)
    4.930457, 4.911899, 4.896629, 4.884946, 4.876993, 4.872725, 4.87191, 
    4.874125, 4.878788, 4.885204, 4.892647, 4.900396, 4.907799, 4.914251, 
    4.919162, 4.918425, 4.926207, 4.925446, 4.92205, 4.916519, 4.909047, 
    4.903338, 4.895158, 4.885455, 4.874131, 4.861706, 4.848792, 4.836337, 
    4.825235, 4.816731, 4.810798, 4.812224, 4.817683, 4.826947, 4.839435, 
    4.854232, 4.870153, 4.885829, 4.899788, 4.910583, 4.91692, 4.917839, 
    4.912915, 4.902449, 4.887573, 4.870214, 4.852869, 4.838229, 4.828725, 
    4.826172,
  // totalHeight(15,41, 0-49)
    4.929952, 4.911724, 4.896721, 4.885202, 4.877274, 4.872872, 4.871749, 
    4.873485, 4.877499, 4.883104, 4.889571, 4.896175, 4.902244, 4.907153, 
    4.910297, 4.909247, 4.917224, 4.914587, 4.909807, 4.903347, 4.895372, 
    4.889627, 4.882048, 4.873604, 4.863957, 4.853662, 4.843232, 4.833522, 
    4.825214, 4.819678, 4.816773, 4.820962, 4.828731, 4.839725, 4.853273, 
    4.868386, 4.883842, 4.898261, 4.910213, 4.918354, 4.921581, 4.919222, 
    4.911222, 4.898285, 4.881907, 4.864242, 4.847815, 4.835123, 4.828254, 
    4.828617,
  // totalHeight(15,42, 0-49)
    4.931294, 4.913325, 4.898424, 4.886817, 4.878589, 4.873669, 4.871818, 
    4.872636, 4.875574, 4.879983, 4.885159, 4.890398, 4.895037, 4.898464, 
    4.900094, 4.898733, 4.906603, 4.902615, 4.896917, 4.88995, 4.881868, 
    4.876405, 4.86973, 4.862811, 4.855051, 4.847018, 4.839118, 4.832088, 
    4.826405, 4.823557, 4.823317, 4.829775, 4.83932, 4.851501, 4.865571, 
    4.880503, 4.89507, 4.907923, 4.917725, 4.923294, 4.923772, 4.918811, 
    4.908726, 4.894571, 4.878089, 4.861507, 4.847205, 4.837363, 4.833653, 
    4.837076,
  // totalHeight(15,43, 0-49)
    4.935475, 4.917697, 4.902711, 4.890727, 4.881828, 4.875952, 4.872892, 
    4.872292, 4.873665, 4.876423, 4.879921, 4.883506, 4.886554, 4.888489, 
    4.888772, 4.887052, 4.894532, 4.889695, 4.883519, 4.876438, 4.868618, 
    4.863738, 4.85823, 4.853035, 4.847303, 4.841592, 4.836183, 4.831695, 
    4.828406, 4.827918, 4.829926, 4.83814, 4.84892, 4.86174, 4.875812, 
    4.89011, 4.90344, 4.914546, 4.922236, 4.925542, 4.923896, 4.917282, 
    4.906342, 4.892384, 4.877251, 4.863077, 4.851962, 4.845681, 4.845468, 
    4.851949,
  // totalHeight(15,44, 0-49)
    4.943389, 4.925753, 4.910508, 4.897867, 4.887924, 4.880651, 4.875891, 
    4.873359, 4.872651, 4.87327, 4.874662, 4.876251, 4.877479, 4.87783, 
    4.876827, 4.87465, 4.881481, 4.876204, 4.869909, 4.863044, 4.855793, 
    4.851745, 4.847598, 4.844251, 4.840609, 4.837198, 4.834173, 4.832032, 
    4.830871, 4.832383, 4.836201, 4.845671, 4.857166, 4.870117, 4.883736, 
    4.897036, 4.908914, 4.918256, 4.924076, 4.925666, 4.922758, 4.91564, 
    4.905199, 4.892863, 4.880429, 4.869793, 4.862683, 4.860432, 4.863861, 
    4.873267,
  // totalHeight(15,45, 0-49)
    4.955724, 4.938224, 4.922591, 4.909056, 4.897744, 4.88868, 4.881776, 
    4.876834, 4.873561, 4.871572, 4.870428, 4.86966, 4.868797, 4.867399, 
    4.865062, 4.862271, 4.868221, 4.862769, 4.856599, 4.850181, 4.843715, 
    4.840663, 4.837982, 4.836504, 4.834927, 4.833717, 4.832911, 4.832884, 
    4.833569, 4.836724, 4.841933, 4.852195, 4.863946, 4.876606, 4.889421, 
    4.901495, 4.911865, 4.919618, 4.924015, 4.924632, 4.921483, 4.915091, 
    4.906478, 4.897058, 4.888436, 4.882178, 4.879595, 4.881592, 4.888622, 
    4.900716,
  // totalHeight(15,46, 0-49)
    4.972857, 4.955551, 4.939471, 4.924886, 4.911969, 4.900812, 4.891409, 
    4.883674, 4.877432, 4.872438, 4.868383, 4.864922, 4.861692, 4.858339, 
    4.854538, 4.850924, 4.855777, 4.850251, 4.844319, 4.838459, 4.832879, 
    4.830882, 4.82966, 4.82997, 4.830338, 4.831164, 4.832362, 4.834197, 
    4.836456, 4.840928, 4.847151, 4.857822, 4.869471, 4.881536, 4.893338, 
    4.904113, 4.913095, 4.919608, 4.923187, 4.923685, 4.921351, 4.916856, 
    4.911235, 4.905757, 4.901744, 4.900376, 4.902549, 4.908782, 4.91922, 
    4.933684,
  // totalHeight(15,47, 0-49)
    4.994822, 4.977833, 4.961337, 4.945648, 4.931002, 4.917567, 4.905441, 
    4.894656, 4.885172, 4.87689, 4.869647, 4.863233, 4.857401, 4.851891, 
    4.846448, 4.841775, 4.845335, 4.839686, 4.833971, 4.828657, 4.82394, 
    4.822939, 4.823054, 4.824963, 4.827073, 4.829704, 4.832666, 4.836111, 
    4.839708, 4.845225, 4.85217, 4.862968, 4.874279, 4.885587, 4.896322, 
    4.905891, 4.913754, 4.9195, 4.922939, 4.92417, 4.923613, 4.921988, 
    4.920238, 4.919398, 4.920445, 4.924166, 4.931067, 4.941337, 4.954875, 
    4.971336,
  // totalHeight(15,48, 0-49)
    5.021287, 5.004817, 4.988027, 4.971284, 4.954903, 4.939142, 4.92421, 
    4.910266, 4.897417, 4.885714, 4.875143, 4.865629, 4.857044, 4.849217, 
    4.841962, 4.835991, 4.838085, 4.832155, 4.826528, 4.821638, 4.817649, 
    4.817477, 4.818703, 4.821928, 4.825503, 4.829668, 4.834137, 4.838961, 
    4.843709, 4.850078, 4.857544, 4.868315, 4.879192, 4.88973, 4.899494, 
    4.908081, 4.915195, 4.920693, 4.92464, 4.927336, 4.929301, 4.931226, 
    4.933884, 4.938024, 4.944261, 4.953, 4.964405, 4.978386, 4.994637, 5.01268,
  // totalHeight(15,49, 0-49)
    5.058356, 5.043217, 5.026606, 5.00895, 4.990648, 4.972076, 4.953585, 
    4.935503, 4.918123, 4.901687, 4.886375, 4.872292, 4.859453, 4.847805, 
    4.837231, 4.829314, 4.83676, 4.82897, 4.82178, 4.815975, 4.811789, 
    4.814678, 4.819662, 4.827548, 4.834721, 4.8415, 4.847211, 4.851875, 
    4.854626, 4.859023, 4.86429, 4.875, 4.885332, 4.89494, 4.903584, 
    4.911133, 4.917612, 4.923219, 4.928326, 4.933444, 4.939155, 4.946041, 
    4.9546, 4.965176, 4.977912, 4.992743, 5.009426, 5.027546, 5.046576, 
    5.065892,
  // totalHeight(16,0, 0-49)
    5.010379, 4.983305, 4.957535, 4.933589, 4.911873, 4.89267, 4.876139, 
    4.862313, 4.851107, 4.842322, 4.835676, 4.830809, 4.827321, 4.824801, 
    4.82285, 4.821224, 4.82087, 4.8188, 4.816489, 4.813863, 4.810887, 
    4.80795, 4.804797, 4.801712, 4.798837, 4.796524, 4.795112, 4.794984, 
    4.796442, 4.799865, 4.805302, 4.813079, 4.822648, 4.833603, 4.845372, 
    4.857257, 4.868512, 4.878438, 4.88649, 4.892384, 4.896164, 4.898243, 
    4.899375, 4.90057, 4.90296, 4.907646, 4.915551, 4.92732, 4.943265, 
    4.963357,
  // totalHeight(16,1, 0-49)
    4.998121, 4.971027, 4.945522, 4.922115, 4.901196, 4.88303, 4.86775, 
    4.855347, 4.845687, 4.838506, 4.833449, 4.830081, 4.827929, 4.826505, 
    4.825345, 4.824247, 4.825438, 4.823134, 4.820419, 4.817234, 4.813533, 
    4.810053, 4.806176, 4.802295, 4.798471, 4.795121, 4.792607, 4.79137, 
    4.791726, 4.794225, 4.798886, 4.806432, 4.81596, 4.827044, 4.839068, 
    4.851271, 4.86282, 4.87292, 4.880921, 4.886435, 4.889426, 4.890259, 
    4.889693, 4.888795, 4.888814, 4.891007, 4.896475, 4.906033, 4.920139, 
    4.938877,
  // totalHeight(16,2, 0-49)
    4.988944, 4.96211, 4.937086, 4.914367, 4.894336, 4.877245, 4.863204, 
    4.852176, 4.84398, 4.838302, 4.834718, 4.832727, 4.831792, 4.831364, 
    4.830914, 4.830249, 4.832897, 4.830378, 4.827298, 4.8236, 4.819216, 
    4.815224, 4.810616, 4.805884, 4.801012, 4.796468, 4.792636, 4.790017, 
    4.788951, 4.790158, 4.793639, 4.800545, 4.809657, 4.82056, 4.832631, 
    4.845079, 4.857021, 4.867584, 4.876018, 4.881814, 4.884809, 4.885249, 
    4.883801, 4.88151, 4.879666, 4.879637, 4.882692, 4.889841, 4.901728, 
    4.918592,
  // totalHeight(16,3, 0-49)
    4.98254, 4.95621, 4.931844, 4.90993, 4.890845, 4.874831, 4.861982, 
    4.852237, 4.845376, 4.841043, 4.838762, 4.837986, 4.838121, 4.838571, 
    4.838752, 4.838411, 4.842396, 4.83975, 4.836403, 4.832302, 4.827349, 
    4.822939, 4.817657, 4.812073, 4.806106, 4.800255, 4.794926, 4.790676, 
    4.787887, 4.787426, 4.789301, 4.795124, 4.80339, 4.813739, 4.82558, 
    4.838131, 4.850492, 4.86174, 4.871041, 4.877756, 4.88156, 4.882516, 
    4.881122, 4.878296, 4.87528, 4.873495, 4.874341, 4.879025, 4.888411, 
    4.902944,
  // totalHeight(16,4, 0-49)
    4.978348, 4.952726, 4.929165, 4.908149, 4.890049, 4.875096, 4.863371, 
    4.854793, 4.849114, 4.845946, 4.844783, 4.845037, 4.846092, 4.847313, 
    4.848078, 4.847959, 4.853121, 4.85051, 4.847063, 4.842731, 4.837382, 
    4.832712, 4.826875, 4.8205, 4.813451, 4.806242, 4.799288, 4.793202, 
    4.788418, 4.785934, 4.785778, 4.790048, 4.797011, 4.806389, 4.817661, 
    4.830092, 4.842803, 4.854854, 4.865345, 4.873514, 4.878854, 4.881207, 
    4.880831, 4.878424, 4.875085, 4.872192, 4.871225, 4.873564, 4.880309, 
    4.89215,
  // totalHeight(16,5, 0-49)
    4.975636, 4.950883, 4.928251, 4.908212, 4.891126, 4.877218, 4.866553, 
    4.859032, 4.85439, 4.852214, 4.851986, 4.853107, 4.85495, 4.856871, 
    4.858217, 4.858232, 4.864367, 4.862026, 4.858702, 4.854363, 4.848849, 
    4.844121, 4.837903, 4.830859, 4.822809, 4.814256, 4.805618, 4.797554, 
    4.790562, 4.785738, 4.78315, 4.785407, 4.790595, 4.798553, 4.808867, 
    4.820886, 4.833784, 4.84663, 4.858483, 4.868478, 4.87593, 4.880437, 
    4.881971, 4.880943, 4.878209, 4.875005, 4.872805, 4.87311, 4.877246, 
    4.886169,
  // totalHeight(16,6, 0-49)
    4.97359, 4.949832, 4.92823, 4.909238, 4.893208, 4.880342, 4.870695, 
    4.864148, 4.860424, 4.859102, 4.859666, 4.861528, 4.864074, 4.866668, 
    4.868656, 4.868736, 4.875587, 4.873809, 4.870874, 4.866787, 4.861371, 
    4.856816, 4.85043, 4.842885, 4.83398, 4.824172, 4.81387, 4.803766, 
    4.794423, 4.787009, 4.781643, 4.781456, 4.784411, 4.790498, 4.799439, 
    4.810699, 4.823528, 4.837036, 4.850263, 4.862264, 4.872192, 4.87941, 
    4.883584, 4.884794, 4.883579, 4.880935, 4.878224, 4.876989, 4.878732, 
    4.884682,
  // totalHeight(16,7, 0-49)
    4.971429, 4.948754, 4.928265, 4.910394, 4.895467, 4.883669, 4.87503, 
    4.869415, 4.866539, 4.865985, 4.867253, 4.869784, 4.872997, 4.876294, 
    4.879041, 4.879138, 4.8864, 4.885508, 4.883248, 4.879677, 4.874628, 
    4.870487, 4.864169, 4.856335, 4.846771, 4.835867, 4.824009, 4.811897, 
    4.800161, 4.789993, 4.781582, 4.778574, 4.778876, 4.782658, 4.789808, 
    4.799926, 4.812365, 4.826291, 4.840752, 4.85474, 4.86728, 4.877518, 
    4.884831, 4.888952, 4.890053, 4.888813, 4.886382, 4.88424, 4.883992, 
    4.887099,
  // totalHeight(16,8, 0-49)
    4.9685, 4.946961, 4.927648, 4.910966, 4.897206, 4.886523, 4.878919, 
    4.874241, 4.872197, 4.872381, 4.874321, 4.877502, 4.881399, 4.885472, 
    4.889145, 4.889234, 4.896564, 4.896873, 4.895561, 4.892765, 4.888341, 
    4.884839, 4.878826, 4.870933, 4.860958, 4.849187, 4.835968, 4.82198, 
    4.807916, 4.794942, 4.783319, 4.777194, 4.774482, 4.775564, 4.780519, 
    4.789104, 4.800787, 4.814806, 4.83023, 4.846014, 4.861082, 4.874398, 
    4.885083, 4.892534, 4.896551, 4.897444, 4.896061, 4.893718, 4.892021, 
    4.892599,
  // totalHeight(16,9, 0-49)
    4.964339, 4.943954, 4.92586, 4.910425, 4.897897, 4.888393, 4.88188, 
    4.878181, 4.876997, 4.87794, 4.88057, 4.88443, 4.889064, 4.894015, 
    4.898808, 4.898908, 4.90595, 4.907724, 4.907599, 4.905803, 4.90224, 
    4.89956, 4.894073, 4.886361, 4.876246, 4.863895, 4.849592, 4.833972, 
    4.817759, 4.802047, 4.787168, 4.777723, 4.771718, 4.769764, 4.772158, 
    4.778826, 4.789371, 4.803106, 4.81913, 4.836383, 4.853708, 4.869932, 
    4.883956, 4.894887, 4.902172, 4.905732, 4.906059, 4.904214, 4.901698, 
    4.900219,
  // totalHeight(16,10, 0-49)
    4.958708, 4.939458, 4.922597, 4.908445, 4.897206, 4.888947, 4.88359, 
    4.880938, 4.880676, 4.882433, 4.885808, 4.890401, 4.895841, 4.901774, 
    4.907865, 4.908079, 4.914513, 4.917924, 4.919169, 4.918551, 4.916037, 
    4.914315, 4.909543, 4.902239, 4.892272, 4.879665, 4.864626, 4.847709, 
    4.829641, 4.811388, 4.793344, 4.780487, 4.770998, 4.76575, 4.765265, 
    4.769666, 4.77869, 4.791737, 4.807944, 4.826241, 4.845419, 4.864198, 
    4.881311, 4.895623, 4.906263, 4.912791, 4.915321, 4.914591, 4.911907, 
    4.908954,
  // totalHeight(16,11, 0-49)
    4.951579, 4.933411, 4.917763, 4.904904, 4.894985, 4.88802, 4.883884, 
    4.882345, 4.883079, 4.88572, 4.889904, 4.895293, 4.901602, 4.9086, 
    4.916114, 4.916668, 4.922263, 4.927371, 4.930091, 4.930777, 4.929453, 
    4.928766, 4.924852, 4.918157, 4.908612, 4.89609, 4.88071, 4.862903, 
    4.84337, 4.822893, 4.801913, 4.785665, 4.77261, 4.763888, 4.760275, 
    4.762101, 4.769247, 4.781209, 4.797158, 4.816027, 4.836568, 4.857426, 
    4.877209, 4.894594, 4.908454, 4.918019, 4.923042, 4.923909, 4.92166, 
    4.917865,
  // totalHeight(16,12, 0-49)
    4.94311, 4.925941, 4.911447, 4.899851, 4.89125, 4.885598, 4.882725, 
    4.882352, 4.884141, 4.887729, 4.892781, 4.899015, 4.906228, 4.914317, 
    4.923285, 4.924597, 4.929274, 4.936002, 4.940219, 4.942276, 4.942241, 
    4.942596, 4.939634, 4.933708, 4.924829, 4.912722, 4.897404, 4.879156, 
    4.858614, 4.836325, 4.812768, 4.793261, 4.776662, 4.764382, 4.757468, 
    4.756468, 4.761423, 4.771923, 4.787184, 4.80614, 4.827521, 4.849919, 
    4.871853, 4.891866, 4.908628, 4.921103, 4.928713, 4.931497, 4.930191, 
    4.926173,
  // totalHeight(16,13, 0-49)
    4.933587, 4.917305, 4.903876, 4.893475, 4.886146, 4.881787, 4.880175, 
    4.88099, 4.883869, 4.888443, 4.894396, 4.901491, 4.909599, 4.918728, 
    4.929043, 4.931781, 4.935657, 4.943816, 4.94947, 4.952912, 4.954217, 
    4.955572, 4.953596, 4.948547, 4.940525, 4.92912, 4.914241, 4.895998, 
    4.874925, 4.8513, 4.825628, 4.803096, 4.783074, 4.767251, 4.756944, 
    4.752938, 4.755445, 4.764153, 4.778327, 4.796912, 4.81862, 4.842006, 
    4.865535, 4.887653, 4.906889, 4.921998, 4.932122, 4.936985, 4.937004, 
    4.933322,
  // totalHeight(16,14, 0-49)
    4.923371, 4.90785, 4.895366, 4.886055, 4.879909, 4.876776, 4.87638, 
    4.87836, 4.882319, 4.887879, 4.894729, 4.902659, 4.9116, 4.921633, 
    4.933037, 4.938135, 4.941565, 4.95087, 4.957839, 4.962636, 4.965298, 
    4.967563, 4.966561, 4.962437, 4.955395, 4.944908, 4.93078, 4.912937, 
    4.891786, 4.867318, 4.84006, 4.814806, 4.791577, 4.772316, 4.758617, 
    4.751506, 4.751376, 4.758027, 4.770776, 4.788579, 4.810141, 4.833998, 
    4.858574, 4.882263, 4.903494, 4.920869, 4.933316, 4.940278, 4.941876, 
    4.938986,
  // totalHeight(16,15, 0-49)
    4.912854, 4.897959, 4.88628, 4.877921, 4.87283, 4.870809, 4.871537, 
    4.874606, 4.87959, 4.886088, 4.893784, 4.90248, 4.912133, 4.922858, 
    4.93496, 4.94358, 4.947157, 4.957278, 4.965407, 4.971506, 4.97552, 
    4.978578, 4.978491, 4.975286, 4.969269, 4.959824, 4.946657, 4.929514, 
    4.908661, 4.883808, 4.855515, 4.827887, 4.801735, 4.779232, 4.762231, 
    4.752002, 4.749129, 4.753531, 4.764589, 4.781275, 4.80229, 4.826159, 
    4.851291, 4.876046, 4.898795, 4.918036, 4.932535, 4.941511, 4.944815, 
    4.943059,
  // totalHeight(16,16, 0-49)
    4.902413, 4.888007, 4.876982, 4.869414, 4.865215, 4.864151, 4.865855, 
    4.869885, 4.87578, 4.883116, 4.891562, 4.900916, 4.911123, 4.922285, 
    4.934649, 4.948032, 4.952551, 4.96318, 4.972324, 4.979673, 4.985033, 
    4.98876, 4.989505, 4.98716, 4.982129, 4.973736, 4.961613, 4.945337, 
    4.92504, 4.900175, 4.871372, 4.841729, 4.81299, 4.787511, 4.767387, 
    4.75412, 4.748487, 4.750541, 4.759723, 4.775039, 4.795194, 4.818704, 
    4.843974, 4.86935, 4.893178, 4.913892, 4.930142, 4.940972, 4.946005, 
    4.945608,
  // totalHeight(16,17, 0-49)
    4.892386, 4.878341, 4.867813, 4.860855, 4.857354, 4.857041, 4.859523, 
    4.864323, 4.870955, 4.878976, 4.88804, 4.897923, 4.908541, 4.919922, 
    4.932185, 4.951418, 4.957764, 4.968699, 4.978784, 4.987378, 4.994099, 
    4.998383, 4.999869, 4.998282, 4.994113, 4.986661, 4.975505, 4.960099, 
    4.940459, 4.915834, 4.886974, 4.855661, 4.824695, 4.796576, 4.773589, 
    4.757456, 4.749144, 4.748833, 4.756054, 4.769843, 4.78891, 4.811782, 
    4.836864, 4.862501, 4.88703, 4.908854, 4.926551, 4.939031, 4.945736, 
    4.946805,
  // totalHeight(16,18, 0-49)
    4.883057, 4.86925, 4.859056, 4.852509, 4.849472, 4.849656, 4.852646, 
    4.857956, 4.865088, 4.873597, 4.88313, 4.893447, 4.904416, 4.91596, 
    4.927983, 4.95368, 4.962641, 4.973895, 4.984979, 4.994907, 5.003065, 
    5.007842, 5.009997, 5.009035, 5.005515, 4.998745, 4.988299, 4.973565, 
    4.954499, 4.930216, 4.901648, 4.868981, 4.836173, 4.805798, 4.780288, 
    4.761552, 4.750729, 4.748141, 4.753402, 4.76559, 4.783442, 4.805486, 
    4.83014, 4.855759, 4.880685, 4.903311, 4.922166, 4.936076, 4.944336, 
    4.946891,
  // totalHeight(16,19, 0-49)
    4.874649, 4.860956, 4.850918, 4.844546, 4.841686, 4.842038, 4.845186, 
    4.850657, 4.857982, 4.866745, 4.876626, 4.887396, 4.898871, 4.910821, 
    4.922827, 4.954803, 4.966801, 4.978681, 4.991045, 5.002561, 5.012359, 
    5.017647, 5.020454, 5.019977, 5.016799, 5.010279, 5.000051, 4.985547, 
    4.966752, 4.942739, 4.9147, 4.880971, 4.846727, 4.814543, 4.786932, 
    4.765944, 4.752872, 4.748176, 4.751559, 4.76216, 4.778742, 4.799853, 
    4.823924, 4.849325, 4.874414, 4.897583, 4.917346, 4.932465, 4.942127, 
    4.946119,
  // totalHeight(16,20, 0-49)
    4.867816, 4.854584, 4.845321, 4.840126, 4.838893, 4.841312, 4.846864, 
    4.85486, 4.864492, 4.874896, 4.885221, 4.894706, 4.902756, 4.909014, 
    4.913389, 30, 4.987489, 4.991956, 4.99765, 5.003873, 5.010102, 5.012218, 
    5.01397, 5.014071, 5.012827, 5.009157, 5.002196, 4.990902, 4.974914, 
    4.953116, 4.927007, 4.893116, 4.858006, 4.824359, 4.79484, 4.771689, 
    4.756392, 4.749557, 4.751001, 4.759923, 4.775121, 4.79516, 4.818483, 
    4.843477, 4.868512, 4.891992, 4.912422, 4.928527, 4.93941, 4.944731,
  // totalHeight(16,21, 0-49)
    4.861976, 4.848943, 4.839874, 4.834837, 4.833697, 4.836112, 4.841539, 
    4.849289, 4.858567, 4.868547, 4.878441, 4.887538, 4.895265, 4.901219, 
    4.905196, 30, 4.992397, 4.997305, 5.003582, 5.010384, 5.017054, 5.017688, 
    5.018337, 5.017498, 5.015707, 5.011953, 5.005382, 4.994881, 4.979984, 
    4.959462, 4.935041, 4.90137, 4.866254, 4.832252, 4.801982, 4.777731, 
    4.761089, 4.752796, 4.752783, 4.760341, 4.774326, 4.793342, 4.815856, 
    4.840277, 4.864996, 4.888429, 4.909086, 4.925674, 4.937243, 4.943362,
  // totalHeight(16,22, 0-49)
    4.857375, 4.844437, 4.83546, 4.830493, 4.82939, 4.83179, 4.837147, 
    4.844765, 4.853857, 4.863614, 4.873266, 4.882125, 4.889603, 4.895244, 
    4.898731, 30, 4.995681, 5.000916, 5.007755, 5.015225, 5.022527, 5.022017, 
    5.021948, 5.020552, 5.018504, 5.014805, 5.008574, 4.99863, 4.984444, 
    4.964725, 4.941484, 4.907679, 4.872356, 4.837974, 4.807092, 4.781999, 
    4.764341, 4.754937, 4.753801, 4.760295, 4.773324, 4.791523, 4.813382, 
    4.837328, 4.86177, 4.885137, 4.905946, 4.922899, 4.935011, 4.941789,
  // totalHeight(16,23, 0-49)
    4.854089, 4.841188, 4.83224, 4.82729, 4.82618, 4.828554, 4.833859, 
    4.841405, 4.850407, 4.860065, 4.869614, 4.878358, 4.885695, 4.891115, 
    4.894202, 30, 4.998227, 5.003655, 5.010888, 5.018858, 5.026659, 5.025187, 
    5.024527, 5.02266, 5.020362, 5.016635, 5.010581, 5.000975, 4.98724, 
    4.968055, 4.945672, 4.911668, 4.876164, 4.841541, 4.810292, 4.784687, 
    4.76639, 4.756265, 4.754383, 4.760154, 4.772521, 4.790148, 4.811541, 
    4.835138, 4.85936, 4.882646, 4.903519, 4.920674, 4.933112, 4.940302,
  // totalHeight(16,24, 0-49)
    4.852131, 4.839238, 4.830288, 4.825319, 4.824179, 4.826513, 4.831777, 
    4.839285, 4.848259, 4.8579, 4.867444, 4.876188, 4.88351, 4.888863, 
    4.891764, 30, 5.000336, 5.005877, 5.013352, 5.021645, 5.029784, 5.027698, 
    5.026659, 5.024476, 5.021976, 5.018165, 5.01214, 5.002656, 4.989122, 
    4.970199, 4.948319, 4.914134, 4.878489, 4.843718, 4.812261, 4.786366, 
    4.767694, 4.757131, 4.754774, 4.760069, 4.771986, 4.789208, 4.810258, 
    4.833585, 4.857615, 4.880801, 4.901666, 4.918907, 4.931514, 4.938937,
  // totalHeight(16,25, 0-49)
    4.85146, 4.838564, 4.829591, 4.824589, 4.823408, 4.825703, 4.830941, 
    4.838443, 4.847441, 4.857141, 4.866776, 4.875635, 4.883084, 4.888557, 
    4.891555, 30, 5.001617, 5.00724, 5.014842, 5.023288, 5.03158, 5.02933, 
    5.02819, 5.025898, 5.02329, 5.019381, 5.01327, 5.003716, 4.990139, 
    4.971201, 4.949409, 4.915092, 4.87936, 4.844524, 4.813005, 4.787022, 
    4.768224, 4.757499, 4.754951, 4.760036, 4.771738, 4.788752, 4.809611, 
    4.83277, 4.856662, 4.879742, 4.900535, 4.917737, 4.930336, 4.937777,
  // totalHeight(16,26, 0-49)
    4.851977, 4.839075, 4.830077, 4.825035, 4.82382, 4.826095, 4.831341, 
    4.838893, 4.847992, 4.857843, 4.867679, 4.876782, 4.884514, 4.890315, 
    4.893711, 30, 5.001983, 5.007671, 5.015292, 5.023718, 5.031972, 5.030043, 
    5.029104, 5.026941, 5.024355, 5.020361, 5.014077, 5.004286, 4.990434, 
    4.971213, 4.949087, 4.914718, 4.878968, 4.844158, 4.812709, 4.786823, 
    4.768129, 4.757494, 4.755009, 4.760123, 4.771822, 4.788801, 4.809599, 
    4.832676, 4.856466, 4.87942, 4.900066, 4.917099, 4.929512, 4.936756,
  // totalHeight(16,27, 0-49)
    4.853549, 4.84063, 4.831599, 4.826528, 4.825302, 4.827601, 4.832926, 
    4.840624, 4.849943, 4.860089, 4.870278, 4.879788, 4.887972, 4.894296, 
    4.898354, 30, 5.001553, 5.007257, 5.014753, 5.022965, 5.030978, 5.02979, 
    5.029314, 5.027491, 5.025039, 5.020969, 5.014422, 5.00423, 4.989888, 
    4.970133, 4.947292, 4.912957, 4.877278, 4.842611, 4.811395, 4.785818, 
    4.767478, 4.757198, 4.755036, 4.760416, 4.772312, 4.789418, 4.810269, 
    4.833325, 4.857021, 4.879806, 4.900201, 4.916908, 4.928932, 4.935752,
  // totalHeight(16,28, 0-49)
    4.855995, 4.843037, 4.833967, 4.828879, 4.827681, 4.830082, 4.835604, 
    4.843608, 4.853339, 4.863991, 4.874754, 4.884873, 4.89369, 4.900697, 
    4.905574, 30, 5.000744, 5.006339, 5.013515, 5.021286, 5.028846, 5.028683, 
    5.02886, 5.027533, 5.025298, 5.021149, 5.014251, 5.003506, 4.988485, 
    4.967993, 4.944139, 4.909925, 4.874425, 4.840048, 4.809262, 4.78423, 
    4.766501, 4.756835, 4.75523, 4.761073, 4.773315, 4.790642, 4.811593, 
    4.834626, 4.858176, 4.88069, 4.900694, 4.916894, 4.928325, 4.934512,
  // totalHeight(16,29, 0-49)
    4.859104, 4.846059, 4.836926, 4.831833, 4.830725, 4.833347, 4.839246, 
    4.847798, 4.858232, 4.869702, 4.881335, 4.892307, 4.901924, 4.909692, 
    4.91538, 30, 4.999225, 5.004516, 5.011139, 5.018236, 5.025145, 5.026101, 
    5.027013, 5.026284, 5.024335, 5.02012, 5.012819, 5.001411, 4.985559, 
    4.964156, 4.939056, 4.904996, 4.869781, 4.835892, 4.805812, 4.781667, 
    4.764914, 4.756218, 4.755496, 4.762076, 4.774881, 4.792583, 4.813718, 
    4.836743, 4.86009, 4.882205, 4.90162, 4.917064, 4.927612, 4.93287,
  // totalHeight(16,30, 0-49)
    4.862476, 4.849107, 4.839384, 4.833349, 4.830894, 4.831782, 4.835658, 
    4.842111, 4.850717, 4.861089, 4.872904, 4.885905, 4.899866, 4.914509, 
    4.92938, 4.966947, 4.978901, 4.992922, 5.007429, 5.020907, 5.032383, 
    5.037577, 5.040587, 5.040208, 5.037008, 5.03027, 5.019615, 5.004519, 
    4.98509, 4.960538, 4.932539, 4.897691, 4.862357, 4.828973, 4.799906, 
    4.777106, 4.761838, 4.754601, 4.75519, 4.762854, 4.776481, 4.794729, 
    4.81613, 4.839152, 4.862225, 4.883802, 4.902434, 4.91689, 4.926324, 
    4.930448,
  // totalHeight(16,31, 0-49)
    4.866781, 4.853611, 4.844128, 4.83839, 4.836299, 4.837609, 4.84195, 
    4.848881, 4.857934, 4.868675, 4.880737, 4.893844, 4.9078, 4.922468, 
    4.937697, 4.967824, 4.977847, 4.991458, 5.004806, 5.016727, 5.02653, 
    5.031267, 5.033574, 5.032618, 5.028995, 5.021968, 5.011114, 4.995862, 
    4.976276, 4.951561, 4.923069, 4.889333, 4.855425, 4.823767, 4.796635, 
    4.775844, 4.762507, 4.756995, 4.759011, 4.767756, 4.782095, 4.800686, 
    4.822061, 4.844687, 4.867003, 4.887477, 4.904691, 4.917486, 4.925124, 
    4.927476,
  // totalHeight(16,32, 0-49)
    4.871303, 4.858335, 4.849073, 4.843582, 4.841766, 4.843366, 4.848002, 
    4.855215, 4.864517, 4.875458, 4.887661, 4.900854, 4.91489, 4.929732, 
    4.945438, 4.968321, 4.976445, 4.989829, 5.002178, 5.012691, 5.02094, 
    5.025236, 5.026824, 5.025161, 5.020825, 5.013091, 5.001563, 4.985727, 
    4.965698, 4.940761, 4.912001, 4.879725, 4.847709, 4.81828, 4.793566, 
    4.775197, 4.764112, 4.760547, 4.764117, 4.773983, 4.788996, 4.807811, 
    4.82897, 4.850946, 4.872193, 4.891208, 4.906636, 4.917415, 4.922964, 
    4.92335,
  // totalHeight(16,33, 0-49)
    4.875925, 4.863193, 4.854173, 4.84893, 4.847354, 4.84918, 4.854009, 
    4.861369, 4.870765, 4.881741, 4.893917, 4.907042, 4.921004, 4.935845, 
    4.951768, 4.968263, 4.974986, 4.988035, 4.999339, 5.008449, 5.015163, 
    5.01895, 5.019767, 5.017297, 5.012066, 5.003394, 4.99095, 4.974339, 
    4.95378, 4.928711, 4.900013, 4.869541, 4.839824, 4.813044, 4.791133, 
    4.775503, 4.766909, 4.765444, 4.770644, 4.78163, 4.797239, 4.816132, 
    4.836852, 4.857888, 4.877718, 4.894889, 4.908136, 4.916543, 4.919724, 
    4.917984,
  // totalHeight(16,34, 0-49)
    4.880545, 4.868095, 4.859358, 4.854384, 4.85305, 4.855068, 4.860024, 
    4.867435, 4.876794, 4.887642, 4.899608, 4.912449, 4.926073, 4.940565, 
    4.956202, 4.967526, 4.973517, 4.985917, 4.996002, 5.003626, 5.008771, 
    5.011938, 5.011914, 5.00858, 5.002374, 4.992685, 4.979272, 4.961896, 
    4.940898, 4.915932, 4.887727, 4.859404, 4.832354, 4.80857, 4.789754, 
    4.777088, 4.771133, 4.771847, 4.778687, 4.790736, 4.806821, 4.825599, 
    4.845624, 4.865399, 4.883441, 4.89837, 4.909048, 4.914743, 4.915324, 
    4.911375,
  // totalHeight(16,35, 0-49)
    4.885081, 4.87296, 4.864542, 4.85986, 4.858766, 4.86095, 4.865981, 
    4.873355, 4.882562, 4.893137, 4.904713, 4.917045, 4.930042, 4.943787, 
    4.95856, 4.96601, 4.971895, 4.98324, 4.991876, 4.997907, 5.001445, 
    5.003863, 5.002946, 4.998738, 4.991569, 4.980916, 4.966636, 4.948666, 
    4.927465, 4.902946, 4.87573, 4.849896, 4.825834, 4.805314, 4.78979, 
    4.780211, 4.776949, 4.779835, 4.788252, 4.801247, 4.817632, 4.836062, 
    4.855099, 4.87327, 4.889144, 4.901443, 4.909194, 4.911911, 4.909752, 
    4.903614,
  // totalHeight(16,36, 0-49)
    4.889462, 4.877706, 4.869629, 4.86524, 4.864367, 4.866679, 4.871722, 
    4.878978, 4.887927, 4.898099, 4.909123, 4.920747, 4.932858, 4.9455, 
    4.958887, 4.963627, 4.969875, 4.979753, 4.986724, 4.99107, 4.992982, 
    4.994537, 4.992704, 4.987673, 4.979637, 4.968187, 4.95327, 4.935, 
    4.913944, 4.890288, 4.86458, 4.841549, 4.820729, 4.803648, 4.791512, 
    4.78504, 4.784429, 4.789392, 4.799244, 4.812998, 4.82945, 4.847256, 
    4.864984, 4.881196, 4.894536, 4.903861, 4.908413, 4.907989, 4.90308, 
    4.894912,
  // totalHeight(16,37, 0-49)
    4.893633, 4.882252, 4.874506, 4.870379, 4.869679, 4.872052, 4.877029, 
    4.88408, 4.892673, 4.902333, 4.912676, 4.923434, 4.934464, 4.94574, 
    4.957366, 4.960308, 4.967186, 4.975255, 4.980393, 4.983005, 4.983312, 
    4.983918, 4.981193, 4.975446, 4.966719, 4.954725, 4.939501, 4.921314, 
    4.900814, 4.878473, 4.854766, 4.834799, 4.817393, 4.803834, 4.79508, 
    4.791636, 4.793539, 4.800397, 4.811465, 4.825723, 4.841955, 4.858814, 
    4.87489, 4.888796, 4.899277, 4.905368, 4.906568, 4.902996, 4.895502, 
    4.885627,
  // totalHeight(16,38, 0-49)
    4.897552, 4.886523, 4.879058, 4.875122, 4.874506, 4.876844, 4.881657, 
    4.888404, 4.896548, 4.905604, 4.915175, 4.924968, 4.934794, 4.944555, 
    4.954224, 4.956, 4.963574, 4.969604, 4.972828, 4.973719, 4.972487, 
    4.972108, 4.968562, 4.962262, 4.953082, 4.940866, 4.925722, 4.908052, 
    4.888546, 4.867952, 4.846678, 4.82996, 4.816054, 4.805999, 4.800521, 
    4.799932, 4.804125, 4.812616, 4.824606, 4.83905, 4.854722, 4.870285, 
    4.884364, 4.895648, 4.903024, 4.905744, 4.903603, 4.897072, 4.887355, 
    4.876265,
  // totalHeight(16,39, 0-49)
    4.901218, 4.89047, 4.88319, 4.879328, 4.878665, 4.880836, 4.885359, 
    4.891698, 4.899304, 4.907685, 4.916423, 4.925197, 4.933774, 4.94198, 
    4.94967, 4.950666, 4.958837, 4.962734, 4.964062, 4.96331, 4.960653, 
    4.959311, 4.955066, 4.948422, 4.939073, 4.926993, 4.912344, 4.89563, 
    4.877538, 4.859074, 4.840569, 4.827199, 4.81678, 4.810116, 4.807721, 
    4.809731, 4.815915, 4.825707, 4.838266, 4.852526, 4.867264, 4.881167, 
    4.892925, 4.901339, 4.905478, 4.904854, 4.89959, 4.890512, 4.879136, 
    4.86748,
  // totalHeight(16,40, 0-49)
    4.904684, 4.894101, 4.886861, 4.882905, 4.882024, 4.883858, 4.887946, 
    4.893749, 4.900727, 4.90837, 4.916239, 4.923985, 4.931323, 4.938021, 
    4.943837, 4.94427, 4.952819, 4.954637, 4.954183, 4.951932, 4.948014, 
    4.94579, 4.941018, 4.934273, 4.925064, 4.913489, 4.89974, 4.884389, 
    4.868077, 4.852043, 4.83653, 4.826512, 4.819475, 4.816006, 4.816424, 
    4.820711, 4.828525, 4.839235, 4.851963, 4.865639, 4.879057, 4.89096, 
    4.900132, 4.905531, 4.906458, 4.902721, 4.89478, 4.883789, 4.871507, 
    4.860053,
  // totalHeight(16,41, 0-49)
    4.908092, 4.897519, 4.89013, 4.885876, 4.884562, 4.88586, 4.889328, 
    4.894451, 4.90069, 4.907524, 4.914495, 4.921216, 4.927366, 4.932658, 
    4.93679, 4.93676, 4.945415, 4.945338, 4.943303, 4.939752, 4.934779, 
    4.93182, 4.926731, 4.920149, 4.911396, 4.900678, 4.888195, 4.874551, 
    4.86031, 4.846904, 4.834485, 4.827735, 4.823891, 4.823347, 4.826247, 
    4.832436, 4.841479, 4.852689, 4.86517, 4.87786, 4.889602, 4.899222, 
    4.905647, 4.908044, 4.905981, 4.899584, 4.889641, 4.877569, 4.865269, 
    4.854838,
  // totalHeight(16,42, 0-49)
    4.911717, 4.900965, 4.893209, 4.888418, 4.886428, 4.886953, 4.889586, 
    4.893843, 4.899196, 4.905123, 4.911144, 4.91684, 4.921854, 4.925863, 
    4.928534, 4.928086, 4.936563, 4.934877, 4.931522, 4.926918, 4.92114, 
    4.917643, 4.912477, 4.906325, 4.89833, 4.888782, 4.877871, 4.866199, 
    4.854226, 4.843546, 4.834213, 4.830557, 4.829648, 4.831701, 4.836706, 
    4.84439, 4.854242, 4.865532, 4.877361, 4.888703, 4.898479, 4.905645, 
    4.909317, 4.908913, 4.904303, 4.895933, 4.88486, 4.872675, 4.861303, 
    4.852696,
  // totalHeight(16,43, 0-49)
    4.915979, 4.904849, 4.896491, 4.890907, 4.887977, 4.887463, 4.889009, 
    4.892169, 4.896441, 4.901309, 4.90628, 4.910909, 4.914815, 4.91765, 
    4.919073, 4.918221, 4.926271, 4.923316, 4.918942, 4.91356, 4.907251, 
    4.903452, 4.898461, 4.892997, 4.886028, 4.877912, 4.868806, 4.859283, 
    4.849682, 4.841722, 4.835365, 4.834563, 4.836274, 4.840557, 4.847266, 
    4.856031, 4.866275, 4.877251, 4.888074, 4.897788, 4.905428, 4.910126, 
    4.911233, 4.908454, 4.901965, 4.892494, 4.881298, 4.870026, 4.860497, 
    4.854419,
  // totalHeight(16,44, 0-49)
    4.921442, 4.909743, 4.900558, 4.893926, 4.889781, 4.887942, 4.888114, 
    4.889902, 4.892839, 4.89643, 4.900186, 4.903648, 4.906418, 4.90814, 
    4.908477, 4.907215, 4.914638, 4.910761, 4.905677, 4.899805, 4.89325, 
    4.8894, 4.884832, 4.880281, 4.874562, 4.868074, 4.860928, 4.853642, 
    4.846432, 4.841105, 4.837529, 4.839285, 4.843264, 4.849389, 4.857398, 
    4.866843, 4.877102, 4.887429, 4.896988, 4.90492, 4.910418, 4.912833, 
    4.911785, 4.907272, 4.89976, 4.890192, 4.879921, 4.87054, 4.863652, 
    4.860648,
  // totalHeight(16,45, 0-49)
    4.928774, 4.916354, 4.906143, 4.89823, 4.892606, 4.889152, 4.887639, 
    4.887737, 4.889032, 4.891066, 4.893369, 4.895489, 4.897025, 4.897626, 
    4.89697, 4.895264, 4.901911, 4.897421, 4.891912, 4.885824, 4.879295, 
    4.875637, 4.871709, 4.868249, 4.863946, 4.85921, 4.854095, 4.849058, 
    4.844183, 4.84133, 4.840287, 4.844272, 4.850154, 4.857734, 4.866662, 
    4.876428, 4.886393, 4.895836, 4.903998, 4.910158, 4.913705, 4.914233, 
    4.911644, 4.906223, 4.898661, 4.890035, 4.881682, 4.875031, 4.871395, 
    4.871812,
  // totalHeight(16,46, 0-49)
    4.93868, 4.925437, 4.914054, 4.904667, 4.897326, 4.891982, 4.888477, 
    4.886553, 4.885867, 4.886013, 4.886566, 4.887105, 4.88724, 4.886635, 
    4.884993, 4.88277, 4.888525, 4.883657, 4.877955, 4.871884, 4.865617, 
    4.862357, 4.859235, 4.856978, 4.854181, 4.851244, 4.848159, 4.845309, 
    4.842661, 4.842082, 4.843284, 4.849162, 4.856587, 4.865265, 4.874779, 
    4.88458, 4.894042, 4.902493, 4.909286, 4.913868, 4.915846, 4.915076, 
    4.911729, 4.906325, 4.899712, 4.892994, 4.887399, 4.884111, 4.884117, 
    4.888099,
  // totalHeight(16,47, 0-49)
    4.951799, 4.937706, 4.925067, 4.914071, 4.904827, 4.897355, 4.891575, 
    4.887312, 4.884302, 4.88222, 4.880702, 4.879376, 4.87789, 4.875928, 
    4.873226, 4.870365, 4.875134, 4.870023, 4.864284, 4.858397, 4.852556, 
    4.849838, 4.847615, 4.846592, 4.845309, 4.844142, 4.843019, 4.842241, 
    4.841671, 4.843141, 4.846299, 4.853746, 4.862389, 4.871863, 4.881702, 
    4.891355, 4.900224, 4.907723, 4.913341, 4.916712, 4.917672, 4.916331, 
    4.913086, 4.908631, 4.903881, 4.899878, 4.897662, 4.89813, 4.901938, 
    4.909441,
  // totalHeight(16,48, 0-49)
    4.968619, 4.953721, 4.939814, 4.927141, 4.915872, 4.906098, 4.897817, 
    4.890945, 4.885314, 4.880691, 4.876794, 4.873322, 4.869973, 4.866468, 
    4.862566, 4.858901, 4.862593, 4.857264, 4.85155, 4.845926, 4.840598, 
    4.838478, 4.837162, 4.837315, 4.837472, 4.837968, 4.838675, 4.839813, 
    4.841158, 4.844455, 4.849295, 4.858031, 4.867624, 4.877662, 4.887666, 
    4.897097, 4.905418, 4.912148, 4.916932, 4.919597, 4.920197, 4.91906, 
    4.916761, 4.914085, 4.911936, 4.911226, 4.912759, 4.917141, 4.92471, 
    4.935537,
  // totalHeight(16,49, 0-49)
    4.997341, 4.981748, 4.96641, 4.95162, 4.937616, 4.924573, 4.9126, 
    4.901742, 4.89198, 4.883229, 4.875348, 4.868152, 4.861418, 4.854907, 
    4.848384, 4.843278, 4.852906, 4.845834, 4.83861, 4.832042, 4.8264, 
    4.827126, 4.82929, 4.833854, 4.837558, 4.840845, 4.843235, 4.844953, 
    4.845376, 4.847987, 4.852074, 4.862319, 4.872993, 4.88364, 4.893794, 
    4.902972, 4.910752, 4.916822, 4.921046, 4.923507, 4.924527, 4.92465, 
    4.9246, 4.925184, 4.927189, 4.931278, 4.93792, 4.947337, 4.959503, 
    4.974175,
  // totalHeight(17,0, 0-49)
    4.932086, 4.910845, 4.892358, 4.876889, 4.864563, 4.855368, 4.849143, 
    4.845583, 4.844279, 4.84473, 4.846404, 4.84877, 4.851345, 4.853716, 
    4.855547, 4.85666, 4.858193, 4.857396, 4.855773, 4.853347, 4.850139, 
    4.846555, 4.84232, 4.837674, 4.832701, 4.827689, 4.822936, 4.818818, 
    4.815685, 4.813998, 4.813952, 4.81605, 4.819995, 4.825649, 4.832704, 
    4.840699, 4.849057, 4.857137, 4.864295, 4.869975, 4.873768, 4.8755, 
    4.875279, 4.87353, 4.870981, 4.868604, 4.867512, 4.868828, 4.873548, 
    4.882422,
  // totalHeight(17,1, 0-49)
    4.927293, 4.906449, 4.888511, 4.873724, 4.862199, 4.853904, 4.848652, 
    4.846119, 4.845862, 4.847353, 4.850029, 4.853331, 4.856744, 4.859819, 
    4.862175, 4.863629, 4.866576, 4.865678, 4.863865, 4.861151, 4.857523, 
    4.853695, 4.849001, 4.843752, 4.837935, 4.831862, 4.825829, 4.820256, 
    4.815511, 4.812222, 4.810579, 4.811505, 4.814435, 4.819283, 4.825787, 
    4.83351, 4.841879, 4.850229, 4.85787, 4.864164, 4.868599, 4.870879, 
    4.870985, 4.869229, 4.866257, 4.863015, 4.860652, 4.860381, 4.863338, 
    4.87043,
  // totalHeight(17,2, 0-49)
    4.925047, 4.904743, 4.887443, 4.873371, 4.862625, 4.855145, 4.85073, 
    4.849032, 4.849593, 4.851871, 4.855292, 4.859291, 4.863336, 4.866961, 
    4.86975, 4.871462, 4.875763, 4.874875, 4.873009, 4.870171, 4.866305, 
    4.862421, 4.857438, 4.851728, 4.845177, 4.838098, 4.830777, 4.823665, 
    4.817146, 4.812004, 4.80843, 4.807797, 4.809296, 4.812929, 4.81851, 
    4.825661, 4.833847, 4.842411, 4.850638, 4.857832, 4.863382, 4.866856, 
    4.868075, 4.867185, 4.864679, 4.861393, 4.858432, 4.857043, 4.85846, 
    4.863751,
  // totalHeight(17,3, 0-49)
    4.924704, 4.905055, 4.888456, 4.875116, 4.865107, 4.858351, 4.854629, 
    4.85358, 4.85474, 4.85757, 4.861506, 4.865989, 4.870497, 4.874556, 
    4.877724, 4.879621, 4.88518, 4.884454, 4.882708, 4.879936, 4.876042, 
    4.872316, 4.867249, 4.861258, 4.854124, 4.846151, 4.837596, 4.828926, 
    4.820539, 4.813347, 4.807551, 4.805, 4.804668, 4.806671, 4.810932, 
    4.817171, 4.824917, 4.833555, 4.842372, 4.850632, 4.85764, 4.862832, 
    4.865854, 4.866643, 4.865483, 4.863023, 4.860238, 4.858329, 4.858582, 
    4.862187,
  // totalHeight(17,4, 0-49)
    4.925554, 4.906652, 4.890803, 4.878195, 4.868879, 4.862763, 4.859605, 
    4.859044, 4.860619, 4.863809, 4.868073, 4.87288, 4.877728, 4.882148, 
    4.885689, 4.887709, 4.894379, 4.894003, 4.892564, 4.890065, 4.886366, 
    4.88302, 4.878093, 4.872019, 4.8645, 4.855797, 4.846127, 4.835956, 
    4.825689, 4.816328, 4.808094, 4.803315, 4.800786, 4.800761, 4.803308, 
    4.808267, 4.815266, 4.823757, 4.833058, 4.842415, 4.85107, 4.858335, 
    4.863684, 4.866829, 4.867804, 4.867007, 4.865207, 4.863475, 4.863067, 
    4.865251,
  // totalHeight(17,5, 0-49)
    4.926895, 4.908814, 4.893754, 4.881882, 4.873228, 4.86768, 4.86499, 
    4.864796, 4.866652, 4.870066, 4.874532, 4.879558, 4.884674, 4.889433, 
    4.893384, 4.89547, 4.903042, 4.903224, 4.902287, 4.900254, 4.896966, 
    4.894212, 4.889642, 4.883701, 4.87602, 4.866802, 4.856206, 4.844675, 
    4.832611, 4.821059, 4.810258, 4.803021, 4.79799, 4.795586, 4.796041, 
    4.799346, 4.805257, 4.813318, 4.822897, 4.833249, 4.843571, 4.853073, 
    4.861067, 4.867047, 4.870778, 4.872372, 4.872322, 4.871489, 4.871013, 
    4.872166,
  // totalHeight(17,6, 0-49)
    4.928093, 4.910898, 4.896666, 4.885541, 4.877535, 4.872518, 4.870237, 
    4.870338, 4.872396, 4.875957, 4.880558, 4.885754, 4.891115, 4.89623, 
    4.900664, 4.902766, 4.910966, 4.911911, 4.911652, 4.910261, 4.907574, 
    4.905591, 4.901582, 4.895983, 4.888383, 4.878903, 4.867634, 4.85497, 
    4.841294, 4.827643, 4.814258, 4.804423, 4.796666, 4.791592, 4.789618, 
    4.790914, 4.795382, 4.802684, 4.812258, 4.823384, 4.835237, 4.84695, 
    4.857692, 4.866757, 4.873649, 4.878177, 4.88052, 4.881258, 4.881336, 
    4.881945,
  // totalHeight(17,7, 0-49)
    4.928635, 4.912382, 4.89902, 4.888669, 4.88132, 4.87683, 4.874942, 
    4.875315, 4.877554, 4.88124, 4.88596, 4.891318, 4.896939, 4.902454, 
    4.907468, 4.909537, 4.918041, 4.919922, 4.920493, 4.919884, 4.91795, 
    4.916876, 4.913595, 4.908529, 4.901253, 4.891789, 4.880151, 4.866659, 
    4.851659, 4.836112, 4.820251, 4.80779, 4.797184, 4.789228, 4.78455, 
    4.783514, 4.786196, 4.792386, 4.801616, 4.813207, 4.826326, 4.840052, 
    4.853444, 4.865614, 4.875832, 4.883608, 4.8888, 4.891662, 4.892874, 
    4.893465,
  // totalHeight(17,8, 0-49)
    4.928143, 4.912886, 4.900441, 4.890904, 4.884245, 4.880311, 4.878841, 
    4.87951, 4.88195, 4.885783, 4.890644, 4.89619, 4.902103, 4.908071, 
    4.913764, 4.915773, 4.92422, 4.927168, 4.928677, 4.928949, 4.927879, 
    4.927794, 4.925365, 4.920992, 4.914267, 4.905104, 4.893435, 4.879482, 
    4.863534, 4.846408, 4.828302, 4.813304, 4.799834, 4.788882, 4.781299, 
    4.777662, 4.778239, 4.782969, 4.791487, 4.803172, 4.817198, 4.83261, 
    4.848373, 4.863461, 4.876935, 4.88804, 4.896313, 4.901678, 4.904503, 
    4.905589,
  // totalHeight(17,9, 0-49)
    4.926387, 4.91217, 4.900692, 4.892024, 4.88611, 4.882786, 4.881791, 
    4.882813, 4.88551, 4.889541, 4.894586, 4.900361, 4.906602, 4.913068, 
    4.919524, 4.921489, 4.929521, 4.933596, 4.936105, 4.937315, 4.937177, 
    4.938101, 4.936598, 4.933035, 4.927056, 4.918464, 4.90711, 4.893102, 
    4.876647, 4.85835, 4.838352, 4.821018, 4.804783, 4.790828, 4.780226, 
    4.773788, 4.771987, 4.774931, 4.782368, 4.793742, 4.808257, 4.824928, 
    4.84266, 4.860311, 4.876772, 4.891061, 4.902427, 4.910475, 4.915247, 
    4.917273,
  // totalHeight(17,10, 0-49)
    4.923273, 4.910128, 4.899665, 4.891922, 4.886822, 4.884184, 4.883743, 
    4.885196, 4.888224, 4.892519, 4.897807, 4.903848, 4.910443, 4.917434, 
    4.924696, 4.92671, 4.934017, 4.939202, 4.942721, 4.944888, 4.945706, 
    4.947608, 4.947049, 4.944363, 4.939278, 4.931495, 4.920787, 4.907132, 
    4.890639, 4.871647, 4.850207, 4.83084, 4.812048, 4.795187, 4.781552, 
    4.772192, 4.767801, 4.768667, 4.774671, 4.785334, 4.799887, 4.817338, 
    4.836549, 4.856289, 4.875316, 4.892464, 4.906739, 4.917458, 4.924351, 
    4.92766,
  // totalHeight(17,11, 0-49)
    4.918819, 4.906762, 4.897353, 4.890594, 4.886381, 4.884509, 4.884711, 
    4.886684, 4.890129, 4.89476, 4.90034, 4.906679, 4.913639, 4.921144, 
    4.929193, 4.931473, 4.937835, 4.944029, 4.948521, 4.951626, 4.953395, 
    4.95619, 4.956545, 4.954758, 4.950663, 4.943872, 4.934094, 4.921172, 
    4.905105, 4.885919, 4.863553, 4.842531, 4.821484, 4.801915, 4.785327, 
    4.773007, 4.765884, 4.764438, 4.768693, 4.778259, 4.792406, 4.810146, 
    4.830305, 4.851591, 4.872667, 4.89222, 4.909069, 4.922284, 4.931321, 
    4.936136,
  // totalHeight(17,12, 0-49)
    4.913151, 4.902174, 4.89384, 4.888111, 4.884847, 4.883822, 4.884756, 
    4.887339, 4.891278, 4.896312, 4.90223, 4.908882, 4.91619, 4.924158, 
    4.932895, 4.935816, 4.941145, 4.948177, 4.953555, 4.957557, 4.960253, 
    4.96382, 4.965019, 4.964102, 4.961035, 4.955356, 4.946728, 4.934856, 
    4.919626, 4.900735, 4.877989, 4.855725, 4.832791, 4.810797, 4.791426, 
    4.776199, 4.766277, 4.762349, 4.764593, 4.772719, 4.786045, 4.803592, 
    4.82417, 4.846443, 4.869005, 4.890441, 4.90943, 4.924849, 4.935921, 
    4.942349,
  // totalHeight(17,13, 0-49)
    4.906466, 4.896542, 4.889278, 4.884605, 4.882339, 4.882226, 4.883963, 
    4.887234, 4.891738, 4.897228, 4.903514, 4.91048, 4.918095, 4.926425, 
    4.93566, 4.939777, 4.944144, 4.951789, 4.95794, 4.962779, 4.966364, 
    4.970561, 4.972504, 4.972393, 4.970335, 4.96582, 4.958477, 4.947888, 
    4.933827, 4.915659, 4.893061, 4.869974, 4.845552, 4.821473, 4.799566, 
    4.781562, 4.768855, 4.762346, 4.762383, 4.768782, 4.78092, 4.797838, 
    4.818337, 4.841057, 4.864547, 4.887329, 4.907979, 4.925239, 4.938151, 
    4.946199,
  // totalHeight(17,14, 0-49)
    4.899024, 4.89009, 4.883871, 4.880249, 4.879004, 4.879846, 4.882438, 
    4.886447, 4.891568, 4.897552, 4.90422, 4.911483, 4.919337, 4.927886, 
    4.937351, 4.943377, 4.947018, 4.955034, 4.961828, 4.967443, 4.971882, 
    4.976558, 4.979132, 4.979733, 4.97862, 4.975255, 4.969245, 4.960069, 
    4.947399, 4.930287, 4.908312, 4.884778, 4.859268, 4.833473, 4.809331, 
    4.788751, 4.773347, 4.764234, 4.761935, 4.766388, 4.777039, 4.792955, 
    4.812939, 4.835619, 4.859524, 4.883137, 4.904978, 4.923697, 4.9382, 
    4.947796,
  // totalHeight(17,15, 0-49)
    4.891112, 4.883087, 4.877852, 4.875248, 4.875012, 4.876813, 4.880279, 
    4.885053, 4.890813, 4.897305, 4.904356, 4.911882, 4.919893, 4.928493, 
    4.93788, 4.946609, 4.949912, 4.958069, 4.965397, 4.97174, 4.97701, 
    4.982026, 4.985116, 4.986323, 4.986053, 4.983757, 4.979042, 4.971297, 
    4.960118, 4.944283, 4.923313, 4.899639, 4.873401, 4.84626, 4.820212, 
    4.797309, 4.779364, 4.767699, 4.763014, 4.76538, 4.774317, 4.788934, 
    4.808044, 4.830278, 4.854156, 4.87815, 4.900752, 4.920557, 4.936386, 
    4.947409,
  // totalHeight(17,16, 0-49)
    4.883029, 4.875806, 4.871468, 4.869812, 4.870532, 4.873254, 4.877571, 
    4.883094, 4.889482, 4.896476, 4.903892, 4.911646, 4.919736, 4.928235, 
    4.937255, 4.949426, 4.952873, 4.96102, 4.968817, 4.975876, 4.981983, 
    4.987225, 4.990734, 4.992444, 4.992887, 4.991526, 4.987975, 4.981569, 
    4.971848, 4.957378, 4.937684, 4.914083, 4.887414, 4.859268, 4.831649, 
    4.806712, 4.786437, 4.772339, 4.765296, 4.765512, 4.772596, 4.785703, 
    4.803671, 4.825141, 4.84864, 4.872643, 4.89564, 4.916207, 4.933103, 
    4.945402,
  // totalHeight(17,17, 0-49)
    4.875055, 4.868514, 4.864955, 4.864135, 4.86571, 4.869261, 4.87435, 
    4.880558, 4.88753, 4.89499, 4.902754, 4.910722, 4.918859, 4.927171, 
    4.935653, 4.951737, 4.955822, 4.963933, 4.972224, 4.980051, 4.987048, 
    4.992446, 4.996313, 4.998434, 4.999444, 4.99883, 4.99623, 4.990953, 
    4.982525, 4.969369, 4.951089, 4.927674, 4.900793, 4.871935, 4.843071, 
    4.816412, 4.794065, 4.777717, 4.768412, 4.766494, 4.771667, 4.783143, 
    4.799794, 4.820279, 4.843141, 4.866875, 4.889984, 4.911039, 4.928771, 
    4.942188,
  // totalHeight(17,18, 0-49)
    4.867438, 4.861432, 4.858498, 4.858359, 4.860627, 4.864854, 4.870573, 
    4.87735, 4.884819, 4.892704, 4.900818, 4.909043, 4.917301, 4.925497, 
    4.93346, 4.953443, 4.958536, 4.966762, 4.975693, 4.984436, 4.992451, 
    4.997995, 5.002215, 5.004687, 5.006111, 5.006001, 5.004041, 4.999564, 
    4.992125, 4.980086, 4.963223, 4.940009, 4.913056, 4.88373, 4.853928, 
    4.825867, 4.801744, 4.783382, 4.771981, 4.768018, 4.771304, 4.781112, 
    4.796357, 4.815728, 4.83779, 4.861065, 4.884079, 4.905415, 4.923792, 
    4.938173,
  // totalHeight(17,19, 0-49)
    4.860362, 4.854715, 4.852209, 4.85253, 4.855262, 4.859932, 4.866065, 
    4.87323, 4.881079, 4.889356, 4.89789, 4.906549, 4.915184, 4.923564, 
    4.931289, 4.954461, 4.960647, 4.969331, 4.979218, 4.989158, 4.998429, 
    5.004205, 5.008854, 5.011667, 5.013352, 5.01345, 5.011711, 5.007554, 
    5.000636, 4.989366, 4.973771, 4.950686, 4.92374, 4.894152, 4.863704, 
    4.834578, 4.809007, 4.788918, 4.775646, 4.769795, 4.771284, 4.77946, 
    4.793291, 4.811497, 4.83268, 4.855388, 4.878173, 4.899641, 4.918513, 
    4.933718,
  // totalHeight(17,20, 0-49)
    4.854655, 4.849918, 4.84861, 4.850455, 4.855026, 4.861779, 4.870096, 
    4.879328, 4.888843, 4.898059, 4.906477, 4.913717, 4.919533, 4.923843, 
    4.926725, 30, 4.976701, 4.980468, 4.985542, 4.99134, 4.997496, 5.000072, 
    5.003079, 5.005518, 5.008004, 5.009818, 5.010391, 5.008807, 5.004483, 
    4.995662, 4.982596, 4.960472, 4.934066, 4.904542, 4.873656, 4.843603, 
    4.816685, 4.794946, 4.779853, 4.772143, 4.771838, 4.778371, 4.790754, 
    4.807751, 4.827991, 4.850053, 4.872515, 4.894001, 4.913239, 4.929135,
  // totalHeight(17,21, 0-49)
    4.849359, 4.844958, 4.844018, 4.846222, 4.851108, 4.858102, 4.866564, 
    4.875849, 4.885345, 4.89451, 4.90289, 4.910137, 4.916014, 4.920402, 
    4.923314, 30, 4.978804, 4.983113, 4.98882, 4.995245, 5.001908, 5.003341, 
    5.005481, 5.007151, 5.009163, 5.010862, 5.011708, 5.010763, 5.007414, 
    4.999859, 4.988595, 4.967202, 4.941577, 4.912706, 4.882171, 4.852049, 
    4.824604, 4.801916, 4.785548, 4.776368, 4.774518, 4.77953, 4.790494, 
    4.806223, 4.825388, 4.846598, 4.868461, 4.889622, 4.908823, 4.924966,
  // totalHeight(17,22, 0-49)
    4.84491, 4.840719, 4.840024, 4.842488, 4.847629, 4.854852, 4.863504, 
    4.872935, 4.882536, 4.891777, 4.900223, 4.907533, 4.913461, 4.917856, 
    4.920673, 30, 4.980448, 4.985187, 4.991485, 4.998569, 5.005846, 5.006361, 
    5.007894, 5.009054, 5.010793, 5.012468, 5.013533, 5.01302, 5.010294, 
    5.003533, 4.9935, 4.972336, 4.947056, 4.918531, 4.888209, 4.858057, 
    4.830273, 4.806931, 4.789643, 4.779356, 4.776308, 4.780115, 4.789931, 
    4.804622, 4.822892, 4.843383, 4.864727, 4.885594, 4.904738, 4.921063,
  // totalHeight(17,23, 0-49)
    4.841343, 4.837268, 4.836722, 4.839362, 4.844692, 4.852111, 4.860959, 
    4.870574, 4.880348, 4.889748, 4.898341, 4.905778, 4.911798, 4.916217, 
    4.918941, 30, 4.982242, 4.987259, 4.993968, 5.001531, 5.009266, 5.00898, 
    5.009981, 5.010692, 5.012161, 5.013753, 5.014909, 5.014637, 5.012286, 
    5.006017, 4.996813, 4.975653, 4.950515, 4.922195, 4.892049, 4.861947, 
    4.834018, 4.810307, 4.792441, 4.781416, 4.77753, 4.780464, 4.789426, 
    4.803322, 4.820889, 4.840794, 4.86169, 4.882262, 4.901279, 4.917653,
  // totalHeight(17,24, 0-49)
    4.838642, 4.834622, 4.834155, 4.836901, 4.842365, 4.849943, 4.858972, 
    4.868788, 4.878774, 4.888392, 4.897195, 4.904826, 4.911006, 4.915524, 
    4.918251, 30, 4.984415, 4.98959, 4.996536, 5.004384, 5.012406, 5.011586, 
    5.012234, 5.012639, 5.013902, 5.015387, 5.016535, 5.016338, 5.014139, 
    5.008089, 4.999325, 4.978053, 4.952898, 4.924624, 4.894527, 4.864416, 
    4.836373, 4.812413, 4.794162, 4.782639, 4.778178, 4.7805, 4.788852, 
    4.80217, 4.819218, 4.838678, 4.859221, 4.879544, 4.898427, 4.914783,
  // totalHeight(17,25, 0-49)
    4.836769, 4.832759, 4.832325, 4.83513, 4.840688, 4.8484, 4.857604, 
    4.867634, 4.877865, 4.887749, 4.896824, 4.904718, 4.911138, 4.915858, 
    4.918736, 30, 4.986551, 4.991792, 4.998822, 5.006766, 5.014881, 5.013883, 
    5.014416, 5.014708, 5.015873, 5.017272, 5.018345, 5.018085, 5.015834, 
    5.009744, 5.001011, 4.979569, 4.954289, 4.925926, 4.895759, 4.865575, 
    4.83743, 4.813322, 4.794866, 4.783079, 4.778309, 4.780292, 4.788291, 
    4.801262, 4.817979, 4.837139, 4.85742, 4.877531, 4.89625, 4.912501,
  // totalHeight(17,26, 0-49)
    4.835672, 4.83165, 4.831218, 4.834058, 4.839693, 4.847535, 4.856926, 
    4.867199, 4.877722, 4.887929, 4.897342, 4.905571, 4.912312, 4.917341, 
    4.920526, 30, 4.988527, 4.993752, 5.000716, 5.008561, 5.016568, 5.015782, 
    5.016457, 5.016857, 5.018059, 5.019417, 5.020375, 5.019933, 5.017445, 
    5.011068, 5.001957, 4.980327, 4.954838, 4.92627, 4.895921, 4.865594, 
    4.837351, 4.813177, 4.794672, 4.782838, 4.778008, 4.779906, 4.787796, 
    4.800632, 4.817194, 4.836185, 4.856286, 4.876206, 4.894732, 4.910787,
  // totalHeight(17,27, 0-49)
    4.835305, 4.831254, 4.830816, 4.833688, 4.83941, 4.847407, 4.857031, 
    4.86761, 4.878496, 4.889104, 4.898934, 4.907572, 4.914705, 4.920119, 
    4.923718, 30, 4.990418, 4.995515, 5.002238, 5.00977, 5.01746, 5.017213, 
    5.018252, 5.01895, 5.020303, 5.021653, 5.022446, 5.021699, 5.018786, 
    5.011879, 5.002003, 4.980161, 4.954391, 4.925523, 4.894915, 4.864421, 
    4.836125, 4.812012, 4.793656, 4.782018, 4.777392, 4.779467, 4.787487, 
    4.800394, 4.816962, 4.835893, 4.855869, 4.875599, 4.893869, 4.909608,
  // totalHeight(17,28, 0-49)
    4.835628, 4.831538, 4.831094, 4.834014, 4.839862, 4.848079, 4.85802, 
    4.869009, 4.880377, 4.891504, 4.90185, 4.910967, 4.91853, 4.924347, 
    4.928369, 30, 4.992599, 4.997404, 5.003668, 5.010651, 5.017807, 5.018314, 
    5.019859, 5.020988, 5.022568, 5.023917, 5.02448, 5.023301, 5.019778, 
    5.01211, 5.00112, 4.979014, 4.952876, 4.923621, 4.892708, 4.862062, 
    4.833807, 4.809922, 4.791938, 4.780753, 4.776589, 4.779086, 4.787449, 
    4.8006, 4.817302, 4.836254, 4.856133, 4.875648, 4.893589, 4.908889,
  // totalHeight(17,29, 0-49)
    4.836607, 4.832465, 4.832018, 4.835017, 4.841056, 4.849597, 4.859998, 
    4.871566, 4.883592, 4.8954, 4.906381, 4.916035, 4.924014, 4.930147, 
    4.934448, 30, 4.994762, 4.999057, 5.004619, 5.010811, 5.01722, 5.01852, 
    5.020604, 5.022212, 5.02405, 5.025388, 5.025658, 5.023925, 5.019612, 
    5.010951, 4.998516, 4.976011, 4.949397, 4.919718, 4.888555, 4.857924, 
    4.829979, 4.806665, 4.789436, 4.779088, 4.77575, 4.778986, 4.787952, 
    4.80154, 4.818505, 4.837532, 4.857296, 4.876508, 4.89396, 4.908601,
  // totalHeight(17,30, 0-49)
    4.837832, 4.833149, 4.831962, 4.833973, 4.838768, 4.84586, 4.854743, 
    4.86493, 4.875998, 4.887613, 4.899509, 4.911485, 4.923332, 4.93478, 
    4.945404, 4.975517, 4.979926, 4.9902, 5.001615, 5.01291, 5.023316, 
    5.028723, 5.033325, 5.036073, 5.037669, 5.037555, 5.035443, 5.030748, 
    5.023216, 5.011344, 4.995587, 4.971336, 4.943355, 4.912786, 4.881282, 
    4.850867, 4.823629, 4.801392, 4.785451, 4.776451, 4.77439, 4.778745, 
    4.788615, 4.802867, 4.820241, 4.839418, 4.859073, 4.87792, 4.894762, 
    4.908581,
  // totalHeight(17,31, 0-49)
    4.840512, 4.836057, 4.835127, 4.837435, 4.842564, 4.85002, 4.85927, 
    4.869801, 4.881155, 4.892956, 4.904926, 4.916868, 4.928643, 4.940125, 
    4.951134, 4.976396, 4.981072, 4.990958, 5.001443, 5.011515, 5.020609, 
    5.025819, 5.029953, 5.032291, 5.033554, 5.033181, 5.03083, 5.025838, 
    5.017842, 5.005279, 4.988306, 4.964038, 4.936157, 4.905926, 4.875092, 
    4.845701, 4.81979, 4.799075, 4.784719, 4.777233, 4.77651, 4.781954, 
    4.792624, 4.80736, 4.824892, 4.843892, 4.863036, 4.881039, 4.896733, 
    4.90915,
  // totalHeight(17,32, 0-49)
    4.84394, 4.839687, 4.838961, 4.84147, 4.8468, 4.854445, 4.863869, 
    4.874544, 4.886004, 4.897867, 4.909857, 4.921802, 4.933619, 4.9453, 
    4.956847, 4.976905, 4.981479, 4.991234, 5.00101, 5.010061, 5.018018, 
    5.023118, 5.026866, 5.028792, 5.02958, 5.028664, 5.025671, 5.019921, 
    5.011018, 4.997434, 4.979104, 4.954812, 4.927166, 4.897542, 4.867736, 
    4.839773, 4.815597, 4.796778, 4.784322, 4.7786, 4.779403, 4.786065, 
    4.797607, 4.812852, 4.830517, 4.849267, 4.867775, 4.88477, 4.899115, 
    4.909908,
  // totalHeight(17,33, 0-49)
    4.848188, 4.844136, 4.843581, 4.846228, 4.851653, 4.859349, 4.868777, 
    4.879411, 4.890791, 4.902544, 4.914413, 4.926251, 4.938032, 4.949833, 
    4.961806, 4.976944, 4.981427, 4.991122, 5.000261, 5.008378, 5.015282, 
    5.02028, 5.023657, 5.025142, 5.025333, 5.023657, 5.019734, 5.012911, 
    5.002809, 4.988014, 4.968327, 4.944061, 4.916827, 4.88808, 4.859641, 
    4.83347, 4.811376, 4.794761, 4.784458, 4.780696, 4.783165, 4.791138, 
    4.803601, 4.819355, 4.837107, 4.855516, 4.87325, 4.889057, 4.901842, 
    4.910791,
  // totalHeight(17,34, 0-49)
    4.853289, 4.849438, 4.849027, 4.851749, 4.857172, 4.864788, 4.874062, 
    4.88448, 4.895594, 4.907053, 4.91862, 4.930174, 4.941731, 4.953428, 
    4.965522, 4.976438, 4.981064, 4.990592, 4.999053, 5.006239, 5.012118, 
    5.01695, 5.019924, 5.020919, 5.020409, 5.017825, 5.01279, 5.004707, 
    4.993249, 4.9772, 4.956297, 4.932189, 4.905595, 4.878024, 4.85128, 
    4.827223, 4.8075, 4.793324, 4.785354, 4.783679, 4.787896, 4.797219, 
    4.810601, 4.826828, 4.844588, 4.862535, 4.879337, 4.893764, 4.904784, 
    4.911689,
  // totalHeight(17,35, 0-49)
    4.859222, 4.855562, 4.855252, 4.857974, 4.863289, 4.870693, 4.879658, 
    4.889689, 4.900362, 4.911344, 4.922421, 4.933497, 4.944608, 4.955915, 
    4.967728, 4.975316, 4.980386, 4.989532, 4.997201, 5.003416, 5.00826, 
    5.012824, 5.015333, 5.015789, 5.014503, 5.010921, 5.004682, 4.995273, 
    4.982435, 4.965222, 4.943371, 4.919636, 4.893962, 4.867884, 4.843148, 
    4.82148, 4.804347, 4.792766, 4.787225, 4.787683, 4.793653, 4.804296, 
    4.81854, 4.835147, 4.852794, 4.870125, 4.885816, 4.898671, 4.907736, 
    4.912441,
  // totalHeight(17,36, 0-49)
    4.865902, 4.862398, 4.862123, 4.86475, 4.869839, 4.876892, 4.885399, 
    4.894885, 4.904952, 4.915292, 4.925711, 4.936127, 4.946576, 4.957216, 
    4.968345, 4.973502, 4.979285, 4.987776, 4.994511, 4.999691, 5.003481, 
    5.007654, 5.009626, 5.009497, 5.007393, 5.002791, 4.995346, 4.984653, 
    4.97054, 4.952381, 4.929957, 4.90688, 4.882451, 4.858187, 4.835741, 
    4.816682, 4.802279, 4.793364, 4.790259, 4.792812, 4.800456, 4.812315, 
    4.827287, 4.844121, 4.861478, 4.877997, 4.892375, 4.903469, 4.910425, 
    4.912837,
  // totalHeight(17,37, 0-49)
    4.873171, 4.869758, 4.869428, 4.871847, 4.876582, 4.883149, 4.891055, 
    4.899855, 4.909174, 4.918733, 4.928355, 4.93796, 4.947573, 4.957314, 
    4.967422, 4.970922, 4.977585, 4.98515, 4.990809, 4.994896, 4.997612, 
    5.001259, 5.002623, 5.001882, 4.998955, 4.993373, 4.984812, 4.972988, 
    4.957819, 4.939039, 4.916505, 4.894428, 4.871589, 4.849447, 4.829532, 
    4.813232, 4.801623, 4.795353, 4.794603, 4.799121, 4.808279, 4.821166, 
    4.836657, 4.853489, 4.870317, 4.885788, 4.898634, 4.907787, 4.91253, 
    4.912643,
  // totalHeight(17,38, 0-49)
    4.880799, 4.877385, 4.876884, 4.878968, 4.88322, 4.889169, 4.896352, 
    4.904349, 4.912816, 4.921493, 4.930215, 4.938902, 4.947552, 4.956231, 
    4.965086, 4.967517, 4.975098, 4.981501, 4.985966, 4.988914, 4.990543, 
    4.993541, 4.994239, 4.992883, 4.989176, 4.982718, 4.973215, 4.960507, 
    4.944603, 4.925617, 4.903484, 4.88278, 4.861875, 4.842131, 4.824929, 
    4.811468, 4.802634, 4.798907, 4.800348, 4.806618, 4.817043, 4.830686, 
    4.846407, 4.862938, 4.878937, 4.893082, 4.904164, 4.911223, 4.913716, 
    4.911637,
  // totalHeight(17,39, 0-49)
    4.8885, 4.884964, 4.884163, 4.885783, 4.889422, 4.894643, 4.901007, 
    4.908122, 4.915665, 4.923398, 4.931163, 4.938869, 4.946483, 4.95401, 
    4.961489, 4.963247, 4.971654, 4.976719, 4.979917, 4.981703, 4.982242, 
    4.984488, 4.984486, 4.982543, 4.978146, 4.970976, 4.960778, 4.947517, 
    4.931282, 4.912557, 4.891349, 4.872391, 4.853734, 4.836616, 4.822244, 
    4.811627, 4.805473, 4.804114, 4.807503, 4.815238, 4.826606, 4.840658, 
    4.856246, 4.87211, 4.886935, 4.899451, 4.908543, 4.913409, 4.913702, 
    4.909656,
  // totalHeight(17,40, 0-49)
    4.895968, 4.892166, 4.890924, 4.891946, 4.894863, 4.899263, 4.90474, 
    4.910928, 4.917522, 4.924296, 4.931087, 4.937795, 4.944351, 4.950702, 
    4.956784, 4.958094, 4.967124, 4.970757, 4.972659, 4.973285, 4.972751, 
    4.974173, 4.973469, 4.971002, 4.966048, 4.958385, 4.947799, 4.934374, 
    4.918255, 4.900277, 4.880496, 4.863629, 4.847486, 4.833153, 4.821659, 
    4.813825, 4.810189, 4.810955, 4.815989, 4.824837, 4.836764, 4.850812, 
    4.865849, 4.880637, 4.893913, 4.904496, 4.911415, 4.914057, 4.912313, 
    4.906664,
  // totalHeight(17,41, 0-49)
    4.902921, 4.898695, 4.89686, 4.897158, 4.899249, 4.902759, 4.907311, 
    4.91256, 4.918214, 4.924046, 4.929891, 4.935626, 4.941149, 4.946351, 
    4.951089, 4.952054, 4.96143, 4.963621, 4.964247, 4.963741, 4.962173, 
    4.962739, 4.96137, 4.958476, 4.95314, 4.945245, 4.934614, 4.921438, 
    4.905893, 4.88913, 4.871221, 4.856738, 4.843309, 4.831854, 4.823215, 
    4.818036, 4.816703, 4.819304, 4.825633, 4.835196, 4.847248, 4.860843, 
    4.874875, 4.888161, 4.899525, 4.907917, 4.912551, 4.913051, 4.909559, 
    4.9028,
  // totalHeight(17,42, 0-49)
    4.909159, 4.904336, 4.901761, 4.901208, 4.902383, 4.904947, 4.90855, 
    4.912868, 4.917612, 4.922549, 4.9275, 4.932313, 4.936859, 4.940983, 
    4.944482, 4.945125, 4.954541, 4.955351, 4.954765, 4.953189, 4.95065, 
    4.950379, 4.948419, 4.945224, 4.939711, 4.931865, 4.921547, 4.909028, 
    4.894497, 4.879364, 4.863691, 4.851813, 4.841222, 4.832664, 4.826799, 
    4.8241, 4.824811, 4.828923, 4.836165, 4.846019, 4.857746, 4.870423, 
    4.883003, 4.894386, 4.903529, 4.90956, 4.911921, 4.910494, 4.905684, 
    4.898421,
  // totalHeight(17,43, 0-49)
    4.914628, 4.909033, 4.905563, 4.904037, 4.904203, 4.905764, 4.908397, 
    4.91179, 4.915656, 4.919752, 4.923867, 4.927831, 4.931473, 4.934608, 
    4.936998, 4.937302, 4.946457, 4.946009, 4.944318, 4.94176, 4.938349, 
    4.937307, 4.934862, 4.93152, 4.926051, 4.91854, 4.908878, 4.897394, 
    4.884263, 4.871099, 4.857931, 4.848797, 4.84109, 4.835384, 4.832156, 
    4.83172, 4.834194, 4.839475, 4.847241, 4.856964, 4.867921, 4.879242, 
    4.889966, 4.899126, 4.905847, 4.909483, 4.909735, 4.906756, 4.901185, 
    4.894104,
  // totalHeight(17,44, 0-49)
    4.919461, 4.912925, 4.908408, 4.905779, 4.904836, 4.90532, 4.90694, 
    4.909394, 4.912395, 4.915678, 4.919009, 4.92218, 4.924991, 4.92723, 
    4.928645, 4.928577, 4.937214, 4.935669, 4.933005, 4.929586, 4.925431, 
    4.923725, 4.920937, 4.917611, 4.91241, 4.905505, 4.896807, 4.88668, 
    4.875265, 4.864319, 4.85382, 4.847488, 4.84264, 4.839678, 4.838911, 
    4.8405, 4.844442, 4.850554, 4.858476, 4.867672, 4.877462, 4.887057, 
    4.895621, 4.902356, 4.906611, 4.907991, 4.906475, 4.902468, 4.896797, 
    4.890616,
  // totalHeight(17,45, 0-49)
    4.924008, 4.916375, 4.910664, 4.906796, 4.904622, 4.903929, 4.904456, 
    4.905918, 4.908018, 4.910478, 4.913033, 4.91544, 4.91747, 4.918889, 
    4.919441, 4.918964, 4.926886, 4.924419, 4.920935, 4.916797, 4.912052, 
    4.909824, 4.906849, 4.903707, 4.898986, 4.892923, 4.885447, 4.876929, 
    4.86746, 4.858889, 4.851131, 4.847575, 4.845493, 4.84512, 4.846608, 
    4.849974, 4.855102, 4.861737, 4.869482, 4.877822, 4.886137, 4.893749, 
    4.899987, 4.904269, 4.906194, 4.90565, 4.902875, 4.898486, 4.893424, 
    4.888831,
  // totalHeight(17,46, 0-49)
    4.928825, 4.919962, 4.912918, 4.90767, 4.904126, 4.902122, 4.90143, 
    4.901784, 4.902892, 4.904456, 4.906185, 4.907807, 4.909061, 4.909698, 
    4.909465, 4.908536, 4.915604, 4.912388, 4.908238, 4.903537, 4.898368, 
    4.895784, 4.892784, 4.88998, 4.885921, 4.880892, 4.874827, 4.868092, 
    4.860718, 4.854588, 4.849548, 4.848677, 4.849215, 4.851243, 4.854764, 
    4.859663, 4.865725, 4.87262, 4.879941, 4.887194, 4.89385, 4.899375, 
    4.903301, 4.905291, 4.905223, 4.903256, 4.899861, 4.895799, 4.892039, 
    4.889628,
  // totalHeight(17,47, 0-49)
    4.934628, 4.924436, 4.915936, 4.909171, 4.904103, 4.900622, 4.898542, 
    4.897622, 4.897577, 4.898103, 4.89889, 4.899638, 4.900064, 4.899903, 
    4.898912, 4.897471, 4.903601, 4.899779, 4.895105, 4.889996, 4.884573, 
    4.881795, 4.878922, 4.876583, 4.873326, 4.869465, 4.864933, 4.860072, 
    4.85486, 4.851156, 4.848743, 4.850405, 4.853375, 4.857594, 4.862926, 
    4.869143, 4.875928, 4.882905, 4.889649, 4.895721, 4.900694, 4.904212, 
    4.906034, 4.906089, 4.904534, 4.901772, 4.898455, 4.895413, 4.893567, 
    4.893793,
  // totalHeight(17,48, 0-49)
    4.942206, 4.930628, 4.920584, 4.912177, 4.905432, 4.900293, 4.896624, 
    4.894217, 4.892807, 4.892093, 4.891754, 4.891472, 4.890954, 4.889923, 
    4.888144, 4.886106, 4.891249, 4.886915, 4.881835, 4.876449, 4.870919, 
    4.868098, 4.865475, 4.863686, 4.861314, 4.858688, 4.855734, 4.852766, 
    4.84971, 4.848352, 4.848417, 4.852421, 4.857611, 4.863803, 4.870745, 
    4.878098, 4.885471, 4.89244, 4.898585, 4.903532, 4.906981, 4.908762, 
    4.908873, 4.907512, 4.905091, 4.902219, 4.899659, 4.898243, 4.898774, 
    4.901918,
  // totalHeight(17,49, 0-49)
    4.959617, 4.946238, 4.934052, 4.923233, 4.913883, 4.906022, 4.89959, 
    4.894449, 4.890389, 4.887144, 4.884412, 4.881876, 4.879222, 4.876143, 
    4.872361, 4.869101, 4.880398, 4.874001, 4.866947, 4.860031, 4.853502, 
    4.852767, 4.852791, 4.85458, 4.855067, 4.854731, 4.853221, 4.850918, 
    4.847435, 4.846223, 4.846673, 4.853611, 4.861576, 4.870242, 4.879228, 
    4.888075, 4.896299, 4.903437, 4.909089, 4.912979, 4.914989, 4.915207, 
    4.913942, 4.911713, 4.909215, 4.907247, 4.906631, 4.908108, 4.91226, 
    4.919442,
  // totalHeight(18,0, 0-49)
    4.884809, 4.871144, 4.860725, 4.853534, 4.849423, 4.848121, 4.849251, 
    4.852354, 4.856926, 4.862458, 4.868456, 4.874484, 4.880164, 4.885192, 
    4.88933, 4.892411, 4.895638, 4.896484, 4.896322, 4.895182, 4.893073, 
    4.890365, 4.886718, 4.882278, 4.87701, 4.871042, 4.864499, 4.857598, 
    4.850573, 4.843819, 4.837571, 4.832456, 4.82845, 4.825788, 4.824625, 
    4.825011, 4.826875, 4.830015, 4.834108, 4.838731, 4.843399, 4.84762, 
    4.850959, 4.853108, 4.853957, 4.853652, 4.852622, 4.851551, 4.851324, 
    4.852911,
  // totalHeight(18,1, 0-49)
    4.884934, 4.871832, 4.862022, 4.855465, 4.85199, 4.851309, 4.853025, 
    4.856676, 4.861752, 4.867746, 4.874176, 4.880609, 4.886672, 4.892051, 
    4.896487, 4.899747, 4.904272, 4.905182, 4.905079, 4.903979, 4.901849, 
    4.899334, 4.895684, 4.891092, 4.885404, 4.878729, 4.871161, 4.862932, 
    4.854278, 4.845744, 4.837555, 4.830768, 4.825129, 4.820971, 4.818543, 
    4.817976, 4.819256, 4.822213, 4.826527, 4.831753, 4.837351, 4.842746, 
    4.847396, 4.850862, 4.852898, 4.853511, 4.853005, 4.851987, 4.851309, 
    4.851967,
  // totalHeight(18,2, 0-49)
    4.886409, 4.873914, 4.864717, 4.858756, 4.855839, 4.85566, 4.857812, 
    4.861832, 4.867219, 4.87348, 4.880151, 4.886819, 4.893123, 4.898752, 
    4.903427, 4.906798, 4.912543, 4.913613, 4.913682, 4.912762, 4.910775, 
    4.908639, 4.905188, 4.900646, 4.894743, 4.887562, 4.879149, 4.869736, 
    4.859549, 4.849249, 4.839058, 4.830468, 4.823002, 4.817106, 4.813138, 
    4.811329, 4.811743, 4.814265, 4.818604, 4.82431, 4.830813, 4.837478, 
    4.84367, 4.848833, 4.852573, 4.854734, 4.855453, 4.855189, 4.854686, 
    4.854899,
  // totalHeight(18,3, 0-49)
    4.888647, 4.876785, 4.868192, 4.862783, 4.86035, 4.860566, 4.863028, 
    4.867271, 4.872816, 4.879192, 4.885966, 4.892745, 4.899195, 4.905011, 
    4.909902, 4.913323, 4.920159, 4.921499, 4.921853, 4.921245, 4.919561, 
    4.917976, 4.914915, 4.910623, 4.904731, 4.897276, 4.888249, 4.877862, 
    4.866318, 4.854356, 4.842188, 4.831735, 4.822308, 4.814471, 4.808708, 
    4.805367, 4.804612, 4.806405, 4.810504, 4.816482, 4.823758, 4.831663, 
    4.839493, 4.846585, 4.852404, 4.856616, 4.859165, 4.860306, 4.860612, 
    4.860924,
  // totalHeight(18,4, 0-49)
    4.89114, 4.879928, 4.871926, 4.867028, 4.865009, 4.865537, 4.868205, 
    4.872565, 4.878159, 4.884547, 4.891326, 4.898142, 4.904681, 4.910653, 
    4.915773, 4.919184, 4.926921, 4.92865, 4.929398, 4.929215, 4.927966, 
    4.927078, 4.924573, 4.920717, 4.91506, 4.907583, 4.898214, 4.887125, 
    4.874485, 4.861058, 4.847029, 4.834742, 4.823296, 4.813377, 4.805604, 
    4.800458, 4.798227, 4.798971, 4.802519, 4.808488, 4.816317, 4.825317, 
    4.834739, 4.843832, 4.851933, 4.858536, 4.863369, 4.866457, 4.868152, 
    4.869117,
  // totalHeight(18,5, 0-49)
    4.893487, 4.882936, 4.875515, 4.871094, 4.869439, 4.870214, 4.873019, 
    4.877421, 4.882993, 4.889328, 4.89606, 4.90287, 4.909472, 4.915598, 
    4.920979, 4.924315, 4.932712, 4.934937, 4.936172, 4.936502, 4.935794, 
    4.935705, 4.933889, 4.930626, 4.925414, 4.918171, 4.908759, 4.897293, 
    4.883885, 4.869284, 4.853611, 4.839611, 4.826176, 4.814109, 4.80417, 
    4.796988, 4.792989, 4.792358, 4.795018, 4.800653, 4.808738, 4.818592, 
    4.829433, 4.840447, 4.85086, 4.860002, 4.867395, 4.872821, 4.876379, 
    4.878513,
  // totalHeight(18,6, 0-49)
    4.895404, 4.88553, 4.878681, 4.874718, 4.873394, 4.874374, 4.877271, 
    4.881673, 4.887185, 4.893434, 4.900091, 4.906876, 4.913533, 4.919827, 
    4.925513, 4.928716, 4.937472, 4.940289, 4.942079, 4.942984, 4.942886, 
    4.94365, 4.942612, 4.940061, 4.935476, 4.928711, 4.919563, 4.908076, 
    4.894294, 4.878877, 4.861876, 4.846375, 4.831077, 4.816886, 4.8047, 
    4.795306, 4.789286, 4.78697, 4.788401, 4.79335, 4.801349, 4.811738, 
    4.823725, 4.836451, 4.849043, 4.860695, 4.870737, 4.878716, 4.884475, 
    4.888203,
  // totalHeight(18,7, 0-49)
    4.896717, 4.887537, 4.881267, 4.877753, 4.876744, 4.877908, 4.880875, 
    4.885259, 4.890693, 4.896843, 4.903419, 4.910171, 4.916884, 4.92336, 
    4.929397, 4.932419, 4.941206, 4.944678, 4.947065, 4.948576, 4.949125, 
    4.950751, 4.950533, 4.948766, 4.944954, 4.938883, 4.930294, 4.919146, 
    4.905412, 4.889598, 4.871658, 4.854958, 4.838015, 4.821816, 4.807391, 
    4.795682, 4.787444, 4.783171, 4.783046, 4.786955, 4.794499, 4.80506, 
    4.81785, 4.831971, 4.846484, 4.860461, 4.873067, 4.88364, 4.891777, 
    4.897409,
  // totalHeight(18,8, 0-49)
    4.897334, 4.888876, 4.8832, 4.880144, 4.879449, 4.880795, 4.88383, 
    4.888193, 4.893551, 4.899602, 4.906095, 4.912813, 4.919581, 4.926244, 
    4.932665, 4.935491, 4.943973, 4.948122, 4.951126, 4.953247, 4.954448, 
    4.956897, 4.957495, 4.956541, 4.953597, 4.948393, 4.940624, 4.930164, 
    4.916898, 4.901135, 4.882703, 4.865164, 4.846878, 4.828883, 4.812316, 
    4.798274, 4.78769, 4.78124, 4.779273, 4.781801, 4.788523, 4.798871, 
    4.812071, 4.82721, 4.843288, 4.859285, 4.874232, 4.887288, 4.897826, 
    4.905539,
  // totalHeight(18,9, 0-49)
    4.897227, 4.889523, 4.884467, 4.881888, 4.881528, 4.883073, 4.886189, 
    4.890546, 4.895837, 4.901796, 4.908204, 4.914883, 4.921696, 4.928542, 
    4.935356, 4.938022, 4.945889, 4.950691, 4.9543, 4.957017, 4.958854, 
    4.962049, 4.963417, 4.963258, 4.96123, 4.957014, 4.950277, 4.940805, 
    4.928404, 4.913132, 4.894676, 4.876698, 4.85743, 4.837928, 4.819408, 
    4.803104, 4.790129, 4.78135, 4.777303, 4.778151, 4.783701, 4.793451, 
    4.806657, 4.822395, 4.839628, 4.857264, 4.874227, 4.889527, 4.902359, 
    4.912195,
  // totalHeight(18,10, 0-49)
    4.896404, 4.88949, 4.885093, 4.883026, 4.883033, 4.884808, 4.888037, 
    4.892411, 4.897654, 4.903532, 4.909855, 4.916485, 4.923323, 4.930325, 
    4.937502, 4.940127, 4.947123, 4.952506, 4.956683, 4.959964, 4.962405, 
    4.966238, 4.968298, 4.968881, 4.967768, 4.964606, 4.959049, 4.950807, 
    4.939605, 4.925227, 4.90721, 4.889191, 4.869336, 4.848673, 4.828465, 
    4.810056, 4.79473, 4.783552, 4.777253, 4.776168, 4.780232, 4.789024, 
    4.80184, 4.817754, 4.835709, 4.854557, 4.873146, 4.890373, 4.905285, 
    4.917168,
  // totalHeight(18,11, 0-49)
    4.894901, 4.888815, 4.885118, 4.88361, 4.884029, 4.886082, 4.889462, 
    4.893889, 4.899112, 4.904922, 4.911164, 4.917727, 4.924558, 4.931664, 
    4.939128, 4.941932, 4.947885, 4.95373, 4.958413, 4.962218, 4.965225, 
    4.969569, 4.972219, 4.97346, 4.973217, 4.971121, 4.966827, 4.95998, 
    4.950234, 4.937087, 4.91993, 4.90224, 4.882188, 4.860743, 4.839166, 
    4.818886, 4.801331, 4.787762, 4.779115, 4.775909, 4.778225, 4.785737, 
    4.797791, 4.813478, 4.831725, 4.851353, 4.87115, 4.889936, 4.906639, 
    4.920398,
  // totalHeight(18,12, 0-49)
    4.892765, 4.88754, 4.884587, 4.88369, 4.884581, 4.886966, 4.890554, 
    4.89508, 4.900316, 4.906077, 4.912237, 4.918715, 4.925493, 4.932621, 
    4.940238, 4.94356, 4.948406, 4.954556, 4.959667, 4.963951, 4.967489, 
    4.972205, 4.97533, 4.977124, 4.977676, 4.976608, 4.973598, 4.968228, 
    4.960105, 4.94844, 4.9325, 4.915447, 4.895557, 4.873702, 4.851109, 
    4.829243, 4.809653, 4.793781, 4.782765, 4.777319, 4.777685, 4.783647, 
    4.794613, 4.809704, 4.827843, 4.847833, 4.868425, 4.888381, 4.906549, 
    4.921947,
  // totalHeight(18,13, 0-49)
    4.890054, 4.885715, 4.88355, 4.883318, 4.884742, 4.887525, 4.891382, 
    4.89606, 4.901348, 4.907085, 4.913165, 4.919536, 4.926205, 4.93325, 
    4.940831, 4.945117, 4.948902, 4.955187, 4.960639, 4.96536, 4.969398, 
    4.97435, 4.977834, 4.980072, 4.981319, 4.981205, 4.979434, 4.975549, 
    4.969117, 4.959093, 4.944644, 4.928452, 4.909022, 4.887101, 4.86384, 
    4.840705, 4.81933, 4.801309, 4.787976, 4.780247, 4.778527, 4.782729, 
    4.792338, 4.806513, 4.824186, 4.844155, 4.865149, 4.885897, 4.905189, 
    4.921952,
  // totalHeight(18,14, 0-49)
    4.886841, 4.883399, 4.882051, 4.882535, 4.884551, 4.887797, 4.891985, 
    4.896872, 4.902257, 4.907996, 4.914003, 4.920245, 4.926744, 4.933584, 
    4.940909, 4.94667, 4.949551, 4.95581, 4.961526, 4.966652, 4.971175, 
    4.976239, 4.979972, 4.982547, 4.984378, 4.98511, 4.984487, 4.982019, 
    4.977257, 4.968933, 4.956161, 4.94096, 4.922206, 4.900504, 4.876897, 
    4.852814, 4.829932, 4.809971, 4.794442, 4.784451, 4.780582, 4.782882, 
    4.790926, 4.803923, 4.820827, 4.840441, 4.861489, 4.882676, 4.90276, 
    4.920603,
  // totalHeight(18,15, 0-49)
    4.883207, 4.880651, 4.880136, 4.881371, 4.884029, 4.887794, 4.892372, 
    4.897519, 4.903045, 4.908817, 4.914763, 4.920861, 4.927134, 4.93365, 
    4.940502, 4.948238, 4.950455, 4.956568, 4.962499, 4.96802, 4.973034, 
    4.978105, 4.982003, 4.984821, 4.987122, 4.988574, 4.988962, 4.987782, 
    4.984583, 4.977922, 4.966918, 4.952744, 4.934793, 4.913519, 4.889838, 
    4.865107, 4.84101, 4.819353, 4.801796, 4.789631, 4.783615, 4.783937, 
    4.790273, 4.801894, 4.817789, 4.836773, 4.857575, 4.878895, 4.899468, 
    4.918118,
  // totalHeight(18,16, 0-49)
    4.879242, 4.87754, 4.87785, 4.879844, 4.883172, 4.887492, 4.892501, 
    4.897952, 4.903658, 4.909498, 4.915406, 4.921362, 4.92738, 4.933488, 
    4.939705, 4.949776, 4.951613, 4.95754, 4.963687, 4.969635, 4.975175, 
    4.98018, 4.984186, 4.987179, 4.989842, 4.991875, 4.993103, 4.993021, 
    4.991203, 4.986084, 4.976843, 4.963641, 4.946527, 4.925811, 4.902266, 
    4.877148, 4.852115, 4.829021, 4.809649, 4.795449, 4.787349, 4.785682, 
    4.790234, 4.800347, 4.815056, 4.8332, 4.853517, 4.874714, 4.895517, 
    4.914725,
  // totalHeight(18,17, 0-49)
    4.875041, 4.874127, 4.875218, 4.87795, 4.881939, 4.886819, 4.892274, 
    4.898053, 4.903974, 4.909922, 4.915837, 4.921696, 4.927484, 4.933181, 
    4.938707, 4.951196, 4.952917, 4.958723, 4.965165, 4.971624, 4.977774, 
    4.982686, 4.986784, 4.989913, 4.992849, 4.995311, 4.997171, 4.997947, 
    4.997252, 4.993465, 4.9859, 4.973534, 4.95721, 4.937099, 4.913828, 
    4.888538, 4.862826, 4.838557, 4.817604, 4.801552, 4.791484, 4.787878, 
    4.790633, 4.799174, 4.812584, 4.829738, 4.849395, 4.870271, 4.891096, 
    4.910655,
  // totalHeight(18,18, 0-49)
    4.870688, 4.87046, 4.872247, 4.875643, 4.880235, 4.885635, 4.891515, 
    4.897624, 4.90379, 4.909906, 4.91592, 4.921796, 4.927487, 4.932893, 
    4.937829, 4.952391, 4.954152, 4.960028, 4.966936, 4.974069, 4.980973, 
    4.985815, 4.99005, 4.993322, 4.99646, 4.999198, 5.001451, 5.002779, 
    5.002877, 5.000129, 4.994055, 4.982319, 4.966665, 4.947137, 4.924218, 
    4.898921, 4.872756, 4.847573, 4.825289, 4.807601, 4.795727, 4.790283, 
    4.791286, 4.798248, 4.810311, 4.826389, 4.84527, 4.865687, 4.886379, 
    4.906126,
  // totalHeight(18,19, 0-49)
    4.86625, 4.86655, 4.868883, 4.872808, 4.877879, 4.883698, 4.889936, 
    4.896357, 4.902807, 4.909202, 4.915492, 4.921624, 4.927492, 4.932897, 
    4.937518, 4.953274, 4.955041, 4.961284, 4.968928, 4.976991, 4.984876, 
    4.989754, 4.994244, 4.997727, 5.001033, 5.003887, 5.006248, 5.007756, 
    5.008227, 5.006122, 5.001248, 4.98988, 4.974717, 4.955695, 4.933158, 
    4.907983, 4.881572, 4.855722, 4.832371, 4.813286, 4.799805, 4.792671, 
    4.792016, 4.797443, 4.808165, 4.823141, 4.841189, 4.861065, 4.881521, 
    4.901341,
  // totalHeight(18,20, 0-49)
    4.862615, 4.864183, 4.867981, 4.873559, 4.880429, 4.888097, 4.896105, 
    4.904039, 4.91155, 4.918352, 4.924236, 4.929071, 4.932817, 4.935514, 
    4.937287, 30, 4.967083, 4.970193, 4.974487, 4.979447, 4.9848, 4.986744, 
    4.989418, 4.992031, 4.995424, 4.999174, 5.003032, 5.006403, 5.008925, 
    5.008933, 5.006418, 4.996209, 4.982046, 4.963815, 4.941799, 4.916811, 
    4.8902, 4.86374, 4.83939, 4.818989, 4.803974, 4.79521, 4.792936, 
    4.796848, 4.806228, 4.820079, 4.837255, 4.856534, 4.87668, 4.896485,
  // totalHeight(18,21, 0-49)
    4.858526, 4.860593, 4.864909, 4.870983, 4.878288, 4.886311, 4.89458, 
    4.902694, 4.910328, 4.917231, 4.923228, 4.928211, 4.932137, 4.935033, 
    4.936998, 30, 4.96749, 4.971151, 4.976059, 4.981626, 4.987492, 4.988534, 
    4.990527, 4.992525, 4.995533, 4.999171, 5.003212, 5.007048, 5.010316, 
    5.011328, 5.010325, 5.000771, 4.987464, 4.970185, 4.949078, 4.924807, 
    4.898589, 4.872103, 4.847268, 4.82596, 4.809701, 4.799472, 4.795639, 
    4.798006, 4.805933, 4.818489, 4.834568, 4.852976, 4.872499, 4.891943,
  // totalHeight(18,22, 0-49)
    4.854605, 4.857058, 4.861805, 4.868328, 4.876069, 4.884493, 4.893115, 
    4.901526, 4.909408, 4.916522, 4.922707, 4.927864, 4.931949, 4.93498, 
    4.937038, 30, 4.968196, 4.972306, 4.977769, 4.98394, 4.990365, 4.990649, 
    4.992125, 4.993677, 4.996429, 5.000011, 5.004191, 5.008338, 5.01208, 
    5.013722, 5.013745, 5.004387, 4.991473, 4.974729, 4.954206, 4.930459, 
    4.904589, 4.878174, 4.853073, 4.831153, 4.813982, 4.802622, 4.797538, 
    4.798625, 4.805327, 4.816769, 4.831888, 4.849522, 4.86848, 4.887581,
  // totalHeight(18,23, 0-49)
    4.850917, 4.853661, 4.858761, 4.865675, 4.873829, 4.882668, 4.891686, 
    4.900468, 4.908682, 4.916094, 4.922538, 4.927917, 4.932185, 4.935344, 
    4.93747, 30, 4.969583, 4.973991, 4.979832, 4.98642, 4.993236, 4.992826, 
    4.993824, 4.99496, 4.99745, 5.000928, 5.005152, 5.009469, 5.013495, 
    5.015525, 5.016229, 5.006853, 4.994095, 4.977653, 4.95752, 4.934175, 
    4.908624, 4.882356, 4.857164, 4.834885, 4.817104, 4.804931, 4.798903, 
    4.798989, 4.804698, 4.81521, 4.8295, 4.846437, 4.864852, 4.883585,
  // totalHeight(18,24, 0-49)
    4.847519, 4.850479, 4.85586, 4.863112, 4.871647, 4.880895, 4.890332, 
    4.899526, 4.908134, 4.915905, 4.92267, 4.928324, 4.932813, 4.936135, 
    4.938357, 30, 4.971826, 4.976392, 4.982431, 4.989242, 4.996271, 4.995375, 
    4.996037, 4.996878, 4.999168, 5.002536, 5.006739, 5.011106, 5.015255, 
    5.017463, 5.018531, 5.009044, 4.996279, 4.979924, 4.959941, 4.936765, 
    4.911347, 4.885115, 4.859817, 4.837259, 4.819028, 4.806264, 4.799543, 
    4.798884, 4.803843, 4.813639, 4.827281, 4.843661, 4.86163, 4.880041,
  // totalHeight(18,25, 0-49)
    4.84447, 4.847589, 4.853196, 4.860741, 4.869628, 4.879272, 4.889136, 
    4.898769, 4.907809, 4.915988, 4.923122, 4.929097, 4.933853, 4.937385, 
    4.939763, 30, 4.974479, 4.979081, 4.985147, 4.991983, 4.999034, 4.997939, 
    4.99846, 4.999179, 5.001375, 5.00467, 5.008821, 5.013151, 5.017279, 
    5.019472, 5.020578, 5.010951, 4.998077, 4.981641, 4.961603, 4.938382, 
    4.91291, 4.88659, 4.861147, 4.838369, 4.819839, 4.806698, 4.799538, 
    4.7984, 4.802862, 4.81217, 4.825348, 4.841312, 4.858924, 4.877048,
  // totalHeight(18,26, 0-49)
    4.841846, 4.845082, 4.850876, 4.858679, 4.867893, 4.877924, 4.888223, 
    4.898314, 4.907815, 4.916437, 4.923976, 4.930305, 4.935359, 4.939139, 
    4.941726, 30, 4.977385, 4.981901, 4.98783, 4.994493, 5.001371, 5.000391, 
    5.000994, 5.001788, 5.004019, 5.007303, 5.01139, 5.015614, 5.019589, 
    5.021584, 5.022406, 5.012643, 4.999584, 4.982924, 4.962636, 4.939158, 
    4.913439, 4.886895, 4.861254, 4.838302, 4.819606, 4.806296, 4.798949, 
    4.797599, 4.801824, 4.810872, 4.823782, 4.839473, 4.856821, 4.874699,
  // totalHeight(18,27, 0-49)
    4.839744, 4.843068, 4.84902, 4.857059, 4.866587, 4.877005, 4.887747, 
    4.898317, 4.908307, 4.917399, 4.925366, 4.932062, 4.937419, 4.941448, 
    4.944248, 30, 4.980576, 4.984866, 4.990472, 4.996755, 5.003257, 5.002659, 
    5.003529, 5.004568, 5.006943, 5.01026, 5.014267, 5.018305, 5.021995, 
    5.023608, 5.023826, 5.013915, 5.000586, 4.983556, 4.962839, 4.938921, 
    4.912803, 4.885948, 4.860112, 4.837081, 4.818402, 4.805168, 4.797915, 
    4.796639, 4.800896, 4.809918, 4.822744, 4.838297, 4.855458, 4.873108,
  // totalHeight(18,28, 0-49)
    4.838279, 4.841671, 4.847761, 4.856022, 4.86586, 4.876674, 4.887884, 
    4.898968, 4.909482, 4.919071, 4.927473, 4.934519, 4.940135, 4.94435, 
    4.94729, 30, 4.984393, 4.988278, 4.993347, 4.999027, 5.004954, 5.004905, 
    5.006158, 5.007552, 5.010141, 5.013506, 5.017393, 5.021155, 5.024417, 
    5.025462, 5.024777, 5.014656, 5.000932, 4.983361, 4.962024, 4.937493, 
    4.910855, 4.883649, 4.857671, 4.834711, 4.816276, 4.803395, 4.796536, 
    4.795633, 4.800196, 4.80943, 4.82236, 4.837905, 4.854949, 4.872379,
  // totalHeight(18,29, 0-49)
    4.837578, 4.841016, 4.847223, 4.855696, 4.865859, 4.8771, 4.888828, 
    4.900484, 4.911574, 4.921689, 4.930514, 4.937848, 4.943614, 4.94786, 
    4.950751, 30, 4.988549, 4.991818, 4.996123, 5.000973, 5.006124, 5.006631, 
    5.00827, 5.010037, 5.012847, 5.016247, 5.019962, 5.023355, 5.02604, 
    5.026312, 5.024417, 5.013925, 4.999619, 4.981328, 4.959243, 4.93405, 
    4.906947, 4.879553, 4.853701, 4.831154, 4.813352, 4.801226, 4.795144, 
    4.794957, 4.800112, 4.80978, 4.822963, 4.83858, 4.855508, 4.872646,
  // totalHeight(18,30, 0-49)
    4.837201, 4.839952, 4.84534, 4.852841, 4.861905, 4.872, 4.882656, 
    4.893489, 4.904216, 4.914642, 4.924639, 4.934104, 4.942914, 4.950874, 
    4.957664, 4.980512, 4.978384, 4.985451, 4.993881, 5.002621, 5.011064, 
    5.015289, 5.019503, 5.022801, 5.026014, 5.028763, 5.03095, 5.032186, 
    5.032328, 5.02988, 5.02498, 5.012665, 4.996644, 4.97683, 4.95351, 
    4.927465, 4.899968, 4.872666, 4.847361, 4.825732, 4.809091, 4.798231, 
    4.793395, 4.794331, 4.800419, 4.81079, 4.824425, 4.840233, 4.8571, 
    4.873925,
  // totalHeight(18,31, 0-49)
    4.838711, 4.841673, 4.847275, 4.855004, 4.864307, 4.874646, 4.885531, 
    4.896559, 4.907419, 4.917896, 4.927857, 4.937228, 4.945951, 4.953948, 
    4.961065, 4.980995, 4.980417, 4.987096, 4.994756, 5.002519, 5.00993, 
    5.014159, 5.018117, 5.021186, 5.024208, 5.026828, 5.028913, 5.029993, 
    5.029801, 5.02675, 5.020671, 5.008065, 4.991631, 4.971384, 4.94774, 
    4.9216, 4.89433, 4.86762, 4.843251, 4.822825, 4.807539, 4.798059, 
    4.794508, 4.796546, 4.803485, 4.814416, 4.828295, 4.844025, 4.860487, 
    4.876597,
  // totalHeight(18,32, 0-49)
    4.841342, 4.844412, 4.850084, 4.857855, 4.867183, 4.877531, 4.888418, 
    4.899436, 4.910273, 4.920713, 4.930632, 4.93998, 4.948754, 4.956964, 
    4.964594, 4.980965, 4.981505, 4.988069, 4.995195, 5.002202, 5.00878, 
    5.013144, 5.016983, 5.019907, 5.02272, 5.025066, 5.026776, 5.02734, 
    5.026409, 5.022374, 5.014822, 5.001704, 4.984722, 4.964009, 4.940114, 
    4.914057, 4.88728, 4.861488, 4.838411, 4.819547, 4.80595, 4.798151, 
    4.796151, 4.799515, 4.807491, 4.819123, 4.833344, 4.849035, 4.865076, 
    4.880392,
  // totalHeight(18,33, 0-49)
    4.845201, 4.848296, 4.853919, 4.861576, 4.870737, 4.880888, 4.891561, 
    4.902365, 4.912999, 4.923262, 4.933043, 4.942318, 4.951126, 4.959552, 
    4.967697, 4.980441, 4.981912, 4.988523, 4.995258, 5.001646, 5.007523, 
    5.012081, 5.015876, 5.018697, 5.021259, 5.023195, 5.024305, 5.02406, 
    5.022061, 5.016749, 5.007536, 4.993733, 4.976113, 4.954939, 4.930896, 
    4.905118, 4.879101, 4.85454, 4.833084, 4.816096, 4.804484, 4.798627, 
    4.798405, 4.803288, 4.812459, 4.824915, 4.839553, 4.855231, 4.870821, 
    4.885258,
  // totalHeight(18,34, 0-49)
    4.850313, 4.853356, 4.858818, 4.866215, 4.875041, 4.884804, 4.895066, 
    4.905462, 4.915716, 4.925641, 4.935148, 4.944232, 4.952967, 4.961494, 
    4.970001, 4.979457, 4.981847, 4.98854, 4.994935, 5.000776, 5.006025, 
    5.010772, 5.014541, 5.01726, 5.019513, 5.020917, 5.02124, 5.019953, 
    5.016633, 5.00984, 4.998881, 4.98429, 4.966008, 4.944437, 4.920403, 
    4.895131, 4.870153, 4.847122, 4.82758, 4.812739, 4.803346, 4.799632, 
    4.801355, 4.8079, 4.818378, 4.831736, 4.846831, 4.862496, 4.877587, 
    4.891049,
  // totalHeight(18,35, 0-49)
    4.85662, 4.859527, 4.864711, 4.871711, 4.880044, 4.889249, 4.898926, 
    4.908741, 4.918445, 4.927876, 4.936965, 4.94572, 4.954232, 4.962675, 
    4.971297, 4.978046, 4.981433, 4.988136, 4.99417, 4.999484, 5.004143, 
    5.009024, 5.012743, 5.015333, 5.017207, 5.017971, 5.017355, 5.014852, 
    5.01003, 5.001642, 4.988949, 4.973538, 4.954648, 4.932821, 4.909005, 
    4.884502, 4.860847, 4.839624, 4.822244, 4.809759, 4.80275, 4.801305, 
    4.805072, 4.813345, 4.825176, 4.839457, 4.855005, 4.870616, 4.885136, 
    4.89752,
  // totalHeight(18,36, 0-49)
    4.863973, 4.866647, 4.871443, 4.877914, 4.885613, 4.894113, 4.903052, 
    4.912133, 4.921141, 4.929941, 4.938475, 4.946762, 4.954895, 4.963057, 
    4.971507, 4.97621, 4.980695, 4.987263, 4.992869, 4.997642, 5.001723, 
    5.006649, 5.010259, 5.012672, 5.014094, 5.014126, 5.01246, 5.008624, 
    5.0022, 4.992191, 4.977875, 4.961699, 4.942339, 4.920467, 4.897135, 
    4.87369, 4.85164, 4.83247, 4.817447, 4.807454, 4.802914, 4.80378, 
    4.809597, 4.819584, 4.832732, 4.847884, 4.863813, 4.879286, 4.893135, 
    4.904335,
  // totalHeight(18,37, 0-49)
    4.872146, 4.874485, 4.878777, 4.884603, 4.891544, 4.899216, 4.907293, 
    4.91552, 4.923715, 4.931767, 4.939631, 4.947328, 4.954942, 4.962633, 
    4.970646, 4.973928, 4.979574, 4.985822, 4.990914, 4.995116, 4.99861, 
    5.003463, 5.006887, 5.00906, 5.009962, 5.009189, 5.006405, 5.001185, 
    4.993144, 4.981586, 4.965855, 4.949062, 4.929453, 4.907815, 4.885276, 
    4.863191, 4.843011, 4.8261, 4.813562, 4.806119, 4.804044, 4.807168, 
    4.814948, 4.826537, 4.840876, 4.856761, 4.872931, 4.888124, 4.901169, 
    4.911073,
  // totalHeight(18,38, 0-49)
    4.880842, 4.882741, 4.886423, 4.891498, 4.897586, 4.904336, 4.911465, 
    4.918751, 4.926048, 4.933264, 4.940367, 4.947376, 4.954354, 4.961426, 
    4.968778, 4.971156, 4.977955, 4.983696, 4.988179, 4.991767, 4.994656, 
    4.999306, 5.002451, 5.004314, 5.004631, 5.003013, 4.999096, 4.992517, 
    4.982934, 4.969998, 4.953146, 4.935975, 4.916419, 4.895351, 4.873941, 
    4.853517, 4.83544, 4.820933, 4.810941, 4.806021, 4.806313, 4.811546, 
    4.821102, 4.834083, 4.849388, 4.86578, 4.881971, 4.896688, 4.908768, 
    4.917272,
  // totalHeight(18,39, 0-49)
    4.889717, 4.891066, 4.894044, 4.898291, 4.903454, 4.909225, 4.915352, 
    4.921652, 4.927999, 4.934326, 4.940608, 4.946858, 4.953117, 4.959458, 
    4.965996, 4.96784, 4.975702, 4.980766, 4.984552, 4.987484, 4.989732, 
    4.99404, 4.996809, 4.998293, 4.997983, 4.995514, 4.990504, 4.982667, 
    4.971714, 4.957668, 4.940073, 4.922842, 4.903699, 4.883575, 4.863635, 
    4.84515, 4.829363, 4.817347, 4.809879, 4.807374, 4.809848, 4.816947, 
    4.827996, 4.842059, 4.858009, 4.874594, 4.890515, 4.904504, 4.915439, 
    4.922453,
  // totalHeight(18,40, 0-49)
    4.8984, 4.899097, 4.90129, 4.904646, 4.908849, 4.913617, 4.91873, 
    4.924032, 4.929419, 4.934838, 4.940274, 4.945725, 4.951211, 4.956755, 
    4.96239, 4.963936, 4.972683, 4.976931, 4.979949, 4.982178, 4.983747, 
    4.987577, 4.989875, 4.990921, 4.989964, 4.98668, 4.98068, 4.971765, 
    4.959704, 4.944898, 4.927004, 4.910091, 4.891764, 4.872965, 4.854824, 
    4.838517, 4.825151, 4.815638, 4.810602, 4.81032, 4.814709, 4.823346, 
    4.835516, 4.850266, 4.866456, 4.882841, 4.898137, 4.911113, 4.920713, 
    4.926178,
  // totalHeight(18,41, 0-49)
    4.906529, 4.906476, 4.907814, 4.910242, 4.91347, 4.917244, 4.921369, 
    4.925701, 4.930154, 4.934687, 4.939281, 4.94393, 4.948625, 4.953344, 
    4.958044, 4.959407, 4.968792, 4.97213, 4.974324, 4.975806, 4.976653, 
    4.979882, 4.981626, 4.98219, 4.980597, 4.976579, 4.969752, 4.960011, 
    4.947186, 4.932035, 4.914319, 4.898144, 4.881041, 4.863939, 4.847887, 
    4.833943, 4.823065, 4.816005, 4.813236, 4.814918, 4.820882, 4.830656, 
    4.843504, 4.858468, 4.874428, 4.890163, 4.904439, 4.916101, 4.924196, 
    4.928107,
  // totalHeight(18,42, 0-49)
    4.913782, 4.912883, 4.913308, 4.914782, 4.917043, 4.919858, 4.923043, 
    4.926467, 4.93005, 4.933751, 4.937549, 4.941423, 4.945343, 4.949245, 
    4.953024, 4.954234, 4.963964, 4.96634, 4.967675, 4.96837, 4.968452, 
    4.970979, 4.972106, 4.972164, 4.969982, 4.965353, 4.957918, 4.947659, 
    4.934467, 4.919428, 4.902383, 4.887368, 4.871888, 4.856811, 4.843086, 
    4.831631, 4.823244, 4.818518, 4.817794, 4.821123, 4.82827, 4.83873, 
    4.851759, 4.866421, 4.881636, 4.896245, 4.9091, 4.919161, 4.925624, 
    4.928048,
  // totalHeight(18,43, 0-49)
    4.919908, 4.918075, 4.917529, 4.918031, 4.919343, 4.921244, 4.923561, 
    4.926164, 4.928969, 4.931925, 4.934999, 4.938159, 4.941349, 4.944471, 
    4.947376, 4.948405, 4.958177, 4.959578, 4.960035, 4.959912, 4.959199, 
    4.960948, 4.961421, 4.960978, 4.958283, 4.953208, 4.945422, 4.934996, 
    4.921866, 4.907401, 4.8915, 4.878047, 4.864542, 4.851766, 4.840542, 
    4.831635, 4.82568, 4.823121, 4.824172, 4.828796, 4.8367, 4.847362, 
    4.860054, 4.873881, 4.887831, 4.900847, 4.911908, 4.920138, 4.924921, 
    4.926015,
  // totalHeight(18,44, 0-49)
    4.924776, 4.921913, 4.92034, 4.91985, 4.920226, 4.921264, 4.92279, 
    4.924667, 4.926798, 4.929115, 4.931567, 4.934095, 4.936621, 4.939024, 
    4.941122, 4.941914, 4.951438, 4.951888, 4.951467, 4.95051, 4.94899, 
    4.94992, 4.94973, 4.948813, 4.945714, 4.940386, 4.932531, 4.9223, 
    4.909667, 4.896218, 4.881884, 4.870344, 4.859107, 4.848838, 4.840219, 
    4.833856, 4.830224, 4.829626, 4.832157, 4.837701, 4.845929, 4.856311, 
    4.868156, 4.880635, 4.89284, 4.903851, 4.912822, 4.91908, 4.922236, 
    4.922259,
  // totalHeight(18,45, 0-49)
    4.928407, 4.924418, 4.921751, 4.920234, 4.919677, 4.919885, 4.920683, 
    4.921923, 4.923484, 4.925271, 4.927204, 4.929194, 4.931141, 4.932897, 
    4.934264, 4.934757, 4.943786, 4.943328, 4.942047, 4.94026, 4.937941, 
    4.93805, 4.937223, 4.935887, 4.932515, 4.927137, 4.9195, 4.909817, 
    4.898086, 4.886047, 4.873634, 4.864293, 4.855537, 4.847908, 4.841933, 
    4.838057, 4.836599, 4.837729, 4.841436, 4.847537, 4.855672, 4.865327, 
    4.875862, 4.886545, 4.896604, 4.9053, 4.912002, 4.916276, 4.917975, 
    4.917284,
  // totalHeight(18,46, 0-49)
    4.931002, 4.925789, 4.921949, 4.919353, 4.917837, 4.917222, 4.917328, 
    4.917989, 4.919061, 4.920411, 4.921917, 4.92346, 4.924904, 4.926087, 
    4.926797, 4.926932, 4.935273, 4.933967, 4.931861, 4.929269, 4.926188, 
    4.925509, 4.924102, 4.922422, 4.918921, 4.9137, 4.906552, 4.897737, 
    4.887263, 4.876956, 4.866735, 4.859797, 4.853657, 4.848723, 4.845367, 
    4.843875, 4.844419, 4.84704, 4.851633, 4.857956, 4.865634, 4.87418, 
    4.883031, 4.891579, 4.899223, 4.905437, 4.90984, 4.912262, 4.912797, 
    4.911825,
  // totalHeight(18,47, 0-49)
    4.932955, 4.926421, 4.921322, 4.91757, 4.91504, 4.913567, 4.912973, 
    4.913074, 4.91369, 4.914652, 4.915792, 4.916949, 4.917954, 4.91862, 
    4.918736, 4.91845, 4.925973, 4.923887, 4.921003, 4.917657, 4.913873, 
    4.912481, 4.910572, 4.908642, 4.905159, 4.900286, 4.893863, 4.88618, 
    4.877249, 4.868914, 4.861065, 4.856644, 4.853178, 4.850926, 4.850114, 
    4.850874, 4.853234, 4.85712, 4.862342, 4.86861, 4.875546, 4.88271, 
    4.88963, 4.895852, 4.900975, 4.904717, 4.906961, 4.907805, 4.907571, 
    4.906791,
  // totalHeight(18,48, 0-49)
    4.934845, 4.9269, 4.920446, 4.915445, 4.911812, 4.909406, 4.908049, 
    4.907547, 4.907685, 4.908252, 4.909031, 4.909818, 4.910404, 4.910583, 
    4.91014, 4.909373, 4.916004, 4.9132, 4.909599, 4.905562, 4.90116, 
    4.899149, 4.896842, 4.894763, 4.891435, 4.887076, 4.881566, 4.875215, 
    4.868028, 4.861816, 4.856431, 4.854557, 4.85374, 4.854105, 4.855721, 
    4.858578, 4.862577, 4.867533, 4.873183, 4.879201, 4.885219, 4.890858, 
    4.895762, 4.899647, 4.902333, 4.903794, 4.904185, 4.903849, 4.903304, 
    4.90318,
  // totalHeight(18,49, 0-49)
    4.943079, 4.933022, 4.92444, 4.917368, 4.911783, 4.907586, 4.904629, 
    4.902708, 4.901586, 4.901, 4.900681, 4.900353, 4.899747, 4.898587, 
    4.896599, 4.894702, 4.907625, 4.902482, 4.896469, 4.890329, 4.884231, 
    4.883526, 4.882961, 4.883486, 4.882074, 4.87913, 4.874318, 4.868094, 
    4.860242, 4.854196, 4.849467, 4.851037, 4.85378, 4.857646, 4.86253, 
    4.868235, 4.874485, 4.880953, 4.887276, 4.893087, 4.898046, 4.901875, 
    4.904406, 4.905601, 4.905601, 4.904716, 4.90344, 4.902396, 4.902278, 
    4.903772,
  // totalHeight(19,0, 0-49)
    4.863467, 4.857262, 4.854007, 4.853439, 4.855211, 4.858918, 4.86413, 
    4.870421, 4.877393, 4.884692, 4.892019, 4.899126, 4.905809, 4.911901, 
    4.917256, 4.921696, 4.926414, 4.929109, 4.930936, 4.931877, 4.931879, 
    4.93122, 4.92947, 4.92665, 4.922586, 4.917221, 4.910484, 4.902398, 
    4.893026, 4.882643, 4.871445, 4.860118, 4.848811, 4.838039, 4.828342, 
    4.820229, 4.814119, 4.8103, 4.808887, 4.80981, 4.812818, 4.817494, 
    4.823306, 4.829645, 4.835906, 4.841548, 4.846171, 4.849586, 4.85186, 
    4.853332,
  // totalHeight(19,1, 0-49)
    4.865608, 4.859947, 4.857208, 4.857111, 4.8593, 4.863361, 4.868865, 
    4.875392, 4.882556, 4.890017, 4.897492, 4.904748, 4.911586, 4.917842, 
    4.923354, 4.927824, 4.933651, 4.936447, 4.938407, 4.939521, 4.939701, 
    4.939492, 4.938069, 4.935489, 4.931462, 4.925898, 4.918675, 4.909807, 
    4.899339, 4.887649, 4.874897, 4.862156, 4.849326, 4.837008, 4.825834, 
    4.816401, 4.809213, 4.804626, 4.802801, 4.803697, 4.807059, 4.812455, 
    4.8193, 4.826921, 4.834619, 4.841738, 4.847753, 4.85234, 4.855436, 
    4.857277,
  // totalHeight(19,2, 0-49)
    4.868079, 4.86294, 4.86067, 4.86098, 4.863502, 4.867823, 4.873523, 
    4.880189, 4.887453, 4.894991, 4.90254, 4.909874, 4.91681, 4.923179, 
    4.928813, 4.933246, 4.940066, 4.942986, 4.945104, 4.946426, 4.946843, 
    4.947165, 4.946175, 4.943969, 4.940157, 4.934615, 4.927167, 4.917808, 
    4.90655, 4.893838, 4.879786, 4.865834, 4.851622, 4.837819, 4.825143, 
    4.814283, 4.805833, 4.800229, 4.7977, 4.798252, 4.801656, 4.807476, 
    4.815114, 4.823852, 4.832918, 4.841565, 4.849153, 4.855217, 4.859553, 
    4.862253,
  // totalHeight(19,3, 0-49)
    4.870552, 4.86591, 4.864064, 4.864718, 4.867503, 4.872014, 4.877833, 
    4.884569, 4.891868, 4.899426, 4.906993, 4.914361, 4.921353, 4.927806, 
    4.93355, 4.937875, 4.945512, 4.948591, 4.950888, 4.952444, 4.953139, 
    4.954044, 4.953572, 4.95185, 4.948418, 4.943113, 4.935712, 4.926178, 
    4.914483, 4.901093, 4.886057, 4.871165, 4.855776, 4.840611, 4.826462, 
    4.814105, 4.804229, 4.797366, 4.793829, 4.793693, 4.796775, 4.802673, 
    4.810785, 4.820376, 4.830633, 4.840738, 4.84995, 4.857678, 4.863564, 
    4.867543,
  // totalHeight(19,4, 0-49)
    4.872817, 4.868643, 4.867184, 4.868135, 4.871129, 4.875768, 4.881651, 
    4.888405, 4.895691, 4.903227, 4.910775, 4.918141, 4.92516, 4.931677, 
    4.937528, 4.941673, 4.949905, 4.953179, 4.955673, 4.957477, 4.958472, 
    4.959987, 4.960082, 4.958926, 4.956011, 4.951143, 4.944056, 4.934675, 
    4.922916, 4.909231, 4.893579, 4.878071, 4.861773, 4.845433, 4.829899, 
    4.816028, 4.804605, 4.796266, 4.79143, 4.790257, 4.792642, 4.798227, 
    4.806442, 4.816557, 4.827739, 4.839124, 4.849892, 4.859341, 4.866971, 
    4.872547,
  // totalHeight(19,5, 0-49)
    4.874774, 4.871048, 4.869942, 4.871148, 4.874307, 4.879029, 4.884934, 
    4.891664, 4.898901, 4.906378, 4.913873, 4.921207, 4.928225, 4.93479, 
    4.940752, 4.944649, 4.953211, 4.956712, 4.959419, 4.961472, 4.962777, 
    4.964893, 4.965576, 4.96503, 4.962738, 4.958478, 4.951951, 4.943034, 
    4.931594, 4.918012, 4.902144, 4.886379, 4.869491, 4.852226, 4.835463, 
    4.820125, 4.807089, 4.797104, 4.790708, 4.788169, 4.789482, 4.79436, 
    4.802285, 4.812552, 4.824332, 4.836738, 4.848891, 4.860003, 4.869445, 
    4.876825,
  // totalHeight(19,6, 0-49)
    4.876401, 4.873109, 4.872334, 4.873767, 4.877055, 4.881827, 4.887718, 
    4.894387, 4.901539, 4.90892, 4.916327, 4.923593, 4.930583, 4.937176, 
    4.943255, 4.946844, 4.955447, 4.959205, 4.962132, 4.964428, 4.966038, 
    4.968722, 4.969982, 4.970057, 4.968456, 4.964935, 4.959171, 4.951004, 
    4.94024, 4.92715, 4.911473, 4.895832, 4.878706, 4.860817, 4.843043, 
    4.826352, 4.811706, 4.799966, 4.7918, 4.78761, 4.787505, 4.791297, 
    4.798542, 4.808578, 4.820599, 4.833713, 4.847009, 4.85963, 4.870845, 
    4.880115,
  // totalHeight(19,7, 0-49)
    4.877742, 4.87488, 4.87442, 4.876059, 4.879453, 4.884243, 4.890086, 
    4.896661, 4.903688, 4.910936, 4.918213, 4.925372, 4.932297, 4.938896, 
    4.945095, 4.948344, 4.956688, 4.960714, 4.963864, 4.966398, 4.968299, 
    4.971492, 4.973291, 4.973963, 4.973082, 4.970386, 4.965547, 4.958364, 
    4.94859, 4.936349, 4.921254, 4.906102, 4.889108, 4.870925, 4.852411, 
    4.83455, 4.818367, 4.804838, 4.79476, 4.78869, 4.78687, 4.789238, 
    4.795435, 4.80487, 4.816771, 4.830261, 4.844414, 4.858326, 4.871181, 
    4.882321,
  // totalHeight(19,8, 0-49)
    4.878867, 4.876438, 4.876289, 4.878121, 4.881602, 4.886387, 4.892151, 
    4.898596, 4.90546, 4.912529, 4.919632, 4.926641, 4.93346, 4.940037, 
    4.946343, 4.94926, 4.957064, 4.961346, 4.964719, 4.967476, 4.969651, 
    4.973279, 4.975556, 4.976775, 4.976603, 4.974774, 4.970967, 4.964946, 
    4.956418, 4.94533, 4.931167, 4.916834, 4.900319, 4.88219, 4.863243, 
    4.844447, 4.826875, 4.811594, 4.799544, 4.791435, 4.787673, 4.788329, 
    4.793161, 4.801657, 4.813101, 4.826638, 4.841345, 4.856289, 4.87059, 
    4.883487,
  // totalHeight(19,9, 0-49)
    4.879853, 4.877869, 4.878036, 4.880059, 4.883614, 4.888375, 4.894034, 
    4.900314, 4.906975, 4.913821, 4.920701, 4.927508, 4.934181, 4.940696, 
    4.94708, 4.94973, 4.956745, 4.961252, 4.964836, 4.967809, 4.970237, 
    4.974212, 4.976891, 4.978584, 4.979081, 4.978118, 4.975397, 4.970651, 
    4.963554, 4.953855, 4.940918, 4.927673, 4.911951, 4.894206, 4.875144, 
    4.855691, 4.836935, 4.820017, 4.80601, 4.795788, 4.789926, 4.788655, 
    4.791863, 4.799135, 4.809819, 4.823099, 4.838062, 4.853761, 4.86927, 
    4.883741,
  // totalHeight(19,10, 0-49)
    4.880766, 4.879248, 4.879743, 4.881961, 4.885587, 4.890312, 4.895844, 
    4.901929, 4.90835, 4.91493, 4.921543, 4.928103, 4.934577, 4.940979, 
    4.947385, 4.949909, 4.955944, 4.960614, 4.964392, 4.967567, 4.970238, 
    4.974462, 4.977457, 4.979537, 4.980639, 4.980505, 4.978874, 4.975456, 
    4.969903, 4.961752, 4.950266, 4.938305, 4.923625, 4.906556, 4.887687, 
    4.867873, 4.848182, 4.829807, 4.813938, 4.801608, 4.79357, 4.79023, 
    4.79162, 4.797441, 4.807114, 4.819869, 4.834813, 4.850992, 4.867447, 
    4.883266,
  // totalHeight(19,11, 0-49)
    4.881644, 4.880621, 4.881466, 4.883892, 4.887596, 4.892278, 4.897672, 
    4.903541, 4.909692, 4.91597, 4.922273, 4.92854, 4.934764, 4.94099, 
    4.94733, 4.949949, 4.954883, 4.959633, 4.963575, 4.966947, 4.969853, 
    4.974226, 4.977445, 4.979825, 4.981448, 4.982079, 4.9815, 4.979406, 
    4.975439, 4.968922, 4.95904, 4.948476, 4.935015, 4.918853, 4.900454, 
    4.880566, 4.860214, 4.840611, 4.823038, 4.80868, 4.798471, 4.792996, 
    4.792449, 4.796651, 4.805115, 4.817122, 4.8318, 4.8482, 4.865337, 4.882246,
  // totalHeight(19,12, 0-49)
    4.882496, 4.881999, 4.883224, 4.885882, 4.889676, 4.894325, 4.899577, 
    4.90522, 4.911082, 4.917034, 4.922996, 4.928931, 4.934853, 4.940827, 
    4.946981, 4.949989, 4.95378, 4.958515, 4.962585, 4.966149, 4.969291, 
    4.973717, 4.977075, 4.979658, 4.981715, 4.983027, 4.983429, 4.982606, 
    4.9802, 4.975337, 4.967144, 4.958006, 4.945863, 4.930773, 4.913065, 
    4.893366, 4.872625, 4.852049, 4.832983, 4.816743, 4.804437, 4.796834, 
    4.794295, 4.796777, 4.803885, 4.814964, 4.829169, 4.845552, 4.863111, 
    4.880845,
  // totalHeight(19,13, 0-49)
    4.883292, 4.883357, 4.884997, 4.887918, 4.891829, 4.896464, 4.901587, 
    4.907006, 4.912575, 4.918189, 4.923789, 4.929358, 4.934927, 4.940565, 
    4.94639, 4.950139, 4.952823, 4.957446, 4.961614, 4.96537, 4.968758, 
    4.973145, 4.976562, 4.979265, 4.981663, 4.983564, 4.98485, 4.985204, 
    4.984283, 4.981029, 4.974552, 4.966794, 4.955986, 4.942058, 4.9252, 
    4.905908, 4.885034, 4.863748, 4.84343, 4.825501, 4.811233, 4.801569, 
    4.797047, 4.797762, 4.803423, 4.813437, 4.826993, 4.84315, 4.86089, 
    4.879182,
  // totalHeight(19,14, 0-49)
    4.883975, 4.884635, 4.886726, 4.889947, 4.894012, 4.898662, 4.903681, 
    4.908897, 4.914186, 4.919464, 4.924696, 4.929881, 4.935049, 4.940267, 
    4.945613, 4.950459, 4.952142, 4.956577, 4.960824, 4.964785, 4.968439, 
    4.972709, 4.976121, 4.978877, 4.981533, 4.983922, 4.985978, 4.987384, 
    4.98782, 4.986081, 4.981294, 4.974806, 4.965281, 4.952532, 4.936615, 
    4.917893, 4.897106, 4.875359, 4.85404, 4.83465, 4.818594, 4.806993, 
    4.800546, 4.799497, 4.803661, 4.812512, 4.825278, 4.841026, 4.858731, 
    4.877334,
  // totalHeight(19,15, 0-49)
    4.884464, 4.885746, 4.888322, 4.891884, 4.896142, 4.900849, 4.905801, 
    4.910846, 4.915881, 4.920848, 4.925724, 4.930517, 4.93526, 4.939989, 
    4.94473, 4.95096, 4.951797, 4.956015, 4.960347, 4.964542, 4.968503, 
    4.972597, 4.97596, 4.978716, 4.981555, 4.984333, 4.987031, 4.989339, 
    4.990971, 4.990606, 4.987436, 4.98206, 4.973706, 4.962089, 4.94714, 
    4.929091, 4.908561, 4.886575, 4.864501, 4.843886, 4.82625, 4.812865, 
    4.804594, 4.801823, 4.804478, 4.812106, 4.823973, 4.83916, 4.856639, 
    4.875334,
  // totalHeight(19,16, 0-49)
    4.884663, 4.88658, 4.889668, 4.893605, 4.898099, 4.902907, 4.907837, 
    4.912756, 4.917584, 4.922279, 4.926834, 4.931263, 4.935582, 4.939795, 
    4.943863, 4.951606, 4.951766, 4.955799, 4.960267, 4.964756, 4.969089, 
    4.972967, 4.976264, 4.978997, 4.981962, 4.985034, 4.988237, 4.991272, 
    4.993902, 4.994734, 4.993072, 4.988607, 4.981264, 4.970675, 4.956662, 
    4.93933, 4.919178, 4.897139, 4.874533, 4.85293, 4.833932, 4.818943, 
    4.808976, 4.804556, 4.805722, 4.812094, 4.822984, 4.837489, 4.854583, 
    4.873177,
  // totalHeight(19,17, 0-49)
    4.884471, 4.887014, 4.890623, 4.894957, 4.899719, 4.904669, 4.909626, 
    4.914478, 4.919161, 4.923654, 4.92796, 4.932091, 4.936043, 4.939777, 
    4.943196, 4.952326, 4.951941, 4.9559, 4.960605, 4.965496, 4.970294, 
    4.973958, 4.977208, 4.979924, 4.982979, 4.986258, 4.989816, 4.993383, 
    4.996779, 4.998592, 4.998283, 4.994504, 4.987976, 4.978271, 4.96511, 
    4.948489, 4.928789, 4.90684, 4.883897, 4.861527, 4.841388, 4.824988, 
    4.813472, 4.8075, 4.807219, 4.81233, 4.822189, 4.835921, 4.852504, 
    4.870842,
  // totalHeight(19,18, 0-49)
    4.883793, 4.886919, 4.891025, 4.895751, 4.900793, 4.905913, 4.910947, 
    4.915798, 4.920425, 4.924825, 4.929009, 4.932978, 4.936702, 4.940094, 
    4.94299, 4.953041, 4.952164, 4.956231, 4.961337, 4.966779, 4.972184, 
    4.975669, 4.978938, 4.981686, 4.984823, 4.988232, 4.991991, 4.995869, 
    4.999767, 5.002297, 5.003136, 4.999793, 4.993859, 4.984858, 4.972429, 
    4.956472, 4.937254, 4.915499, 4.892387, 4.869453, 4.848384, 4.830771, 
    4.817868, 4.810457, 4.808792, 4.812659, 4.821465, 4.834362, 4.850341, 
    4.868311,
  // totalHeight(19,19, 0-49)
    4.882538, 4.886151, 4.890681, 4.895749, 4.901048, 4.906345, 4.911496, 
    4.916429, 4.921131, 4.92561, 4.929882, 4.933926, 4.937669, 4.94096, 
    4.943571, 4.95371, 4.952253, 4.956655, 4.962374, 4.968572, 4.974777, 
    4.978183, 4.981593, 4.984472, 4.987724, 4.991202, 4.994999, 4.998935, 
    5.003021, 5.00595, 5.007671, 5.004481, 4.998894, 4.990393, 4.978553, 
    4.963183, 4.944447, 4.922963, 4.899824, 4.876513, 4.854719, 4.836087, 
    4.821965, 4.813243, 4.810278, 4.812939, 4.820692, 4.832723, 4.848042, 
    4.865566,
  // totalHeight(19,20, 0-49)
    4.881588, 4.886601, 4.892593, 4.899169, 4.905969, 4.912692, 4.919097, 
    4.924998, 4.930258, 4.934787, 4.938541, 4.941516, 4.943758, 4.94535, 
    4.946416, 30, 4.960864, 4.963375, 4.966852, 4.970822, 4.975077, 4.975944, 
    4.977604, 4.979422, 4.982367, 4.986216, 4.99093, 4.996161, 5.00179, 
    5.006393, 5.010077, 5.007852, 5.003162, 4.995485, 4.98438, 4.969624, 
    4.951338, 4.930086, 4.906902, 4.883231, 4.860764, 4.841182, 4.825912, 
    4.815937, 4.811708, 4.813176, 4.819865, 4.831002, 4.845614, 4.862631,
  // totalHeight(19,21, 0-49)
    4.87942, 4.884988, 4.891505, 4.898539, 4.905715, 4.912723, 4.919326, 
    4.92536, 4.930717, 4.935334, 4.939191, 4.942301, 4.944708, 4.946493, 
    4.947779, 30, 4.960035, 4.963074, 4.967126, 4.971672, 4.976431, 4.976584, 
    4.977723, 4.979072, 4.98174, 4.985524, 4.990396, 4.995993, 5.002195, 
    5.007564, 5.012428, 5.010612, 5.006535, 4.999634, 4.989399, 4.975526, 
    4.958041, 4.937399, 4.914538, 4.890834, 4.867946, 4.84758, 4.831234, 
    4.819987, 4.814397, 4.814506, 4.819916, 4.829904, 4.843533, 4.859751,
  // totalHeight(19,22, 0-49)
    4.876799, 4.882879, 4.889917, 4.897455, 4.905089, 4.912499, 4.919439, 
    4.925747, 4.931327, 4.936132, 4.940154, 4.943415, 4.945968, 4.947898, 
    4.949335, 30, 4.959913, 4.963387, 4.967949, 4.973043, 4.978314, 4.977839, 
    4.978555, 4.979537, 4.982003, 4.985746, 4.990732, 4.996574, 5.003149, 
    5.009007, 5.014683, 5.012933, 5.009101, 5.002608, 4.992905, 4.97964, 
    4.962763, 4.942643, 4.920128, 4.896511, 4.873403, 4.852501, 4.835343, 
    4.823078, 4.816355, 4.815298, 4.819583, 4.828539, 4.841269, 4.856745,
  // totalHeight(19,23, 0-49)
    4.873835, 4.880381, 4.887924, 4.895979, 4.904121, 4.912008, 4.91938, 
    4.926068, 4.931972, 4.937049, 4.941298, 4.944747, 4.947457, 4.949518, 
    4.951072, 30, 4.960715, 4.964478, 4.969381, 4.974841, 4.980453, 4.979389, 
    4.979692, 4.980315, 4.982558, 4.986212, 4.991232, 4.997212, 5.004019, 
    5.010185, 5.016409, 5.014583, 5.010819, 5.004539, 4.995176, 4.982343, 
    4.96594, 4.946269, 4.924097, 4.900642, 4.877457, 4.856218, 4.838474, 
    4.825424, 4.817783, 4.815747, 4.819055, 4.827091, 4.838994, 4.853765,
  // totalHeight(19,24, 0-49)
    4.870672, 4.877634, 4.885653, 4.894224, 4.902894, 4.911297, 4.91916, 
    4.926295, 4.932595, 4.93801, 4.94254, 4.946218, 4.949106, 4.951304, 
    4.952971, 30, 4.962595, 4.966502, 4.971569, 4.977206, 4.982986, 4.981498, 
    4.981503, 4.981868, 4.98394, 4.987504, 4.992511, 4.998539, 5.005456, 
    5.011777, 5.018311, 5.016373, 5.012581, 5.006359, 4.997128, 4.984486, 
    4.968306, 4.948847, 4.926829, 4.903417, 4.880123, 4.858602, 4.840403, 
    4.826757, 4.818415, 4.815626, 4.818173, 4.82548, 4.836718, 4.850913,
  // totalHeight(19,25, 0-49)
    4.867481, 4.874813, 4.883271, 4.892335, 4.901527, 4.91046, 4.918839, 
    4.926459, 4.933195, 4.938988, 4.943835, 4.947769, 4.950856, 4.953206, 
    4.954986, 30, 4.965112, 4.969028, 4.974089, 4.979712, 4.985476, 4.983797, 
    4.983668, 4.983923, 4.985918, 4.989429, 4.994407, 5.000427, 5.007351, 
    5.013689, 5.020282, 5.018254, 5.014394, 5.008122, 4.998861, 4.986204, 
    4.970013, 4.950536, 4.92847, 4.904962, 4.881504, 4.859735, 4.841204, 
    4.827145, 4.818328, 4.815025, 4.817045, 4.823834, 4.834585, 4.848341,
  // totalHeight(19,26, 0-49)
    4.864459, 4.87211, 4.880964, 4.890482, 4.900172, 4.909622, 4.918519, 
    4.926631, 4.933817, 4.940006, 4.945184, 4.949382, 4.952669, 4.955164, 
    4.957052, 30, 4.968115, 4.971904, 4.97679, 4.98221, 4.987775, 4.986162, 
    4.986086, 4.986403, 4.988436, 4.991954, 4.996908, 5.002874, 5.009715, 
    5.015938, 5.022344, 5.020271, 5.016323, 5.009913, 5.00047, 4.98759, 
    4.971152, 4.951414, 4.929086, 4.905328, 4.881636, 4.859649, 4.840906, 
    4.826628, 4.817581, 4.814027, 4.815778, 4.822286, 4.832751, 4.846226,
  // totalHeight(19,27, 0-49)
    4.861812, 4.869731, 4.878926, 4.888848, 4.898993, 4.908931, 4.918322, 
    4.926916, 4.934547, 4.941125, 4.946622, 4.951062, 4.954522, 4.957128, 
    4.959073, 30, 4.97163, 4.975142, 4.979673, 4.984694, 4.989872, 4.988544, 
    4.988675, 4.989195, 4.991359, 4.994929, 4.999852, 5.005712, 5.012372, 
    5.018343, 5.024315, 5.022226, 5.018149, 5.011499, 5.001717, 4.988418, 
    4.971513, 4.951303, 4.928545, 4.904437, 4.880499, 4.858378, 4.839594, 
    4.825338, 4.816338, 4.812825, 4.814583, 4.821054, 4.831435, 4.844779,
  // totalHeight(19,28, 0-49)
    4.859741, 4.867873, 4.877347, 4.887616, 4.898163, 4.908547, 4.918406, 
    4.927459, 4.935514, 4.942453, 4.948228, 4.952856, 4.956412, 4.959038, 
    4.960937, 30, 4.975993, 4.979054, 4.983034, 4.987453, 4.992063, 4.991148, 
    4.991572, 4.99238, 4.994724, 4.998356, 5.003215, 5.008902, 5.015275, 
    5.020853, 5.026161, 5.024028, 5.019733, 5.012695, 5.002378, 4.988438, 
    4.970845, 4.949972, 4.926649, 4.90214, 4.87801, 4.8559, 4.837305, 
    4.823361, 4.814726, 4.811572, 4.813638, 4.820332, 4.830835, 4.844201,
  // totalHeight(19,29, 0-49)
    4.858432, 4.866712, 4.876399, 4.88695, 4.897851, 4.908648, 4.918948, 
    4.92844, 4.936892, 4.944144, 4.950123, 4.95483, 4.958349, 4.960835, 
    4.962511, 30, 4.980938, 4.983357, 4.986584, 4.990198, 4.994048, 4.993536, 
    4.994227, 4.995311, 4.997817, 5.001482, 5.006229, 5.011665, 5.017635, 
    5.022667, 5.027061, 5.024763, 5.020088, 5.012481, 5.00145, 4.986721, 
    4.968343, 4.946784, 4.922968, 4.898229, 4.874156, 4.852381, 4.834337, 
    4.821075, 4.813166, 4.810695, 4.81334, 4.820467, 4.831241, 4.8447,
  // totalHeight(19,30, 0-49)
    4.857325, 4.864811, 4.87362, 4.883223, 4.89315, 4.903017, 4.912543, 
    4.921545, 4.929926, 4.937651, 4.944711, 4.951098, 4.956753, 4.961548, 
    4.965257, 4.981699, 4.974598, 4.979191, 4.985151, 4.991585, 4.998013, 
    5.000706, 5.003804, 5.006528, 5.009774, 5.013294, 5.017124, 5.021049, 
    5.02509, 5.027961, 5.029866, 5.026049, 5.019855, 5.010766, 4.998342, 
    4.982376, 4.962988, 4.940724, 4.916574, 4.891904, 4.868294, 4.847318, 
    4.830311, 4.818207, 4.811459, 4.810057, 4.813608, 4.821434, 4.832671, 
    4.846352,
  // totalHeight(19,31, 0-49)
    4.858174, 4.865802, 4.874738, 4.884463, 4.894507, 4.904485, 4.9141, 
    4.923157, 4.931543, 4.939215, 4.946176, 4.952444, 4.958014, 4.962843, 
    4.966795, 4.981744, 4.976817, 4.98103, 4.986337, 4.99197, 4.997562, 
    5.000377, 5.003357, 5.005968, 5.009114, 5.01259, 5.016417, 5.020319, 
    5.02421, 5.026711, 5.027736, 5.023791, 5.017277, 5.007711, 4.994723, 
    4.978187, 4.958328, 4.935792, 4.911653, 4.88733, 4.8644, 4.844378, 
    4.828509, 4.817608, 4.812016, 4.811631, 4.815988, 4.824363, 4.835867, 
    4.849523,
  // totalHeight(19,32, 0-49)
    4.860078, 4.867659, 4.876506, 4.886116, 4.896039, 4.905897, 4.915404, 
    4.924363, 4.932662, 4.940258, 4.947163, 4.953413, 4.959052, 4.964091, 
    4.968487, 4.981169, 4.978074, 4.982155, 4.987026, 4.992065, 4.997014, 
    5.000091, 5.003103, 5.005722, 5.008819, 5.012202, 5.015869, 5.019507, 
    5.02294, 5.024753, 5.024618, 5.020299, 5.013247, 5.003031, 4.989363, 
    4.972216, 4.95193, 4.929254, 4.905345, 4.881649, 4.859718, 4.840992, 
    4.826592, 4.817206, 4.813052, 4.813928, 4.819293, 4.828377, 4.840262, 
    4.853956,
  // totalHeight(19,33, 0-49)
    4.863094, 4.870475, 4.879053, 4.888352, 4.897948, 4.907487, 4.916703, 
    4.925407, 4.9335, 4.940943, 4.947758, 4.953999, 4.959738, 4.965044, 
    4.969951, 4.980079, 4.97859, 4.982728, 4.987326, 4.991925, 4.996374, 
    4.999796, 5.002942, 5.005651, 5.008716, 5.011941, 5.015303, 5.018456, 
    5.021159, 5.022017, 5.020511, 5.015593, 5.007808, 4.996795, 4.982359, 
    4.964593, 4.943953, 4.921297, 4.897847, 4.875063, 4.854445, 4.837331, 
    4.824705, 4.817112, 4.814642, 4.816987, 4.823531, 4.833456, 4.845809, 
    4.859584,
  // totalHeight(19,34, 0-49)
    4.867206, 4.874252, 4.882409, 4.891233, 4.900333, 4.909385, 4.918148, 
    4.926455, 4.934219, 4.941414, 4.948065, 4.954243, 4.960041, 4.96557, 
    4.970939, 4.978593, 4.978584, 4.98288, 4.987299, 4.991557, 4.995606, 
    4.999401, 5.002732, 5.005574, 5.008594, 5.011591, 5.014505, 5.016977, 
    5.018713, 5.018397, 5.015368, 5.009659, 5.000988, 4.989071, 4.973829, 
    4.955482, 4.934607, 4.912163, 4.889425, 4.867839, 4.848833, 4.833615, 
    4.823024, 4.817452, 4.816856, 4.820828, 4.828676, 4.839528, 4.852401, 
    4.86627,
  // totalHeight(19,35, 0-49)
    4.872328, 4.878919, 4.886526, 4.89474, 4.903203, 4.911632, 4.919809, 
    4.927599, 4.934926, 4.941772, 4.948174, 4.954204, 4.959976, 4.965626, 
    4.971318, 4.976828, 4.978239, 4.982703, 4.986978, 4.990948, 4.99466, 
    4.998809, 5.002337, 5.005319, 5.008259, 5.010948, 5.01328, 5.014896, 
    5.015461, 5.013795, 5.009148, 5.002493, 4.992821, 4.979948, 4.963921, 
    4.945088, 4.92415, 4.90215, 4.880391, 4.860284, 4.843158, 4.83008, 
    4.821725, 4.818338, 4.819746, 4.825438, 4.834654, 4.84647, 4.859871, 
    4.873812,
  // totalHeight(19,36, 0-49)
    4.878319, 4.884347, 4.891294, 4.898786, 4.906506, 4.914204, 4.921698, 
    4.928871, 4.935667, 4.942079, 4.948146, 4.953941, 4.95958, 4.965217, 
    4.97104, 4.974863, 4.977667, 4.982239, 4.986354, 4.99006, 4.993469, 
    4.997919, 5.001616, 5.004714, 5.007523, 5.009817, 5.011443, 5.012049, 
    5.011275, 5.008129, 5.00182, 4.994109, 4.98338, 4.969563, 4.952835, 
    4.933675, 4.912894, 4.891598, 4.871095, 4.852732, 4.837718, 4.826962, 
    4.820982, 4.819872, 4.823338, 4.830776, 4.841359, 4.854115, 4.868001, 
    4.881951,
  // totalHeight(19,37, 0-49)
    4.884991, 4.890361, 4.896557, 4.903244, 4.910141, 4.917033, 4.923767, 
    4.930253, 4.936448, 4.942355, 4.948011, 4.953487, 4.958893, 4.964376, 
    4.97013, 4.972736, 4.976905, 4.981477, 4.985387, 4.988821, 4.991942, 
    4.996607, 5.000417, 5.003583, 5.006192, 5.008002, 5.008813, 5.008285, 
    5.006043, 5.001339, 4.993384, 4.98456, 4.972786, 4.958107, 4.940834, 
    4.921567, 4.901206, 4.880898, 4.861922, 4.845537, 4.832814, 4.824502, 
    4.820959, 4.822139, 4.827637, 4.836768, 4.848647, 4.862257, 4.876529, 
    4.890384,
  // totalHeight(19,38, 0-49)
    4.892121, 4.896754, 4.902132, 4.907953, 4.913973, 4.920011, 4.92594, 
    4.931687, 4.937231, 4.942576, 4.947761, 4.952847, 4.957928, 4.963131, 
    4.968633, 4.970451, 4.975925, 4.980362, 4.984005, 4.987148, 4.989974, 
    4.994747, 4.99859, 5.001753, 5.004083, 5.005324, 5.005226, 5.003472, 
    4.999688, 4.993407, 4.983876, 4.973956, 4.96122, 4.945838, 4.928244, 
    4.909145, 4.889503, 4.870472, 4.853275, 4.839058, 4.828744, 4.82292, 
    4.821793, 4.825191, 4.832617, 4.843311, 4.856339, 4.870652, 4.885157, 
    4.898771,
  // totalHeight(19,39, 0-49)
    4.899467, 4.903297, 4.907806, 4.912726, 4.917843, 4.923001, 4.928099, 
    4.933086, 4.937946, 4.942693, 4.947358, 4.951997, 4.95668, 4.961504, 
    4.966603, 4.967971, 4.974646, 4.978811, 4.982118, 4.984936, 4.987445, 
    4.992202, 4.995981, 4.999056, 5.00102, 5.001617, 5.000542, 4.997513, 
    4.99217, 4.984358, 4.973391, 4.962465, 4.948932, 4.93308, 4.915452, 
    4.896836, 4.878227, 4.860754, 4.845551, 4.833638, 4.825777, 4.822405, 
    4.823591, 4.829056, 4.838219, 4.850267, 4.864228, 4.879025, 4.893557, 
    4.906746,
  // totalHeight(19,40, 0-49)
    4.906766, 4.909746, 4.913357, 4.917359, 4.921566, 4.925843, 4.930111, 
    4.934331, 4.938495, 4.942622, 4.94674, 4.950891, 4.95512, 4.959492, 
    4.964085, 4.965239, 4.97296, 4.976724, 4.979627, 4.98208, 4.984232, 
    4.988842, 4.992447, 4.995337, 4.996855, 4.996744, 4.994654, 4.990354, 
    4.983506, 4.974283, 4.962084, 4.950325, 4.936236, 4.920212, 4.902885, 
    4.885092, 4.867829, 4.852161, 4.839121, 4.829577, 4.824143, 4.823107, 
    4.82642, 4.833713, 4.844347, 4.857467, 4.872072, 4.887079, 4.901387, 
    4.913939,
  // totalHeight(19,41, 0-49)
    4.913755, 4.915848, 4.918544, 4.921631, 4.924941, 4.928359, 4.931815, 
    4.935283, 4.938761, 4.942267, 4.945827, 4.949466, 4.953209, 4.957081, 
    4.961106, 4.962186, 4.970744, 4.974006, 4.976444, 4.97848, 4.980226, 
    4.984553, 4.987868, 4.990473, 4.991469, 4.990608, 4.987513, 4.982002, 
    4.973772, 4.963334, 4.950175, 4.93783, 4.923496, 4.90765, 4.890987, 
    4.874359, 4.858728, 4.845076, 4.8343, 4.827125, 4.824011, 4.825119, 
    4.830297, 4.839108, 4.850871, 4.864708, 4.879611, 4.894502, 4.908296, 
    4.919983,
  // totalHeight(19,42, 0-49)
    4.92017, 4.921348, 4.923127, 4.925314, 4.927758, 4.930353, 4.933038, 
    4.935792, 4.938614, 4.94152, 4.944527, 4.94765, 4.950894, 4.954247, 
    4.957675, 4.958741, 4.967895, 4.970575, 4.972492, 4.974058, 4.975332, 
    4.979243, 4.982157, 4.984379, 4.984793, 4.983174, 4.979122, 4.97252, 
    4.963109, 4.951718, 4.937935, 4.92532, 4.911098, 4.895811, 4.880182, 
    4.865045, 4.851295, 4.839802, 4.83133, 4.826448, 4.825478, 4.828466, 
    4.835182, 4.845138, 4.857627, 4.871772, 4.886574, 4.900981, 4.913953, 
    4.924549,
  // totalHeight(19,43, 0-49)
    4.925763, 4.926003, 4.926868, 4.928182, 4.929801, 4.931626, 4.933599, 
    4.935696, 4.937914, 4.94026, 4.942748, 4.945375, 4.948125, 4.950956, 
    4.953793, 4.954841, 4.96433, 4.966375, 4.967723, 4.968758, 4.969495, 
    4.972867, 4.975272, 4.977025, 4.97682, 4.974465, 4.969556, 4.962043, 
    4.951717, 4.939699, 4.925668, 4.913147, 4.899427, 4.885087, 4.87084, 
    4.857475, 4.845798, 4.836551, 4.830351, 4.827622, 4.828561, 4.833115, 
    4.840987, 4.851663, 4.86443, 4.878427, 4.892694, 4.906231, 4.91807, 
    4.927366,
  // totalHeight(19,44, 0-49)
    4.930317, 4.929597, 4.929554, 4.930022, 4.930867, 4.931989, 4.933323, 
    4.934839, 4.936524, 4.938376, 4.940395, 4.942565, 4.944849, 4.94718, 
    4.949445, 4.950438, 4.960001, 4.961379, 4.962115, 4.96256, 4.962694, 
    4.965418, 4.967226, 4.968439, 4.967605, 4.964572, 4.95895, 4.950758, 
    4.93984, 4.927562, 4.913687, 4.901648, 4.888824, 4.875793, 4.863242, 
    4.85188, 4.842403, 4.835417, 4.831395, 4.830625, 4.833188, 4.838951, 
    4.847569, 4.85851, 4.87108, 4.884458, 4.897746, 4.910027, 4.920442, 
    4.928277,
  // totalHeight(19,45, 0-49)
    4.933671, 4.931966, 4.931014, 4.930665, 4.930786, 4.931273, 4.932052, 
    4.933077, 4.934319, 4.935762, 4.937385, 4.939156, 4.941019, 4.942884, 
    4.944615, 4.945492, 4.954885, 4.955587, 4.955676, 4.955476, 4.954947, 
    4.956939, 4.958081, 4.958708, 4.957262, 4.953647, 4.947495, 4.938894, 
    4.92774, 4.915594, 4.902283, 4.89111, 4.879552, 4.868159, 4.857555, 
    4.848358, 4.841139, 4.836369, 4.834379, 4.835332, 4.839209, 4.845804, 
    4.854742, 4.86549, 4.877389, 4.889682, 4.901563, 4.912237, 4.920988, 
    4.927265,
  // totalHeight(19,46, 0-49)
    4.935753, 4.933025, 4.931156, 4.930007, 4.929449, 4.929368, 4.929675, 
    4.930304, 4.931202, 4.932328, 4.933641, 4.935088, 4.936592, 4.938042, 
    4.939281, 4.939974, 4.948993, 4.949016, 4.948432, 4.947545, 4.946309, 
    4.947513, 4.947949, 4.947968, 4.945961, 4.941886, 4.935413, 4.926697, 
    4.915676, 4.904049, 4.89169, 4.881741, 4.871771, 4.862283, 4.853815, 
    4.846878, 4.841915, 4.83926, 4.839114, 4.841527, 4.846392, 4.853445, 
    4.862292, 4.872415, 4.883203, 4.893989, 4.904093, 4.912873, 4.919795, 
    4.924508,
  // totalHeight(19,47, 0-49)
    4.936611, 4.932811, 4.929999, 4.92805, 4.926839, 4.926242, 4.92615, 
    4.92647, 4.927119, 4.928027, 4.929121, 4.930323, 4.931534, 4.932622, 
    4.93342, 4.933862, 4.942347, 4.941703, 4.94043, 4.938825, 4.936858, 
    4.937251, 4.936972, 4.936396, 4.933905, 4.929514, 4.922946, 4.914406, 
    4.903878, 4.893131, 4.882066, 4.873648, 4.86553, 4.858142, 4.851929, 
    4.847281, 4.844512, 4.843832, 4.84532, 4.848924, 4.854459, 4.861622, 
    4.870004, 4.879118, 4.888425, 4.897368, 4.905418, 4.912122, 4.917159, 
    4.920394,
  // totalHeight(19,48, 0-49)
    4.936437, 4.931505, 4.927708, 4.924939, 4.923077, 4.921989, 4.921544, 
    4.921619, 4.922096, 4.922868, 4.923826, 4.924857, 4.925838, 4.926618, 
    4.92702, 4.927145, 4.934983, 4.93369, 4.931725, 4.929393, 4.926692, 
    4.926288, 4.925319, 4.924188, 4.921313, 4.916768, 4.910326, 4.90224, 
    4.892526, 4.88297, 4.87348, 4.866836, 4.860761, 4.855598, 4.851686, 
    4.849298, 4.848623, 4.849751, 4.852652, 4.857186, 4.863106, 4.870075, 
    4.877688, 4.885501, 4.89306, 4.89994, 4.905788, 4.910366, 4.913583, 
    4.915535,
  // totalHeight(19,49, 0-49)
    4.939479, 4.932686, 4.927199, 4.922946, 4.919828, 4.917706, 4.916431, 
    4.915837, 4.915757, 4.916022, 4.916465, 4.916909, 4.91717, 4.917032, 
    4.916247, 4.915366, 4.929752, 4.926197, 4.921779, 4.917198, 4.912539, 
    4.913105, 4.913378, 4.914213, 4.912521, 4.90855, 4.901885, 4.89297, 
    4.881677, 4.871408, 4.861761, 4.857852, 4.85482, 4.852896, 4.852281, 
    4.853092, 4.855345, 4.858965, 4.86378, 4.869527, 4.875886, 4.882484, 
    4.888945, 4.894903, 4.900057, 4.904189, 4.907223, 4.909227, 4.910436, 
    4.91124,
  // totalHeight(20,0, 0-49)
    4.860252, 4.86001, 4.861908, 4.865577, 4.870636, 4.876714, 4.883478, 
    4.890644, 4.897981, 4.905314, 4.912512, 4.919477, 4.926129, 4.932405, 
    4.938227, 4.943402, 4.949084, 4.953224, 4.956752, 4.959602, 4.961658, 
    4.963098, 4.963417, 4.962541, 4.960215, 4.956271, 4.950531, 4.9429, 
    4.933327, 4.921966, 4.908915, 4.894793, 4.879703, 4.864185, 4.848875, 
    4.834458, 4.821619, 4.810974, 4.803027, 4.798102, 4.796328, 4.797613, 
    4.801653, 4.80796, 4.815895, 4.82473, 4.833702, 4.842091, 4.849298, 
    4.854918,
  // totalHeight(20,1, 0-49)
    4.862436, 4.862621, 4.86489, 4.86887, 4.874181, 4.880456, 4.887374, 
    4.894657, 4.902087, 4.909499, 4.91677, 4.923805, 4.93053, 4.936876, 
    4.94276, 4.947818, 4.954359, 4.958505, 4.962062, 4.965001, 4.967188, 
    4.969077, 4.969801, 4.969337, 4.967341, 4.963618, 4.957946, 4.950209, 
    4.94033, 4.92852, 4.914805, 4.900119, 4.884272, 4.867824, 4.851451, 
    4.835898, 4.821912, 4.810189, 4.8013, 4.795636, 4.793375, 4.794456, 
    4.798588, 4.805271, 4.813842, 4.823527, 4.833501, 4.842969, 4.851245, 
    4.857827,
  // totalHeight(20,2, 0-49)
    4.864428, 4.86499, 4.867573, 4.871808, 4.877315, 4.883739, 4.890766, 
    4.898131, 4.905627, 4.913094, 4.920412, 4.927494, 4.934264, 4.94065, 
    4.946568, 4.951439, 4.958696, 4.962821, 4.966372, 4.969354, 4.971641, 
    4.973957, 4.97509, 4.97507, 4.97349, 4.970134, 4.964743, 4.957186, 
    4.947346, 4.935463, 4.921481, 4.90663, 4.890397, 4.873343, 4.856158, 
    4.839617, 4.824526, 4.811648, 4.801634, 4.794953, 4.791851, 4.792322, 
    4.79611, 4.802735, 4.811536, 4.821715, 4.832422, 4.842813, 4.852137, 
    4.85981,
  // totalHeight(20,3, 0-49)
    4.866155, 4.86705, 4.869899, 4.874338, 4.879996, 4.886528, 4.893631, 
    4.90105, 4.908585, 4.916081, 4.923425, 4.930527, 4.937315, 4.943715, 
    4.949641, 4.954255, 4.962042, 4.966132, 4.969641, 4.972626, 4.974976, 
    4.977679, 4.979204, 4.979639, 4.978534, 4.975669, 4.970754, 4.963642, 
    4.954173, 4.94259, 4.928738, 4.914125, 4.897903, 4.880599, 4.862891, 
    4.845562, 4.829454, 4.815392, 4.804106, 4.796156, 4.791875, 4.791333, 
    4.794338, 4.800455, 4.809047, 4.819333, 4.830458, 4.841559, 4.851843, 
    4.860661,
  // totalHeight(20,4, 0-49)
    4.867635, 4.868824, 4.871896, 4.876496, 4.882263, 4.888866, 4.896011, 
    4.903454, 4.910999, 4.918499, 4.925837, 4.932927, 4.939702, 4.946087, 
    4.952006, 4.956291, 4.964385, 4.968431, 4.971873, 4.974825, 4.977198, 
    4.980241, 4.982126, 4.982999, 4.982406, 4.980123, 4.975844, 4.969408, 
    4.960617, 4.949678, 4.936331, 4.922343, 4.906526, 4.889344, 4.871434, 
    4.85356, 4.836578, 4.82136, 4.808711, 4.799289, 4.793529, 4.791602, 
    4.793405, 4.798576, 4.80653, 4.816529, 4.827738, 4.8393, 4.850401, 
    4.860345,
  // totalHeight(20,5, 0-49)
    4.868941, 4.870391, 4.873652, 4.878376, 4.884216, 4.890854, 4.898007, 
    4.905436, 4.912956, 4.920418, 4.927711, 4.934752, 4.941473, 4.947814, 
    4.953711, 4.957606, 4.965757, 4.969759, 4.973117, 4.976005, 4.978372, 
    4.981693, 4.983891, 4.98517, 4.985097, 4.983453, 4.979932, 4.97436, 
    4.966503, 4.956503, 4.944001, 4.930983, 4.915935, 4.899241, 4.881466, 
    4.863327, 4.845665, 4.82938, 4.815343, 4.80431, 4.796834, 4.793207, 
    4.793438, 4.797264, 4.804183, 4.813521, 4.824488, 4.836249, 4.84799, 
    4.858978,
  // totalHeight(20,6, 0-49)
    4.870184, 4.871867, 4.875287, 4.880104, 4.885983, 4.892617, 4.899735, 
    4.907109, 4.914557, 4.921935, 4.929136, 4.936078, 4.942703, 4.948964, 
    4.95482, 4.958287, 4.966236, 4.970192, 4.97346, 4.976264, 4.978598, 
    4.982133, 4.984593, 4.986225, 4.986656, 4.985677, 4.982993, 4.978419, 
    4.971696, 4.962874, 4.95149, 4.939726, 4.925767, 4.9099, 4.892593, 
    4.874488, 4.856383, 4.83918, 4.823804, 4.8111, 4.801749, 4.796178, 
    4.794536, 4.796683, 4.802223, 4.810569, 4.820991, 4.832695, 4.844877, 
    4.856782,
  // totalHeight(20,7, 0-49)
    4.871486, 4.873385, 4.876938, 4.881816, 4.887699, 4.894289, 4.901329, 
    4.908598, 4.915922, 4.923161, 4.930209, 4.936997, 4.943477, 4.949618, 
    4.955414, 4.958443, 4.965936, 4.969844, 4.97302, 4.975732, 4.978019, 
    4.981705, 4.984363, 4.986288, 4.987187, 4.986865, 4.985055, 4.981565, 
    4.976113, 4.968638, 4.958585, 4.948279, 4.935663, 4.92091, 4.904378, 
    4.886606, 4.868324, 4.850407, 4.833809, 4.819458, 4.808159, 4.800493, 
    4.796761, 4.796972, 4.800858, 4.807934, 4.81755, 4.828959, 4.841378, 
    4.854039,
  // totalHeight(20,8, 0-49)
    4.872965, 4.875064, 4.878729, 4.883643, 4.889493, 4.895999, 4.902913, 
    4.910024, 4.917163, 4.924199, 4.931038, 4.937615, 4.943896, 4.949877, 
    4.955583, 4.958203, 4.965009, 4.968857, 4.971947, 4.974571, 4.976808, 
    4.980578, 4.983373, 4.98552, 4.986834, 4.987137, 4.986202, 4.983829, 
    4.979728, 4.973704, 4.965117, 4.956395, 4.945295, 4.931881, 4.916384, 
    4.899226, 4.88104, 4.862648, 4.845007, 4.829113, 4.815887, 4.806065, 
    4.800118, 4.798223, 4.800258, 4.805854, 4.81445, 4.825356, 4.837813, 
    4.851048,
  // totalHeight(20,9, 0-49)
    4.874715, 4.877008, 4.88077, 4.885693, 4.891478, 4.897859, 4.904594, 
    4.911492, 4.918387, 4.925161, 4.931726, 4.938032, 4.944063, 4.949836, 
    4.955409, 4.957707, 4.963628, 4.967393, 4.970406, 4.972955, 4.975152, 
    4.978941, 4.981811, 4.984108, 4.985774, 4.98665, 4.986557, 4.985291, 
    4.982565, 4.978032, 4.970989, 4.96389, 4.954402, 4.942473, 4.928211, 
    4.911908, 4.894079, 4.87547, 4.857014, 4.839749, 4.824699, 4.812755, 
    4.804565, 4.800483, 4.800548, 4.804519, 4.811933, 4.82216, 4.834473, 
    4.848091,
  // totalHeight(20,10, 0-49)
    4.876799, 4.879285, 4.883133, 4.888045, 4.893735, 4.899947, 4.906461, 
    4.913087, 4.919682, 4.926131, 4.932365, 4.938345, 4.944074, 4.949587, 
    4.954967, 4.957089, 4.961978, 4.965627, 4.968569, 4.971067, 4.973243, 
    4.97699, 4.979874, 4.98225, 4.984199, 4.985584, 4.986276, 4.986076, 
    4.984701, 4.981645, 4.976162, 4.970654, 4.962789, 4.952418, 4.939521, 
    4.924259, 4.907021, 4.88845, 4.869433, 4.851023, 4.834328, 4.82038, 
    4.810005, 4.803736, 4.801787, 4.804056, 4.810177, 4.819589, 4.831591, 
    4.845403,
  // totalHeight(20,11, 0-49)
    4.879239, 4.881923, 4.885851, 4.890735, 4.896304, 4.902315, 4.908561, 
    4.91487, 4.921111, 4.927186, 4.933039, 4.938643, 4.944018, 4.949213, 
    4.954324, 4.956469, 4.960239, 4.963728, 4.966609, 4.969083, 4.971266, 
    4.974913, 4.977757, 4.980145, 4.982306, 4.984129, 4.985535, 4.986328, 
    4.986242, 4.98461, 4.980663, 4.976647, 4.97035, 4.961532, 4.950062, 
    4.935967, 4.919504, 4.901208, 4.881889, 4.862591, 4.844482, 4.828718, 
    4.816289, 4.807916, 4.80398, 4.804524, 4.80929, 4.81778, 4.829328, 
    4.843155,
  // totalHeight(20,12, 0-49)
    4.88201, 4.884904, 4.888915, 4.893763, 4.899191, 4.904974, 4.910917, 
    4.916871, 4.922716, 4.928374, 4.933802, 4.938989, 4.943964, 4.948782, 
    4.953533, 4.95595, 4.958569, 4.961857, 4.964685, 4.967168, 4.969397, 
    4.972889, 4.975645, 4.977991, 4.980297, 4.982482, 4.984518, 4.986214, 
    4.987322, 4.987028, 4.984559, 4.981891, 4.977048, 4.969718, 4.959666, 
    4.946801, 4.93125, 4.913426, 4.894051, 4.874133, 4.854875, 4.837531, 
    4.823242, 4.812902, 4.807063, 4.805912, 4.809299, 4.816798, 4.827771, 
    4.841449,
  // totalHeight(20,13, 0-49)
    4.885045, 4.888165, 4.892267, 4.897079, 4.902358, 4.907895, 4.913514, 
    4.919086, 4.924509, 4.929721, 4.934696, 4.939434, 4.943967, 4.948348, 
    4.952642, 4.955595, 4.957088, 4.960145, 4.962937, 4.965468, 4.967791, 
    4.971079, 4.973709, 4.975964, 4.978357, 4.980833, 4.98341, 4.985902, 
    4.98809, 4.989025, 4.987952, 4.986454, 4.982911, 4.976952, 4.968254, 
    4.956622, 4.942061, 4.92486, 4.905646, 4.885368, 4.865235, 4.846574, 
    4.830656, 4.818532, 4.810918, 4.808143, 4.810166, 4.816629, 4.826932, 
    4.840311,
  // totalHeight(20,14, 0-49)
    4.888229, 4.8916, 4.895807, 4.900593, 4.905726, 4.911015, 4.916304, 
    4.921482, 4.92647, 4.931225, 4.935732, 4.940003, 4.944067, 4.947958, 
    4.951711, 4.955437, 4.955875, 4.958696, 4.961479, 4.964108, 4.966577, 
    4.969624, 4.9721, 4.974234, 4.976667, 4.979364, 4.98239, 4.985562, 
    4.988698, 4.990733, 4.990968, 4.99044, 4.988013, 4.983267, 4.975816, 
    4.965367, 4.951819, 4.935346, 4.916467, 4.896061, 4.875321, 4.855616, 
    4.838318, 4.824619, 4.815388, 4.811089, 4.811786, 4.817195, 4.826753, 
    4.839705,
  // totalHeight(20,15, 0-49)
    4.891417, 4.895063, 4.899403, 4.904181, 4.909182, 4.914233, 4.919199, 
    4.923991, 4.928551, 4.932856, 4.936903, 4.940707, 4.944289, 4.947664, 
    4.950818, 4.955467, 4.954948, 4.957564, 4.96039, 4.963179, 4.965862, 
    4.968639, 4.970955, 4.972952, 4.975391, 4.978249, 4.981628, 4.985358, 
    4.989294, 4.99229, 4.993727, 4.993963, 4.99245, 4.988739, 4.982389, 
    4.973036, 4.96048, 4.944787, 4.926372, 4.906035, 4.884928, 4.864438, 
    4.846014, 4.830963, 4.820285, 4.814578, 4.81401, 4.818363, 4.827119, 
    4.839538,
  // totalHeight(20,16, 0-49)
    4.894438, 4.898385, 4.902883, 4.90768, 4.912577, 4.917415, 4.922084, 
    4.926518, 4.93068, 4.934565, 4.938181, 4.941544, 4.944665, 4.94753, 
    4.950081, 4.955651, 4.954271, 4.956758, 4.959707, 4.962741, 4.965721, 
    4.968219, 4.970386, 4.972255, 4.974681, 4.977648, 4.981289, 4.985443, 
    4.990022, 4.993821, 4.99635, 4.997137, 4.996331, 4.993463, 4.98805, 
    4.97967, 4.968042, 4.953138, 4.935272, 4.915156, 4.893888, 4.87285, 
    4.853538, 4.837351, 4.825407, 4.818417, 4.816652, 4.819967, 4.827884, 
    4.839682,
  // totalHeight(20,17, 0-49)
    4.897111, 4.901378, 4.906057, 4.910903, 4.915725, 4.920388, 4.924805, 
    4.92893, 4.93275, 4.936276, 4.939528, 4.942516, 4.945239, 4.947652, 
    4.949658, 4.955938, 4.95375, 4.956237, 4.959424, 4.962814, 4.966193, 
    4.968428, 4.970485, 4.972262, 4.974679, 4.977714, 4.981524, 4.985966, 
    4.991012, 4.995444, 4.99893, 5.000061, 4.999754, 4.997528, 4.992876, 
    4.985324, 4.974533, 4.960389, 4.943113, 4.92333, 4.90207, 4.880688, 
    4.860705, 4.843585, 4.830546, 4.822402, 4.819518, 4.82182, 4.828876, 
    4.839989,
  // totalHeight(20,18, 0-49)
    4.899259, 4.903844, 4.908713, 4.913628, 4.918412, 4.922945, 4.927167, 
    4.931057, 4.934627, 4.9379, 4.940901, 4.943637, 4.946083, 4.948168, 
    4.94976, 4.956294, 4.953275, 4.955921, 4.959491, 4.963376, 4.967283, 
    4.969299, 4.971318, 4.973071, 4.97551, 4.97859, 4.98248, 4.987064, 
    4.992386, 4.997256, 5.001545, 5.002809, 5.002788, 5.001004, 4.996927, 
    4.990052, 4.979986, 4.966546, 4.949867, 4.930487, 4.909364, 4.887812, 
    4.867347, 4.849483, 4.83551, 4.826337, 4.822413, 4.823737, 4.829926, 
    4.840314,
  // totalHeight(20,19, 0-49)
    4.900722, 4.905582, 4.910621, 4.915603, 4.920366, 4.924819, 4.928921, 
    4.932685, 4.936142, 4.939328, 4.942264, 4.944942, 4.947306, 4.949254, 
    4.950626, 4.956723, 4.952731, 4.955709, 4.959822, 4.964365, 4.968961, 
    4.970843, 4.972939, 4.974776, 4.977301, 4.980426, 4.984317, 4.988889, 
    4.994273, 4.99935, 5.004237, 5.005415, 5.005468, 5.00392, 5.000231, 
    4.993872, 4.984408, 4.971598, 4.9555, 4.936566, 4.915679, 4.894096, 
    4.873318, 4.854876, 4.840123, 4.83004, 4.825162, 4.825555, 4.830888, 
    4.840529,
  // totalHeight(20,20, 0-49)
    4.90239, 4.908547, 4.914843, 4.921025, 4.926898, 4.932327, 4.937214, 
    4.9415, 4.945158, 4.948183, 4.950596, 4.952441, 4.953793, 4.954744, 
    4.955407, 30, 4.958249, 4.960236, 4.962961, 4.965996, 4.969181, 4.968955, 
    4.969491, 4.97025, 4.972277, 4.975456, 4.979868, 4.985317, 4.991841, 
    4.998215, 5.004694, 5.006587, 5.007314, 5.006402, 5.00332, 4.997553, 
    4.988664, 4.976397, 4.960779, 4.942212, 4.921516, 4.899904, 4.878851, 
    4.859899, 4.844436, 4.83351, 4.827723, 4.827208, 4.831687, 4.840559,
  // totalHeight(20,21, 0-49)
    4.902546, 4.909152, 4.915813, 4.922264, 4.928308, 4.93382, 4.938725, 
    4.942987, 4.946609, 4.949608, 4.952027, 4.953918, 4.955361, 4.956449, 
    4.957307, 30, 4.95625, 4.958742, 4.96202, 4.965616, 4.96931, 4.968532, 
    4.968688, 4.969118, 4.970976, 4.974154, 4.978734, 4.984498, 4.991485, 
    4.998459, 5.005868, 5.007966, 5.009057, 5.008655, 5.006201, 5.001147, 
    4.99302, 4.981514, 4.966591, 4.948582, 4.928237, 4.906707, 4.885434, 
    4.865964, 4.849724, 4.837832, 4.830966, 4.829334, 4.832719, 4.840568,
  // totalHeight(20,22, 0-49)
    4.902033, 4.909122, 4.916215, 4.92303, 4.929366, 4.935092, 4.940144, 
    4.944501, 4.948182, 4.951223, 4.953678, 4.955619, 4.957127, 4.958311, 
    4.959311, 30, 4.955119, 4.958027, 4.96179, 4.965904, 4.970087, 4.968813, 
    4.968649, 4.968804, 4.970531, 4.973706, 4.978404, 4.984384, 4.991682, 
    4.999045, 5.007104, 5.009167, 5.010358, 5.010189, 5.00809, 5.003501, 
    4.995925, 4.985018, 4.970692, 4.953214, 4.933263, 4.911923, 4.89059, 
    4.870792, 4.853981, 4.841319, 4.833551, 4.830953, 4.833365, 4.84028,
  // totalHeight(20,23, 0-49)
    4.900946, 4.908532, 4.916096, 4.92334, 4.930048, 4.936085, 4.941385, 
    4.945931, 4.949752, 4.952897, 4.955433, 4.95744, 4.959013, 4.96027, 
    4.961375, 30, 4.954969, 4.958154, 4.962238, 4.966699, 4.971208, 4.969459, 
    4.96897, 4.968847, 4.970413, 4.973536, 4.978281, 4.984387, 4.991886, 
    4.999502, 5.008006, 5.009949, 5.011131, 5.011066, 5.009185, 5.00492, 
    4.99776, 4.987338, 4.973525, 4.956533, 4.936977, 4.915878, 4.894584, 
    4.874597, 4.857371, 4.844103, 4.835588, 4.832156, 4.833704, 4.839765,
  // totalHeight(20,24, 0-49)
    4.899428, 4.907504, 4.915555, 4.92326, 4.930388, 4.936795, 4.942407, 
    4.947209, 4.951232, 4.95453, 4.957183, 4.959279, 4.96092, 4.962241, 
    4.963425, 30, 4.95597, 4.959291, 4.963529, 4.968157, 4.972827, 4.970741, 
    4.970021, 4.969701, 4.971145, 4.974215, 4.978966, 4.985128, 4.992729, 
    5.000482, 5.009243, 5.011076, 5.012208, 5.012159, 5.010361, 5.006243, 
    4.999289, 4.98912, 4.975582, 4.958858, 4.939522, 4.918553, 4.897259, 
    4.877122, 4.859592, 4.845881, 4.836812, 4.832757, 4.833642, 4.839036,
  // totalHeight(20,25, 0-49)
    4.897653, 4.906196, 4.91472, 4.922887, 4.93045, 4.937253, 4.943209, 
    4.948304, 4.952564, 4.956049, 4.958841, 4.961037, 4.962751, 4.964127, 
    4.965363, 30, 4.957728, 4.961046, 4.96527, 4.969884, 4.974544, 4.972311, 
    4.971497, 4.971106, 4.972506, 4.975554, 4.980302, 4.986476, 4.994102, 
    5.001885, 5.010712, 5.012488, 5.013579, 5.013506, 5.011698, 5.007585, 
    5.000655, 4.990522, 4.977032, 4.960351, 4.941041, 4.920062, 4.898702, 
    4.878432, 4.860693, 4.846697, 4.837277, 4.832819, 4.833266, 4.838201,
  // totalHeight(20,26, 0-49)
    4.895818, 4.904783, 4.913742, 4.922344, 4.930325, 4.937515, 4.943821, 
    4.949216, 4.953726, 4.957407, 4.960343, 4.962636, 4.964409, 4.965817, 
    4.967063, 30, 4.960133, 4.963308, 4.967357, 4.971776, 4.976251, 4.974082, 
    4.973327, 4.973009, 4.974462, 4.977538, 4.982289, 4.98844, 4.996022, 
    5.003737, 5.012439, 5.014235, 5.015309, 5.015183, 5.013282, 5.009041, 
    5.001948, 4.99163, 4.97794, 4.961062, 4.941566, 4.920424, 4.898925, 
    4.878536, 4.860688, 4.846581, 4.837034, 4.832421, 4.832682, 4.8374,
  // totalHeight(20,27, 0-49)
    4.894114, 4.903435, 4.912771, 4.921757, 4.930116, 4.937665, 4.944301, 
    4.949985, 4.954732, 4.958596, 4.961658, 4.964022, 4.965817, 4.967206, 
    4.968397, 30, 4.96324, 4.966122, 4.969824, 4.973864, 4.97798, 4.976048, 
    4.975473, 4.975338, 4.976915, 4.98005, 4.984796, 4.990885, 4.998345, 
    5.00589, 5.014274, 5.016143, 5.01721, 5.016988, 5.014902, 5.010391, 
    5.002958, 4.992247, 4.978143, 4.960862, 4.941015, 4.919603, 4.897938, 
    4.87749, 4.859674, 4.845661, 4.836235, 4.831735, 4.832074, 4.836821,
  // totalHeight(20,28, 0-49)
    4.892716, 4.902316, 4.911954, 4.921258, 4.92994, 4.937809, 4.94474, 
    4.950686, 4.955645, 4.959659, 4.962801, 4.965176, 4.966919, 4.9682, 
    4.969231, 30, 4.967395, 4.969824, 4.972999, 4.976473, 4.980055, 4.978459, 
    4.97812, 4.978223, 4.979947, 4.983134, 4.987837, 4.993802, 5.001053, 
    5.008318, 5.016205, 5.018162, 5.019183, 5.018777, 5.016371, 5.011417, 
    5.00344, 4.992121, 4.977393, 4.95953, 4.939205, 4.917471, 4.895676, 
    4.875288, 4.8577, 4.844033, 4.835011, 4.830916, 4.831614, 4.836638,
  // totalHeight(20,29, 0-49)
    4.891768, 4.901561, 4.91142, 4.920973, 4.929929, 4.938075, 4.945275, 
    4.951451, 4.956579, 4.960682, 4.963824, 4.966108, 4.967679, 4.968717, 
    4.969442, 30, 4.972353, 4.974166, 4.976633, 4.979355, 4.982222, 4.980926, 
    4.980772, 4.981068, 4.982892, 4.986081, 4.990681, 4.996451, 5.003397, 
    5.010265, 5.017463, 5.019434, 5.020311, 5.019595, 5.016734, 5.011202, 
    5.002559, 4.990538, 4.975133, 4.956691, 4.935954, 4.914032, 4.892297, 
    4.872213, 4.855128, 4.842093, 4.833755, 4.830319, 4.831594, 4.837072,
  // totalHeight(20,30, 0-49)
    4.890552, 4.899473, 4.908428, 4.917069, 4.925149, 4.932522, 4.939125, 
    4.94497, 4.950115, 4.954631, 4.958583, 4.961999, 4.964857, 4.967066, 
    4.968472, 4.979602, 4.96907, 4.971892, 4.976008, 4.980648, 4.98542, 
    4.986781, 4.988743, 4.990612, 4.993301, 4.996634, 5.000715, 5.005429, 
    5.010921, 5.01609, 5.021275, 5.022079, 5.021772, 5.019878, 5.015864, 
    5.009229, 4.99956, 4.986626, 4.970476, 4.951515, 4.930534, 4.90868, 
    4.887331, 4.867914, 4.851709, 4.839678, 4.832371, 4.829907, 4.832027, 
    4.838179,
  // totalHeight(20,31, 0-49)
    4.890921, 4.899925, 4.908952, 4.91766, 4.925797, 4.93321, 4.939828, 
    4.945653, 4.950732, 4.95514, 4.958956, 4.962236, 4.965003, 4.967213, 
    4.968752, 4.979363, 4.971177, 4.97361, 4.977141, 4.98109, 4.985148, 
    4.986675, 4.988585, 4.990395, 4.993023, 4.996342, 5.00046, 5.005226, 
    5.010689, 5.015679, 5.020274, 5.021196, 5.02085, 5.01876, 5.014407, 
    5.007318, 4.997122, 4.983652, 4.967027, 4.947731, 4.926632, 4.904924, 
    4.883998, 4.865252, 4.849897, 4.83881, 4.832448, 4.830843, 4.833675, 
    4.840341,
  // totalHeight(20,32, 0-49)
    4.891858, 4.900726, 4.909607, 4.918174, 4.926184, 4.933486, 4.940012, 
    4.945757, 4.950766, 4.955113, 4.958885, 4.962158, 4.964985, 4.967364, 
    4.969228, 4.978518, 4.972463, 4.974708, 4.977826, 4.98125, 4.984755, 
    4.986572, 4.988569, 4.990442, 4.993085, 4.996394, 5.000472, 5.005139, 
    5.010365, 5.014951, 5.01875, 5.019603, 5.019039, 5.016583, 5.011744, 
    5.004078, 4.993276, 4.979236, 4.962163, 4.942626, 4.921564, 4.900208, 
    4.879947, 4.86213, 4.847888, 4.837993, 4.832799, 4.832254, 4.835965, 
    4.843286,
  // totalHeight(20,33, 0-49)
    4.893402, 4.901961, 4.910522, 4.918782, 4.926514, 4.933579, 4.93991, 
    4.945505, 4.950407, 4.954688, 4.958445, 4.961763, 4.964719, 4.96735, 
    4.96964, 4.977197, 4.973083, 4.975312, 4.978167, 4.981205, 4.984287, 
    4.986477, 4.98866, 4.990693, 4.993394, 4.996678, 5.000629, 5.005051, 
    5.009844, 5.013827, 5.016671, 5.017282, 5.016326, 5.013347, 5.00788, 
    4.999536, 4.988063, 4.973445, 4.955978, 4.936319, 4.915467, 4.894683, 
    4.87533, 4.858694, 4.845803, 4.83732, 4.833489, 4.834168, 4.838899, 
    4.846986,
  // totalHeight(20,34, 0-49)
    4.89555, 4.903658, 4.911766, 4.919588, 4.926923, 4.933646, 4.939695, 
    4.945072, 4.949821, 4.954011, 4.957741, 4.961105, 4.964197, 4.967091, 
    4.969819, 4.975549, 4.97322, 4.975553, 4.978248, 4.981001, 4.983756, 
    4.986354, 4.988786, 4.991036, 4.993814, 4.997042, 5.000778, 5.004812, 
    5.008993, 5.012204, 5.01397, 5.014173, 5.01267, 5.009023, 5.002813, 
    4.993709, 4.981535, 4.966369, 4.9486, 4.928967, 4.908524, 4.88854, 
    4.870338, 4.855117, 4.843793, 4.836905, 4.834589, 4.836618, 4.842463, 
    4.851387,
  // totalHeight(20,35, 0-49)
    4.898267, 4.905814, 4.913355, 4.920641, 4.92749, 4.933788, 4.939488, 
    4.944591, 4.949139, 4.953203, 4.956876, 4.960257, 4.963455, 4.966567, 
    4.969674, 4.973719, 4.973058, 4.975548, 4.978137, 4.98067, 4.983167, 
    4.986171, 4.988875, 4.991373, 4.994223, 4.997348, 5.000774, 5.004288, 
    5.007689, 5.009979, 5.010575, 5.010211, 5.008013, 5.003575, 4.996533, 
    4.986623, 4.973759, 4.958113, 4.940172, 4.920749, 4.900939, 4.881996, 
    4.865181, 4.851587, 4.842009, 4.83686, 4.836168, 4.83962, 4.846628, 
    4.856417,
  // totalHeight(20,36, 0-49)
    4.901495, 4.908389, 4.915284, 4.921958, 4.92825, 4.934066, 4.939364, 
    4.944149, 4.948456, 4.952359, 4.955939, 4.959299, 4.962548, 4.965801, 
    4.969179, 4.971826, 4.972733, 4.975375, 4.977877, 4.980225, 4.982509, 
    4.985884, 4.988856, 4.991599, 4.994495, 4.99746, 5.00048, 5.003342, 
    5.005812, 5.007051, 5.006406, 5.005326, 5.002304, 4.996975, 4.989042, 
    4.97832, 4.964816, 4.948807, 4.930867, 4.911874, 4.892938, 4.87528, 
    4.860076, 4.848299, 4.84061, 4.837299, 4.838289, 4.843188, 4.85136, 
    4.861993,
  // totalHeight(20,37, 0-49)
    4.905167, 4.911334, 4.917521, 4.923526, 4.929215, 4.934506, 4.939363, 
    4.943795, 4.947833, 4.95154, 4.954994, 4.958288, 4.961529, 4.964836, 
    4.968349, 4.969948, 4.972336, 4.975077, 4.977478, 4.979656, 4.981754, 
    4.985441, 4.988646, 4.991607, 4.994504, 4.99724, 4.999755, 5.001844, 
    5.003247, 5.003323, 5.001387, 4.999458, 4.995503, 4.989217, 4.980371, 
    4.968874, 4.954834, 4.938624, 4.9209, 4.902584, 4.884777, 4.868644, 
    4.855253, 4.845448, 4.839749, 4.838326, 4.841006, 4.847328, 4.856611, 
    4.868018,
  // totalHeight(20,38, 0-49)
    4.909193, 4.914583, 4.920015, 4.925317, 4.930371, 4.935106, 4.939497, 
    4.943548, 4.947289, 4.950776, 4.954073, 4.957259, 4.960435, 4.96371, 
    4.967225, 4.968122, 4.971893, 4.974655, 4.976923, 4.97893, 4.980852, 
    4.984771, 4.988155, 4.991285, 4.994119, 4.996551, 4.998464, 4.999669, 
    4.999884, 4.99871, 4.995449, 4.992558, 4.987595, 4.98032, 4.970589, 
    4.958406, 4.943982, 4.927779, 4.910518, 4.893145, 4.876726, 4.862342, 
    4.85094, 4.84322, 4.839568, 4.840035, 4.844362, 4.852028, 4.862319, 
    4.874377,
  // totalHeight(20,39, 0-49)
    4.913477, 4.918053, 4.922704, 4.927279, 4.931678, 4.93584, 4.939745, 
    4.943396, 4.946823, 4.950062, 4.953173, 4.956218, 4.959277, 4.962446, 
    4.965847, 4.966341, 4.971383, 4.974071, 4.976166, 4.977993, 4.979737, 
    4.983795, 4.987283, 4.990516, 4.993211, 4.995252, 4.99647, 4.996691, 
    4.995628, 4.99314, 4.988544, 4.984612, 4.978605, 4.970356, 4.959818, 
    4.94709, 4.932482, 4.916533, 4.900011, 4.883851, 4.869068, 4.856631, 
    4.847351, 4.841784, 4.840184, 4.842492, 4.848373, 4.857256, 4.868401, 
    4.880943,
  // totalHeight(20,40, 0-49)
    4.917906, 4.921646, 4.925501, 4.929339, 4.933074, 4.936653, 4.940061, 
    4.9433, 4.946392, 4.949367, 4.952266, 4.955137, 4.958039, 4.961041, 
    4.964238, 4.964564, 4.970736, 4.97326, 4.975143, 4.976772, 4.978323, 
    4.982419, 4.985922, 4.989172, 4.991644, 4.993212, 4.993649, 4.99281, 
    4.990404, 4.98657, 4.980658, 4.975645, 4.968606, 4.959457, 4.948241, 
    4.93516, 4.920611, 4.905192, 4.889691, 4.87501, 4.86208, 4.851747, 
    4.844676, 4.84128, 4.841683, 4.845729, 4.853019, 4.862945, 4.874746, 
    4.887564,
  // totalHeight(20,41, 0-49)
    4.922345, 4.925241, 4.928298, 4.9314, 4.934471, 4.937466, 4.940372, 
    4.943191, 4.945935, 4.948627, 4.951293, 4.953965, 4.956676, 4.95947, 
    4.9624, 4.962718, 4.969854, 4.972135, 4.973769, 4.975179, 4.976512, 
    4.980538, 4.983962, 4.987133, 4.989291, 4.9903, 4.98989, 4.987938, 
    4.984165, 4.978992, 4.971818, 4.965739, 4.957735, 4.94781, 4.936104, 
    4.92291, 4.908694, 4.894094, 4.879889, 4.866925, 4.856025, 4.847902, 
    4.84307, 4.841802, 4.844105, 4.849738, 4.858246, 4.868992, 4.881212, 
    4.894058,
  // totalHeight(20,42, 0-49)
    4.926642, 4.928699, 4.930964, 4.93334, 4.935758, 4.938178, 4.940584, 
    4.942979, 4.945368, 4.947763, 4.950179, 4.95263, 4.955127, 4.957681, 
    4.960309, 4.96071, 4.96862, 4.970598, 4.971952, 4.973114, 4.974197, 
    4.978046, 4.981288, 4.98428, 4.986035, 4.986415, 4.985108, 4.982025, 
    4.976905, 4.970449, 4.962109, 4.955034, 4.946192, 4.935675, 4.923714, 
    4.910677, 4.897085, 4.88359, 4.870934, 4.859879, 4.851132, 4.845262, 
    4.842635, 4.843394, 4.847439, 4.854456, 4.863945, 4.875252, 4.887619, 
    4.900222,
  // totalHeight(20,43, 0-49)
    4.930626, 4.931849, 4.933344, 4.935014, 4.936798, 4.938658, 4.940579, 
    4.942554, 4.944587, 4.94668, 4.948834, 4.951047, 4.953313, 4.955612, 
    4.957922, 4.958442, 4.966921, 4.968552, 4.9696, 4.970482, 4.971275, 
    4.974844, 4.977806, 4.980515, 4.981785, 4.981482, 4.979256, 4.975064, 
    4.968668, 4.961029, 4.951668, 4.943729, 4.934234, 4.923361, 4.911418, 
    4.898832, 4.886153, 4.874021, 4.86312, 4.854114, 4.847578, 4.843935, 
    4.843416, 4.846041, 4.851618, 4.85977, 4.869962, 4.881538, 4.893755, 
    4.905829,
  // totalHeight(20,44, 0-49)
    4.93411, 4.934515, 4.935261, 4.936253, 4.937433, 4.938762, 4.940217, 
    4.941791, 4.943477, 4.94527, 4.94716, 4.949131, 4.951157, 4.953195, 
    4.955183, 4.955816, 4.964656, 4.965913, 4.966628, 4.967195, 4.967651, 
    4.970848, 4.973435, 4.975765, 4.976482, 4.975461, 4.972332, 4.967094, 
    4.959548, 4.950883, 4.940692, 4.93208, 4.922171, 4.911213, 4.89958, 
    4.887739, 4.876243, 4.865695, 4.856701, 4.849814, 4.845474, 4.843967, 
    4.845396, 4.84967, 4.856519, 4.865516, 4.876104, 4.887634, 4.899394, 
    4.910653,
  // totalHeight(20,45, 0-49)
    4.936903, 4.936502, 4.936521, 4.936871, 4.937485, 4.938321, 4.939349, 
    4.940551, 4.941915, 4.943424, 4.945058, 4.946791, 4.948578, 4.950358, 
    4.952039, 4.952745, 4.961742, 4.962612, 4.962971, 4.963184, 4.963254, 
    4.965993, 4.968124, 4.96999, 4.970107, 4.968362, 4.964381, 4.958209, 
    4.949688, 4.940206, 4.929422, 4.920379, 4.910328, 4.899585, 4.888559, 
    4.877738, 4.867655, 4.858856, 4.851855, 4.847086, 4.844861, 4.845332, 
    4.848487, 4.854145, 4.861969, 4.87149, 4.882148, 4.893308, 4.904304, 
    4.914479,
  // totalHeight(20,46, 0-49)
    4.938819, 4.937624, 4.936943, 4.936685, 4.936779, 4.93717, 4.937817, 
    4.938693, 4.939772, 4.94103, 4.942434, 4.943947, 4.945509, 4.947042, 
    4.948433, 4.949158, 4.958127, 4.958603, 4.958583, 4.958401, 4.958039, 
    4.960252, 4.961856, 4.963193, 4.962687, 4.960245, 4.955501, 4.948549, 
    4.939279, 4.929226, 4.918125, 4.908927, 4.899035, 4.888804, 4.878668, 
    4.869109, 4.860616, 4.853668, 4.848677, 4.845958, 4.845698, 4.847935, 
    4.852553, 4.859291, 4.86776, 4.877473, 4.887864, 4.898334, 4.908283, 
    4.91715,
  // totalHeight(20,47, 0-49)
    4.93972, 4.937729, 4.936366, 4.935534, 4.935153, 4.935151, 4.935477, 
    4.936083, 4.936932, 4.937986, 4.939202, 4.940526, 4.941891, 4.9432, 
    4.944324, 4.945001, 4.953781, 4.953864, 4.95344, 4.952825, 4.951988, 
    4.953621, 4.954652, 4.955418, 4.954295, 4.951216, 4.945836, 4.938297, 
    4.928536, 4.918194, 4.907071, 4.898016, 4.888585, 4.879151, 4.870152, 
    4.862043, 4.85526, 4.850199, 4.847168, 4.84637, 4.847877, 4.851622, 
    4.857403, 4.864896, 4.873673, 4.883236, 4.893039, 4.902533, 4.911198, 
    4.918588,
  // totalHeight(20,48, 0-49)
    4.939519, 4.93672, 4.934682, 4.933303, 4.932487, 4.932148, 4.932213, 
    4.932616, 4.933301, 4.934213, 4.935294, 4.936477, 4.937681, 4.938794, 
    4.939677, 4.940239, 4.948703, 4.94839, 4.94754, 4.946457, 4.945107, 
    4.946132, 4.946567, 4.946746, 4.945043, 4.94142, 4.935561, 4.927656, 
    4.917686, 4.907351, 4.896503, 4.88789, 4.879201, 4.870818, 4.863158, 
    4.856635, 4.85162, 4.848419, 4.847244, 4.848188, 4.851223, 4.856192, 
    4.862821, 4.870739, 4.879495, 4.888591, 4.89752, 4.905799, 4.913006, 
    4.918834,
  // totalHeight(20,49, 0-49)
    4.940613, 4.936409, 4.933164, 4.930776, 4.929138, 4.928135, 4.927667, 
    4.927631, 4.927937, 4.928491, 4.9292, 4.92996, 4.930647, 4.931097, 
    4.931102, 4.930818, 4.946164, 4.943949, 4.940964, 4.937904, 4.934816, 
    4.936986, 4.938692, 4.94071, 4.939893, 4.93633, 4.929495, 4.919771, 
    4.907046, 4.894641, 4.882136, 4.8747, 4.867539, 4.861034, 4.855579, 
    4.851521, 4.849131, 4.84859, 4.849968, 4.853214, 4.858169, 4.864559, 
    4.872037, 4.88018, 4.888537, 4.896647, 4.90409, 4.910515, 4.915682, 
    4.919499,
  // totalHeight(21,0, 0-49)
    4.867756, 4.87136, 4.876185, 4.881904, 4.888227, 4.894917, 4.901782, 
    4.908686, 4.915534, 4.922264, 4.928842, 4.935246, 4.941461, 4.947464, 
    4.953222, 4.958513, 4.964422, 4.96916, 4.973463, 4.977247, 4.98037, 
    4.982961, 4.984521, 4.984962, 4.984047, 4.981614, 4.977492, 4.971577, 
    4.963781, 4.95417, 4.942726, 4.929893, 4.915575, 4.900093, 4.883879, 
    4.867457, 4.851445, 4.836494, 4.823259, 4.812335, 4.804196, 4.799148, 
    4.797297, 4.798529, 4.802532, 4.808812, 4.816741, 4.82561, 4.834689, 
    4.843285,
  // totalHeight(21,1, 0-49)
    4.869227, 4.873135, 4.878213, 4.88414, 4.890633, 4.897455, 4.904428, 
    4.911416, 4.918332, 4.925114, 4.931731, 4.938162, 4.944387, 4.950385, 
    4.956112, 4.961147, 4.967659, 4.972268, 4.976444, 4.980152, 4.983257, 
    4.986171, 4.988067, 4.988924, 4.988447, 4.98646, 4.982759, 4.977232, 
    4.969764, 4.960455, 4.949201, 4.93672, 4.922586, 4.907089, 4.890637, 
    4.87375, 4.857055, 4.841236, 4.827, 4.815002, 4.805791, 4.799745, 
    4.797029, 4.797587, 4.801143, 4.807224, 4.815208, 4.824379, 4.833981, 
    4.843285,
  // totalHeight(21,2, 0-49)
    4.87042, 4.874584, 4.879874, 4.885972, 4.892601, 4.899534, 4.906593, 
    4.913648, 4.920613, 4.927431, 4.934066, 4.940497, 4.946706, 4.952666, 
    4.958333, 4.963048, 4.970029, 4.974471, 4.978471, 4.982044, 4.985077, 
    4.988253, 4.990441, 4.991687, 4.991656, 4.99017, 4.987002, 4.982033, 
    4.97512, 4.966384, 4.955632, 4.943846, 4.930265, 4.915128, 4.898799, 
    4.881767, 4.864641, 4.848114, 4.832927, 4.819794, 4.809337, 4.802019, 
    4.798089, 4.79757, 4.800246, 4.805697, 4.813336, 4.822461, 4.832316, 
    4.842153,
  // totalHeight(21,3, 0-49)
    4.871417, 4.875794, 4.881257, 4.88749, 4.894225, 4.90124, 4.90836, 
    4.91546, 4.922452, 4.92928, 4.935906, 4.942309, 4.948469, 4.954359, 
    4.959938, 4.964278, 4.971559, 4.975809, 4.979591, 4.982981, 4.985889, 
    4.989264, 4.991691, 4.993279, 4.993685, 4.992729, 4.990175, 4.985899, 
    4.979735, 4.971802, 4.96182, 4.951028, 4.938334, 4.923909, 4.908056, 
    4.891205, 4.873922, 4.856891, 4.840857, 4.826586, 4.81477, 4.805964, 
    4.800524, 4.798568, 4.799973, 4.804396, 4.811304, 4.820037, 4.829866, 
    4.840038,
  // totalHeight(21,4, 0-49)
    4.872332, 4.876885, 4.882481, 4.888814, 4.895623, 4.902688, 4.909839, 
    4.916954, 4.923941, 4.930746, 4.937329, 4.943668, 4.949744, 4.955535, 
    4.961005, 4.964917, 4.972301, 4.976346, 4.979885, 4.983051, 4.985792, 
    4.989301, 4.991906, 4.993781, 4.994592, 4.994171, 4.992283, 4.9888, 
    4.983535, 4.976586, 4.967588, 4.958031, 4.946498, 4.933095, 4.91804, 
    4.90169, 4.884544, 4.867239, 4.850518, 4.835167, 4.821952, 4.811521, 
    4.804342, 4.800659, 4.800459, 4.8035, 4.809333, 4.817359, 4.826887, 
    4.837183,
  // totalHeight(21,5, 0-49)
    4.873298, 4.87799, 4.883683, 4.890078, 4.896924, 4.904002, 4.91115, 
    4.91824, 4.925184, 4.931925, 4.938425, 4.94466, 4.950615, 4.956275, 
    4.961616, 4.965065, 4.972339, 4.976171, 4.979454, 4.982371, 4.984913, 
    4.988491, 4.99121, 4.993308, 4.994482, 4.994578, 4.993377, 4.990749, 
    4.986489, 4.980652, 4.972798, 4.964639, 4.954481, 4.942347, 4.928371, 
    4.912815, 4.896089, 4.878769, 4.861557, 4.845256, 4.830675, 4.818562, 
    4.809506, 4.803884, 4.801821, 4.803196, 4.807662, 4.8147, 4.823673, 
    4.833878,
  // totalHeight(21,6, 0-49)
    4.874443, 4.879241, 4.884993, 4.891414, 4.898254, 4.905306, 4.912405, 
    4.919427, 4.926284, 4.932917, 4.939289, 4.945377, 4.951174, 4.956671, 
    4.961865, 4.964837, 4.971784, 4.975398, 4.97842, 4.981078, 4.983403, 
    4.986985, 4.989758, 4.992006, 4.993488, 4.994068, 4.99355, 4.991801, 
    4.988611, 4.983963, 4.977353, 4.970687, 4.962039, 4.951355, 4.938675, 
    4.924161, 4.908125, 4.891047, 4.87358, 4.856506, 4.840674, 4.826908, 
    4.815924, 4.808243, 4.804142, 4.803638, 4.806506, 4.812325, 4.820523, 
    4.830435,
  // totalHeight(21,7, 0-49)
    4.87588, 4.880752, 4.88653, 4.892937, 4.899731, 4.90671, 4.913714, 
    4.920619, 4.927339, 4.933815, 4.940012, 4.945911, 4.951509, 4.956812, 
    4.961838, 4.964347, 4.970757, 4.97415, 4.976916, 4.979318, 4.981421, 
    4.98495, 4.987716, 4.990044, 4.991772, 4.992788, 4.992926, 4.992055, 
    4.989957, 4.986527, 4.981206, 4.976059, 4.968983, 4.959855, 4.948626, 
    4.93535, 4.92023, 4.903647, 4.886172, 4.868548, 4.851635, 4.836328, 
    4.823456, 4.813686, 4.807459, 4.804945, 4.806056, 4.810474, 4.81771, 
    4.82715,
  // totalHeight(21,8, 0-49)
    4.8777, 4.882618, 4.888388, 4.894741, 4.901444, 4.908303, 4.915162, 
    4.9219, 4.928433, 4.934703, 4.940678, 4.946343, 4.951704, 4.95678, 
    4.961609, 4.963711, 4.969393, 4.972557, 4.975082, 4.977241, 4.979133, 
    4.982553, 4.985257, 4.987593, 4.989506, 4.990901, 4.99165, 4.991627, 
    4.990613, 4.988391, 4.984363, 4.980696, 4.975188, 4.967651, 4.957954, 
    4.946052, 4.932031, 4.916164, 4.898924, 4.880996, 4.863228, 4.846558, 
    4.831919, 4.82012, 4.811763, 4.807185, 4.806442, 4.80934, 4.81547, 
    4.824277,
  // totalHeight(21,9, 0-49)
    4.879959, 4.884899, 4.890628, 4.89689, 4.903462, 4.910154, 4.916817, 
    4.923337, 4.929632, 4.935648, 4.941355, 4.946746, 4.951833, 4.956645, 
    4.961241, 4.963027, 4.967825, 4.970748, 4.97305, 4.974993, 4.976692, 
    4.979956, 4.982547, 4.98483, 4.986863, 4.988575, 4.989882, 4.990657, 
    4.99069, 4.989635, 4.986869, 4.984592, 4.98059, 4.974617, 4.966471, 
    4.956012, 4.943221, 4.928251, 4.911475, 4.893493, 4.87512, 4.857318, 
    4.8411, 4.827405, 4.816993, 4.810369, 4.807745, 4.80905, 4.813972, 
    4.822018,
  // totalHeight(21,10, 0-49)
    4.882683, 4.887622, 4.893283, 4.899419, 4.905817, 4.912298, 4.918719, 
    4.924973, 4.930984, 4.936702, 4.942099, 4.947176, 4.951952, 4.956465, 
    4.960778, 4.962388, 4.966177, 4.968843, 4.970945, 4.972705, 4.974249, 
    4.977313, 4.979748, 4.98192, 4.984013, 4.985978, 4.98778, 4.989291, 
    4.99031, 4.990362, 4.988803, 4.987789, 4.985182, 4.980694, 4.97406, 
    4.965057, 4.953567, 4.939633, 4.923513, 4.905717, 4.887003, 4.868331, 
    4.85077, 4.835371, 4.823044, 4.814457, 4.809978, 4.809673, 4.813326, 
    4.820508,
  // totalHeight(21,11, 0-49)
    4.885859, 4.890782, 4.896351, 4.902331, 4.90852, 4.914749, 4.920887, 
    4.926834, 4.932517, 4.937896, 4.942946, 4.947676, 4.952104, 4.956275, 
    4.960248, 4.961854, 4.964558, 4.966954, 4.968882, 4.970501, 4.971934, 
    4.974759, 4.977002, 4.979015, 4.981116, 4.983275, 4.985504, 4.987677, 
    4.989609, 4.990688, 4.990268, 4.990361, 4.989007, 4.985883, 4.980674, 
    4.973091, 4.962924, 4.950112, 4.934801, 4.917403, 4.898602, 4.879333, 
    4.860695, 4.843828, 4.829777, 4.819361, 4.813109, 4.811215, 4.813574, 
    4.819819,
  // totalHeight(21,12, 0-49)
    4.88944, 4.894337, 4.899799, 4.905598, 4.911548, 4.917494, 4.923313, 
    4.928915, 4.934238, 4.939242, 4.943916, 4.948267, 4.952316, 4.956103, 
    4.959673, 4.961469, 4.963051, 4.965169, 4.966954, 4.968485, 4.96986, 
    4.972414, 4.974438, 4.976257, 4.978319, 4.980617, 4.983204, 4.985958, 
    4.988717, 4.990734, 4.99138, 4.99241, 4.992143, 4.990234, 4.986331, 
    4.980086, 4.971216, 4.959564, 4.945173, 4.928348, 4.909691, 4.890091, 
    4.870652, 4.852578, 4.837027, 4.824958, 4.81705, 4.813632, 4.814701, 
    4.819964,
  // totalHeight(21,13, 0-49)
    4.893345, 4.898217, 4.90356, 4.909164, 4.914856, 4.920492, 4.925966, 
    4.931196, 4.936131, 4.94074, 4.945012, 4.948959, 4.952602, 4.955966, 
    4.959073, 4.961245, 4.961709, 4.963559, 4.96524, 4.96674, 4.96812, 
    4.970376, 4.972166, 4.973768, 4.975757, 4.978142, 4.981021, 4.984272, 
    4.987758, 4.990619, 4.99226, 4.994047, 4.99469, 4.993832, 4.991089, 
    4.98607, 4.978432, 4.967936, 4.954527, 4.93841, 4.920095, 4.900408, 
    4.880437, 4.861424, 4.844614, 4.831095, 4.821679, 4.816827, 4.816639, 
    4.820898,
  // totalHeight(21,14, 0-49)
    4.897468, 4.902321, 4.907547, 4.912951, 4.918373, 4.923688, 4.928799, 
    4.93364, 4.93817, 4.942365, 4.946223, 4.949754, 4.95297, 4.95588, 
    4.958479, 4.961169, 4.960548, 4.962161, 4.963795, 4.965333, 4.966787, 
    4.968728, 4.97028, 4.971656, 4.973548, 4.975982, 4.979085, 4.982744, 
    4.986854, 4.990458, 4.993018, 4.995389, 4.996763, 4.99678, 4.995036, 
    4.991111, 4.98461, 4.975227, 4.962822, 4.947505, 4.929689, 4.910128, 
    4.889874, 4.870183, 4.852361, 4.837605, 4.826849, 4.820671, 4.819281, 
    4.822535,
  // totalHeight(21,15, 0-49)
    4.901683, 4.906533, 4.911652, 4.916859, 4.922011, 4.927, 4.931743, 
    4.936191, 4.94031, 4.944088, 4.94753, 4.950641, 4.953424, 4.955871, 
    4.957943, 4.96121, 4.959546, 4.960984, 4.962644, 4.9643, 4.965909, 
    4.967529, 4.968853, 4.970014, 4.971802, 4.974249, 4.977513, 4.981489, 
    4.986113, 4.990354, 4.993762, 4.996544, 4.998473, 4.999189, 4.998278, 
    4.995298, 4.989818, 4.981478, 4.970063, 4.955593, 4.938392, 4.919131, 
    4.898813, 4.878683, 4.860091, 4.844313, 4.832389, 4.825014, 4.822492, 
    4.824755,
  // totalHeight(21,16, 0-49)
    4.905852, 4.910719, 4.915746, 4.92077, 4.925663, 4.930331, 4.934713, 
    4.938773, 4.942492, 4.945868, 4.948905, 4.951612, 4.953979, 4.955981, 
    4.95755, 4.961321, 4.958642, 4.960001, 4.961782, 4.963653, 4.965511, 
    4.966817, 4.967943, 4.968918, 4.970611, 4.973051, 4.976418, 4.980618, 
    4.985636, 4.9904, 4.994579, 4.99761, 4.999923, 5.001165, 5.00092, 
    4.99873, 4.994142, 4.986749, 4.976277, 4.962667, 4.946156, 4.927331, 
    4.907132, 4.886779, 4.86764, 4.851046, 4.838132, 4.82969, 4.826118, 
    4.82742,
  // totalHeight(21,17, 0-49)
    4.909837, 4.914738, 4.919692, 4.924548, 4.929195, 4.93356, 4.9376, 
    4.941293, 4.944641, 4.947648, 4.950324, 4.95267, 4.954671, 4.956281, 
    4.957415, 4.961463, 4.957752, 4.959157, 4.961174, 4.963372, 4.965584, 
    4.966605, 4.967587, 4.968428, 4.970053, 4.97248, 4.975895, 4.980227, 
    4.985517, 4.99068, 4.995541, 4.998661, 5.001194, 5.002797, 5.003052, 
    5.001498, 4.997662, 4.991107, 4.98151, 4.968741, 4.95296, 4.934667, 
    4.914736, 4.894343, 4.874856, 4.857644, 4.843911, 4.834536, 4.83, 4.830382,
  // totalHeight(21,18, 0-49)
    4.913497, 4.918441, 4.923331, 4.928032, 4.932451, 4.936535, 4.940263, 
    4.943635, 4.946665, 4.949371, 4.951762, 4.953833, 4.955557, 4.956873, 
    4.957686, 4.961622, 4.956789, 4.958377, 4.96076, 4.963412, 4.9661, 
    4.966885, 4.967799, 4.968584, 4.970194, 4.972615, 4.97604, 4.980412, 
    4.985839, 4.991264, 4.996696, 4.999753, 5.002348, 5.004149, 5.004743, 
    5.003669, 5.000443, 4.994608, 4.985798, 4.973829, 4.958785, 4.94109, 
    4.921543, 4.901266, 4.881607, 4.863956, 4.849568, 4.839391, 4.833985, 
    4.833497,
  // totalHeight(21,19, 0-49)
    4.9167, 4.921665, 4.926477, 4.931019, 4.93522, 4.939054, 4.942522, 
    4.945646, 4.948455, 4.950972, 4.953205, 4.955136, 4.956722, 4.957885, 
    4.958528, 4.961836, 4.95568, 4.957586, 4.960464, 4.963702, 4.967002, 
    4.967633, 4.968585, 4.96942, 4.971097, 4.973547, 4.976954, 4.981276, 
    4.986701, 4.992226, 4.998084, 5.00092, 5.003414, 5.00525, 5.006023, 
    5.005275, 5.00252, 4.997281, 4.989166, 4.977938, 4.963619, 4.94656, 
    4.927482, 4.90745, 4.887774, 4.869849, 4.854956, 4.84411, 4.837931, 
    4.836633,
  // totalHeight(21,20, 0-49)
    4.920373, 4.926408, 4.932198, 4.937615, 4.942574, 4.947017, 4.95092, 
    4.954266, 4.957061, 4.959322, 4.961086, 4.962402, 4.963344, 4.963996, 
    4.96446, 30, 4.958336, 4.959911, 4.962055, 4.964373, 4.966731, 4.965669, 
    4.965298, 4.965133, 4.966242, 4.968559, 4.972223, 4.977122, 4.983384, 
    4.989923, 4.997092, 5.000469, 5.003476, 5.005798, 5.007044, 5.006776, 
    5.004527, 4.999839, 4.992319, 4.981717, 4.96802, 4.951524, 4.932887, 
    4.913119, 4.893489, 4.875374, 4.860076, 4.848648, 4.841766, 4.839701,
  // totalHeight(21,21, 0-49)
    4.922716, 4.928973, 4.934875, 4.9403, 4.945176, 4.949471, 4.95318, 
    4.956317, 4.958914, 4.96101, 4.962654, 4.963908, 4.964848, 4.965567, 
    4.966182, 30, 4.955145, 4.957202, 4.959885, 4.962759, 4.965636, 4.964164, 
    4.963536, 4.963161, 4.964198, 4.966575, 4.970424, 4.975614, 4.982278, 
    4.989311, 4.997245, 5.000715, 5.003937, 5.006592, 5.008276, 5.008539, 
    5.006902, 5.002893, 4.996096, 4.986228, 4.97323, 4.957343, 4.939162, 
    4.919639, 4.900001, 4.881614, 4.865797, 4.85364, 4.845881, 4.842846,
  // totalHeight(21,22, 0-49)
    4.924577, 4.931123, 4.937216, 4.942735, 4.947618, 4.951845, 4.955435, 
    4.958422, 4.960857, 4.962803, 4.964324, 4.965492, 4.966395, 4.967139, 
    4.967857, 30, 4.952854, 4.955309, 4.958461, 4.96184, 4.965202, 4.963355, 
    4.962503, 4.961944, 4.962914, 4.96533, 4.96931, 4.974701, 4.981636, 
    4.988995, 4.997468, 5.000855, 5.004099, 5.006884, 5.008801, 5.009401, 
    5.008202, 5.004722, 4.998529, 4.989316, 4.976982, 4.961714, 4.944051, 
    4.92488, 4.905382, 4.886895, 4.870741, 4.858034, 4.849556, 4.845685,
  // totalHeight(21,23, 0-49)
    4.925975, 4.932854, 4.939191, 4.944864, 4.949818, 4.954044, 4.957575, 
    4.960462, 4.962778, 4.964598, 4.966004, 4.967083, 4.967932, 4.968668, 
    4.969452, 30, 4.951511, 4.954235, 4.957705, 4.961428, 4.965119, 4.962908, 
    4.961822, 4.961064, 4.961936, 4.964339, 4.968385, 4.973899, 4.98101, 
    4.988581, 4.997424, 5.000678, 5.003872, 5.006702, 5.008762, 5.009603, 
    5.008744, 5.0057, 5.000029, 4.9914, 4.97968, 4.96501, 4.947873, 4.929098, 
    4.909818, 4.891339, 4.874972, 4.861847, 4.852779, 4.848183,
  // totalHeight(21,24, 0-49)
    4.926955, 4.934186, 4.940796, 4.946662, 4.951729, 4.956, 4.959518, 
    4.962349, 4.964579, 4.966302, 4.96761, 4.968601, 4.969385, 4.970094, 
    4.970906, 30, 4.951337, 4.954191, 4.957818, 4.961719, 4.965586, 4.963124, 
    4.961879, 4.96099, 4.961792, 4.964177, 4.968248, 4.973822, 4.981027, 
    4.988714, 4.997774, 5.000921, 5.004061, 5.006891, 5.009009, 5.009973, 
    5.009304, 5.006517, 5.001168, 4.992916, 4.981607, 4.967354, 4.950599, 
    4.932136, 4.913054, 4.894632, 4.878164, 4.864782, 4.855316, 4.850201,
  // totalHeight(21,25, 0-49)
    4.927581, 4.93516, 4.94205, 4.948121, 4.953326, 4.957671, 4.961206, 
    4.964014, 4.96619, 4.967835, 4.969058, 4.969966, 4.970678, 4.971337, 
    4.972132, 30, 4.951993, 4.954841, 4.958466, 4.962369, 4.966248, 4.963695, 
    4.962402, 4.961487, 4.962284, 4.964675, 4.968763, 4.974359, 4.981592, 
    4.989312, 4.998431, 5.001542, 5.004662, 5.007491, 5.009628, 5.010636, 
    5.010038, 5.007354, 5.002141, 4.994059, 4.982945, 4.968903, 4.952358, 
    4.934081, 4.915137, 4.896785, 4.880301, 4.866809, 4.857136, 4.851721,
  // totalHeight(21,26, 0-49)
    4.927925, 4.935825, 4.942978, 4.949254, 4.954605, 4.959037, 4.962613, 
    4.965418, 4.967557, 4.969142, 4.970285, 4.971105, 4.971728, 4.972306, 
    4.973034, 30, 4.953425, 4.95613, 4.959591, 4.963326, 4.96705, 4.964577, 
    4.963362, 4.962536, 4.963402, 4.965837, 4.969944, 4.975535, 4.982742, 
    4.990416, 4.999442, 5.002605, 5.005761, 5.008602, 5.010732, 5.011711, 
    5.011069, 5.008329, 5.003057, 4.994917, 4.983764, 4.969701, 4.953165, 
    4.934923, 4.91604, 4.89776, 4.881342, 4.867894, 4.858222, 4.852753,
  // totalHeight(21,27, 0-49)
    4.92806, 4.936237, 4.943624, 4.950087, 4.955577, 4.960105, 4.963733, 
    4.96655, 4.968665, 4.970191, 4.971249, 4.971961, 4.972464, 4.972912, 
    4.973501, 30, 4.955719, 4.958138, 4.961273, 4.964661, 4.968061, 4.965804, 
    4.964757, 4.964105, 4.965088, 4.967585, 4.971696, 4.977244, 4.98436, 
    4.99191, 5.000689, 5.003982, 5.007212, 5.01007, 5.012156, 5.013031, 
    5.01223, 5.009284, 5.00377, 4.995371, 4.983961, 4.969677, 4.952976, 
    4.93465, 4.915774, 4.897588, 4.881337, 4.868097, 4.85864, 4.853362,
  // totalHeight(21,28, 0-49)
    4.928054, 4.936454, 4.944035, 4.950661, 4.956285, 4.960913, 4.964603, 
    4.967442, 4.969531, 4.970989, 4.971935, 4.972499, 4.972823, 4.973068, 
    4.973427, 30, 4.959241, 4.961226, 4.963868, 4.966732, 4.969642, 4.967668, 
    4.96682, 4.966366, 4.967466, 4.969997, 4.974066, 4.979512, 4.986459, 
    4.993795, 5.002191, 5.005653, 5.008963, 5.011804, 5.013775, 5.014439, 
    5.013337, 5.010012, 5.004061, 4.995199, 4.983335, 4.968651, 4.951647, 
    4.933157, 4.914279, 4.896254, 4.880302, 4.867464, 4.858457, 4.853627,
  // totalHeight(21,29, 0-49)
    4.92797, 4.936532, 4.944271, 4.951048, 4.956806, 4.961545, 4.965309, 
    4.968172, 4.970227, 4.971584, 4.972364, 4.972703, 4.972755, 4.972694, 
    4.972711, 30, 4.963769, 4.965175, 4.967158, 4.969325, 4.971568, 4.96982, 
    4.969094, 4.968768, 4.969911, 4.972406, 4.976363, 4.981632, 4.988328, 
    4.995357, 5.003223, 5.006826, 5.010169, 5.01293, 5.014711, 5.015079, 
    5.013591, 5.0098, 5.003335, 4.99394, 4.981572, 4.966462, 4.949168, 
    4.930563, 4.911772, 4.894035, 4.878546, 4.866288, 4.85792, 4.853728,
  // totalHeight(21,30, 0-49)
    4.926956, 4.934618, 4.941468, 4.947391, 4.952364, 4.956439, 4.959708, 
    4.962296, 4.964333, 4.965935, 4.967184, 4.968123, 4.968738, 4.968968, 
    4.968709, 4.975595, 4.962874, 4.964472, 4.967275, 4.970613, 4.974156, 
    4.97453, 4.975579, 4.976661, 4.978667, 4.98145, 4.985137, 4.989669, 
    4.995262, 5.000958, 5.007199, 5.009936, 5.012409, 5.014312, 5.015257, 
    5.014821, 5.012557, 5.008026, 5.000863, 4.990838, 4.977942, 4.962452, 
    4.944969, 4.926406, 4.9079, 4.890683, 4.875904, 4.864484, 4.857009, 
    4.853695,
  // totalHeight(21,31, 0-49)
    4.926929, 4.934672, 4.941601, 4.947601, 4.95264, 4.956754, 4.960025, 
    4.962573, 4.964523, 4.965997, 4.967094, 4.96788, 4.968374, 4.968542, 
    4.968293, 4.975252, 4.964764, 4.96593, 4.968161, 4.970851, 4.97374, 
    4.974269, 4.975286, 4.976324, 4.978278, 4.981052, 4.98479, 4.98941, 
    4.995051, 5.0007, 5.006574, 5.009628, 5.012319, 5.014328, 5.015259, 
    5.014685, 5.012158, 5.007254, 4.999632, 4.989102, 4.975713, 4.959807, 
    4.942053, 4.923415, 4.905064, 4.888221, 4.874006, 4.863276, 4.856546, 
    4.853962,
  // totalHeight(21,32, 0-49)
    4.926838, 4.934477, 4.941327, 4.947276, 4.952287, 4.956389, 4.959658, 
    4.962198, 4.964133, 4.965584, 4.966657, 4.967435, 4.967957, 4.968214, 
    4.968139, 4.974419, 4.966065, 4.966943, 4.968725, 4.970888, 4.973237, 
    4.974019, 4.975111, 4.976216, 4.978195, 4.980991, 4.984751, 4.989377, 
    4.994931, 5.000389, 5.005764, 5.009021, 5.011818, 5.013818, 5.014621, 
    5.013795, 5.0109, 5.005525, 4.997361, 4.986272, 4.972367, 4.956063, 
    4.938097, 4.919488, 4.901426, 4.885119, 4.871639, 4.861775, 4.855964, 
    4.854273,
  // totalHeight(21,33, 0-49)
    4.926754, 4.934147, 4.940796, 4.946594, 4.951506, 4.955551, 4.958797, 
    4.961343, 4.963299, 4.964785, 4.96591, 4.966764, 4.967407, 4.967854, 
    4.968068, 4.973201, 4.966861, 4.967598, 4.969047, 4.970792, 4.972705, 
    4.973806, 4.97506, 4.976316, 4.978374, 4.981203, 4.984944, 4.989483, 
    4.994825, 4.999962, 5.004738, 5.008092, 5.010881, 5.012757, 5.013318, 
    5.012129, 5.00876, 5.002823, 4.994051, 4.982362, 4.967942, 4.951282, 
    4.93319, 4.914731, 4.897108, 4.881502, 4.868926, 4.86009, 4.855348, 
    4.854691,
  // totalHeight(21,34, 0-49)
    4.926736, 4.933774, 4.940129, 4.945702, 4.950455, 4.954404, 4.95761, 
    4.960158, 4.962151, 4.9637, 4.964916, 4.96589, 4.966699, 4.967385, 
    4.967942, 4.971733, 4.967276, 4.967985, 4.969195, 4.970612, 4.972173, 
    4.973621, 4.975093, 4.976563, 4.978733, 4.98159, 4.98526, 4.989622, 
    4.994627, 4.999331, 5.003438, 5.006778, 5.009446, 5.011085, 5.011292, 
    5.009635, 5.005699, 4.999127, 4.989699, 4.977401, 4.962496, 4.945557, 
    4.927455, 4.909292, 4.892269, 4.877531, 4.866017, 4.858353, 4.854806, 
    4.855289,
  // totalHeight(21,35, 0-49)
    4.926836, 4.933433, 4.939422, 4.944709, 4.949258, 4.953081, 4.956228, 
    4.95877, 4.960804, 4.96243, 4.96375, 4.964861, 4.965849, 4.966776, 
    4.967676, 4.970145, 4.967444, 4.968202, 4.969242, 4.970393, 4.971665, 
    4.973465, 4.975183, 4.976903, 4.979197, 4.982062, 4.985603, 4.989695, 
    4.994246, 4.998414, 5.001794, 5.005006, 5.007436, 5.008721, 5.008463, 
    5.00624, 5.001657, 4.994396, 4.984295, 4.971416, 4.9561, 4.938995, 
    4.921033, 4.903339, 4.887095, 4.873391, 4.863085, 4.856715, 4.854457, 
    4.856152,
  // totalHeight(21,36, 0-49)
    4.927101, 4.933189, 4.938755, 4.943709, 4.948019, 4.951687, 4.954755, 
    4.957284, 4.959356, 4.961058, 4.962487, 4.963735, 4.964891, 4.966037, 
    4.967238, 4.96855, 4.967488, 4.968328, 4.969235, 4.970166, 4.9712, 
    4.973329, 4.975299, 4.977283, 4.979695, 4.982537, 4.985882, 4.989611, 
    4.993591, 4.997127, 4.999732, 5.00269, 5.004757, 5.005571, 5.00474, 
    5.00186, 4.996566, 4.988592, 4.977838, 4.964443, 4.948833, 4.931724, 
    4.91409, 4.897061, 4.881786, 4.869282, 4.860319, 4.855337, 4.85443, 
    4.857368,
  // totalHeight(21,37, 0-49)
    4.927572, 4.933101, 4.938197, 4.942782, 4.946818, 4.950309, 4.95328, 
    4.955783, 4.957885, 4.959661, 4.961193, 4.962566, 4.963869, 4.965193, 
    4.966624, 4.967034, 4.967501, 4.96842, 4.969209, 4.969953, 4.970782, 
    4.9732, 4.975408, 4.97765, 4.980156, 4.982931, 4.986008, 4.989279, 
    4.992575, 4.995385, 4.997163, 4.999734, 5.00131, 5.001532, 5.000024, 
    4.996412, 4.990367, 4.981685, 4.970336, 4.956542, 4.940803, 4.923894, 
    4.906811, 4.890669, 4.876559, 4.865418, 4.857912, 4.854388, 4.854856, 
    4.859026,
  // totalHeight(21,38, 0-49)
    4.928286, 4.933214, 4.937806, 4.941989, 4.945725, 4.949013, 4.951869, 
    4.954332, 4.956453, 4.95829, 4.959915, 4.9614, 4.962823, 4.964279, 
    4.965862, 4.965644, 4.967535, 4.968503, 4.969175, 4.969752, 4.970407, 
    4.97306, 4.975472, 4.977946, 4.980508, 4.983161, 4.985892, 4.988606, 
    4.991111, 4.993099, 4.993998, 4.996039, 4.99699, 4.996502, 4.994226, 
    4.989821, 4.983016, 4.97367, 4.961834, 4.947803, 4.932146, 4.915679, 
    4.899399, 4.884381, 4.87164, 4.86201, 4.856055, 4.854027, 4.85586, 
    4.861211,
  // totalHeight(21,39, 0-49)
    4.929265, 4.933565, 4.937625, 4.941379, 4.944791, 4.947852, 4.950571, 
    4.952974, 4.955095, 4.95698, 4.958681, 4.960257, 4.961775, 4.963317, 
    4.964976, 4.964395, 4.967595, 4.96857, 4.969121, 4.969549, 4.97005, 
    4.972878, 4.975447, 4.978108, 4.980676, 4.983141, 4.985444, 4.987503, 
    4.989108, 4.990186, 4.990143, 4.991511, 4.991702, 4.990395, 4.987274, 
    4.982047, 4.974504, 4.964581, 4.952405, 4.938348, 4.923028, 4.907279, 
    4.892075, 4.878423, 4.867244, 4.859259, 4.854925, 4.8544, 4.857553, 
    4.863996,
  // totalHeight(21,40, 0-49)
    4.930509, 4.934163, 4.937672, 4.940976, 4.944041, 4.946851, 4.949409, 
    4.951728, 4.953829, 4.95574, 4.957498, 4.959143, 4.96073, 4.962318, 
    4.963991, 4.96327, 4.967656, 4.968591, 4.969017, 4.969309, 4.969671, 
    4.972606, 4.975278, 4.97807, 4.980577, 4.982781, 4.984569, 4.985875, 
    4.986485, 4.986562, 4.985514, 4.986065, 4.985376, 4.983157, 4.979137, 
    4.973087, 4.964869, 4.954496, 4.942178, 4.928343, 4.913644, 4.898909, 
    4.885057, 4.873009, 4.86357, 4.857339, 4.854666, 4.855622, 4.860014, 
    4.867422,
  // totalHeight(21,41, 0-49)
    4.931998, 4.934996, 4.937942, 4.94078, 4.943478, 4.946014, 4.948385, 
    4.950592, 4.952645, 4.954556, 4.956345, 4.958038, 4.959667, 4.961271, 
    4.962908, 4.962221, 4.967657, 4.968509, 4.968806, 4.968975, 4.969211, 
    4.972187, 4.974899, 4.977754, 4.980126, 4.981987, 4.983173, 4.983639, 
    4.983162, 4.982157, 4.980039, 4.979643, 4.977969, 4.974769, 4.969831, 
    4.962996, 4.954207, 4.943558, 4.931327, 4.917993, 4.904217, 4.890792, 
    4.878562, 4.868335, 4.860787, 4.856392, 4.855388, 4.857768, 4.863286, 
    4.8715,
  // totalHeight(21,42, 0-49)
    4.933681, 4.93602, 4.938399, 4.940762, 4.943074, 4.945315, 4.947473, 
    4.949539, 4.951512, 4.953393, 4.955186, 4.9569, 4.958545, 4.960138, 
    4.961708, 4.961169, 4.967508, 4.968248, 4.968419, 4.968473, 4.968589, 
    4.971543, 4.97423, 4.977072, 4.979232, 4.980669, 4.981169, 4.980713, 
    4.979079, 4.976922, 4.973677, 4.972228, 4.969491, 4.965276, 4.95944, 
    4.951901, 4.942686, 4.931967, 4.920083, 4.907539, 4.894986, 4.883152, 
    4.872786, 4.864562, 4.859018, 4.856503, 4.857143, 4.860859, 4.867363, 
    4.876194,
  // totalHeight(21,43, 0-49)
    4.935478, 4.937166, 4.938977, 4.940857, 4.942774, 4.9447, 4.946618, 
    4.948514, 4.950376, 4.952195, 4.953959, 4.955664, 4.957301, 4.958864, 
    4.960346, 4.960024, 4.967107, 4.967718, 4.967767, 4.967717, 4.967713, 
    4.970584, 4.973182, 4.975931, 4.977798, 4.978734, 4.978477, 4.977031, 
    4.974191, 4.970835, 4.966425, 4.963848, 4.960012, 4.95479, 4.948117, 
    4.939998, 4.930539, 4.919984, 4.908716, 4.897247, 4.886191, 4.876195, 
    4.867887, 4.861801, 4.858331, 4.857696, 4.859924, 4.86486, 4.87218, 
    4.88142,
  // totalHeight(21,44, 0-49)
    4.937275, 4.938323, 4.939574, 4.940974, 4.942487, 4.944084, 4.945742, 
    4.947441, 4.949162, 4.950884, 4.95259, 4.954257, 4.955863, 4.957377, 
    4.958764, 4.958681, 4.966344, 4.966816, 4.966756, 4.966607, 4.966479, 
    4.969213, 4.971659, 4.974236, 4.975735, 4.976098, 4.975027, 4.972552, 
    4.968484, 4.96391, 4.958328, 4.954591, 4.949665, 4.943493, 4.936093, 
    4.927554, 4.91806, 4.907915, 4.897525, 4.887393, 4.878069, 4.8701, 
    4.863985, 4.860114, 4.858732, 4.859934, 4.863651, 4.869663, 4.877614, 
    4.887039,
  // totalHeight(21,45, 0-49)
    4.938926, 4.939353, 4.940056, 4.940982, 4.942094, 4.943354, 4.944736, 
    4.946219, 4.947771, 4.949369, 4.950988, 4.952592, 4.954145, 4.955598, 
    4.956888, 4.957033, 4.965114, 4.965453, 4.965286, 4.965036, 4.964778, 
    4.967328, 4.969562, 4.97189, 4.972956, 4.972693, 4.970773, 4.967258, 
    4.961981, 4.956205, 4.949481, 4.944608, 4.938652, 4.931637, 4.923662, 
    4.914896, 4.905593, 4.896097, 4.886826, 4.878241, 4.870824, 4.865007, 
    4.861149, 4.859497, 4.860159, 4.863107, 4.868181, 4.875099, 4.883481, 
    4.892863,
  // totalHeight(21,46, 0-49)
    4.940262, 4.940084, 4.940259, 4.940728, 4.941444, 4.942371, 4.943476, 
    4.944729, 4.946098, 4.947554, 4.949063, 4.950583, 4.952066, 4.953447, 
    4.954642, 4.95498, 4.963323, 4.963535, 4.963268, 4.96291, 4.962506, 
    4.964828, 4.9668, 4.968812, 4.969393, 4.968471, 4.965699, 4.961167, 
    4.954741, 4.947829, 4.940039, 4.934107, 4.927235, 4.919528, 4.911165, 
    4.902386, 4.893498, 4.884871, 4.876911, 4.870032, 4.864622, 4.861, 
    4.859388, 4.859892, 4.862491, 4.867044, 4.873307, 4.880941, 4.889546, 
    4.898666,
  // totalHeight(21,47, 0-49)
    4.941096, 4.940332, 4.939998, 4.940029, 4.940372, 4.940979, 4.941815, 
    4.942842, 4.944026, 4.945332, 4.94672, 4.948144, 4.949549, 4.950854, 
    4.951961, 4.952435, 4.960899, 4.960996, 4.960621, 4.960141, 4.959572, 
    4.961631, 4.963296, 4.964937, 4.965001, 4.963412, 4.959817, 4.954334, 
    4.946867, 4.938931, 4.930195, 4.923338, 4.915718, 4.907512, 4.898972, 
    4.890397, 4.882132, 4.874554, 4.868045, 4.862955, 4.859578, 4.858113, 
    4.858655, 4.861183, 4.865554, 4.871528, 4.878778, 4.886925, 4.895541, 
    4.904192,
  // totalHeight(21,48, 0-49)
    4.941243, 4.939906, 4.939085, 4.938703, 4.938699, 4.939013, 4.939602, 
    4.940422, 4.941435, 4.942599, 4.943874, 4.945204, 4.946529, 4.947761, 
    4.948786, 4.949333, 4.957789, 4.957774, 4.957283, 4.956659, 4.955901, 
    4.95767, 4.958993, 4.960226, 4.959764, 4.95753, 4.953178, 4.946849, 
    4.938492, 4.929691, 4.920184, 4.91259, 4.904428, 4.895942, 4.887444, 
    4.879278, 4.871814, 4.865419, 4.860435, 4.857142, 4.855741, 4.856319, 
    4.858856, 4.863209, 4.869135, 4.876301, 4.884318, 4.892757, 4.901187, 
    4.909195,
  // totalHeight(21,49, 0-49)
    4.941844, 4.93949, 4.937799, 4.936679, 4.936049, 4.935833, 4.935967, 
    4.936391, 4.937048, 4.937884, 4.938838, 4.939832, 4.94078, 4.941552, 
    4.941981, 4.941836, 4.957452, 4.955976, 4.953788, 4.951624, 4.94955, 
    4.952877, 4.955788, 4.959049, 4.959525, 4.957204, 4.951482, 4.942688, 
    4.930685, 4.918662, 4.906098, 4.898111, 4.889776, 4.881432, 4.873471, 
    4.866293, 4.860284, 4.855782, 4.853061, 4.852297, 4.853556, 4.856781, 
    4.861804, 4.868344, 4.876037, 4.88445, 4.893135, 4.901632, 4.909525, 
    4.916467,
  // totalHeight(22,0, 0-49)
    4.880537, 4.886049, 4.892055, 4.89834, 4.90474, 4.911143, 4.917471, 
    4.923685, 4.92976, 4.935697, 4.941501, 4.947173, 4.952713, 4.958113, 
    4.963342, 4.968148, 4.973527, 4.977929, 4.981947, 4.985516, 4.988526, 
    4.991129, 4.992905, 4.993828, 4.99375, 4.992583, 4.990228, 4.986621, 
    4.981689, 4.975449, 4.967793, 4.959002, 4.948776, 4.937156, 4.924249, 
    4.910238, 4.895406, 4.880136, 4.864914, 4.850298, 4.836879, 4.825234, 
    4.815861, 4.809134, 4.805259, 4.804258, 4.805966, 4.810053, 4.816054, 
    4.823408,
  // totalHeight(22,1, 0-49)
    4.881404, 4.887128, 4.893311, 4.899741, 4.906262, 4.912758, 4.919157, 
    4.925417, 4.93152, 4.937462, 4.943248, 4.948881, 4.954358, 4.959669, 
    4.964782, 4.969224, 4.975, 4.979175, 4.982958, 4.986339, 4.989226, 
    4.992044, 4.994077, 4.995368, 4.995728, 4.995061, 4.993247, 4.99022, 
    4.985889, 4.980306, 4.973286, 4.96537, 4.95594, 4.94499, 4.932577, 
    4.918843, 4.904028, 4.888497, 4.872729, 4.857299, 4.842846, 4.830007, 
    4.819363, 4.81137, 4.806323, 4.804312, 4.805237, 4.808805, 4.814574, 
    4.821985,
  // totalHeight(22,2, 0-49)
    4.882138, 4.888039, 4.894367, 4.900916, 4.907531, 4.914097, 4.920544, 
    4.926829, 4.932936, 4.938857, 4.944596, 4.950159, 4.955542, 4.960733, 
    4.965704, 4.969741, 4.975807, 4.979735, 4.983255, 4.986413, 4.989146, 
    4.992136, 4.994386, 4.996001, 4.99677, 4.996595, 4.995338, 4.992937, 
    4.989284, 4.984453, 4.978187, 4.971295, 4.962846, 4.952787, 4.941124, 
    4.927945, 4.913436, 4.897918, 4.881842, 4.865784, 4.850403, 4.836392, 
    4.824409, 4.815003, 4.808563, 4.805276, 4.805117, 4.807853, 4.813084, 
    4.820271,
  // totalHeight(22,3, 0-49)
    4.88286, 4.888899, 4.895341, 4.901977, 4.908658, 4.915267, 4.921736, 
    4.92802, 4.9341, 4.93997, 4.945633, 4.951095, 4.956351, 4.961398, 
    4.966206, 4.969803, 4.976026, 4.979697, 4.982938, 4.98585, 4.988398, 
    4.991513, 4.99393, 4.995817, 4.996953, 4.997241, 4.996539, 4.994784, 
    4.991858, 4.987838, 4.982406, 4.976634, 4.969298, 4.960302, 4.949604, 
    4.937222, 4.923286, 4.908053, 4.891929, 4.875461, 4.859316, 4.844221, 
    4.830904, 4.820007, 4.812023, 4.807248, 4.80575, 4.807377, 4.811787, 
    4.818478,
  // totalHeight(22,4, 0-49)
    4.883684, 4.889828, 4.896346, 4.903038, 4.90975, 4.916372, 4.922831, 
    4.929082, 4.935105, 4.940893, 4.946448, 4.951777, 4.956883, 4.96176, 
    4.966392, 4.969527, 4.975749, 4.97916, 4.982116, 4.984766, 4.987107, 
    4.990293, 4.992825, 4.99492, 4.996367, 4.997078, 4.996912, 4.995807, 
    4.993631, 4.990452, 4.985897, 4.981287, 4.975144, 4.96733, 4.957751, 
    4.94637, 4.93324, 4.918549, 4.902637, 4.886006, 4.869302, 4.853272, 
    4.838696, 4.826305, 4.8167, 4.810288, 4.807254, 4.807538, 4.810874, 
    4.816814,
  // totalHeight(22,5, 0-49)
    4.884719, 4.890928, 4.897486, 4.904196, 4.910906, 4.917505, 4.92392, 
    4.930103, 4.936036, 4.941709, 4.947129, 4.952298, 4.957226, 4.961914, 
    4.96636, 4.969028, 4.97508, 4.978233, 4.980904, 4.983284, 4.985404, 
    4.98861, 4.991196, 4.993429, 4.995127, 4.99621, 4.996547, 4.996074, 
    4.994657, 4.992321, 4.988653, 4.985206, 4.980282, 4.973714, 4.96536, 
    4.955123, 4.942988, 4.929064, 4.913613, 4.897071, 4.880046, 4.86328, 
    4.847586, 4.833769, 4.822536, 4.814412, 4.809701, 4.80846, 4.81051, 
    4.815478,
  // totalHeight(22,6, 0-49)
    4.886049, 4.892287, 4.898846, 4.905535, 4.912204, 4.918742, 4.925076, 
    4.931158, 4.936968, 4.942498, 4.947752, 4.952737, 4.957466, 4.961949, 
    4.9662, 4.968412, 4.974121, 4.97702, 4.979414, 4.981527, 4.983417, 
    4.986587, 4.98917, 4.991468, 4.99335, 4.994747, 4.995544, 4.99568, 
    4.995009, 4.993502, 4.990707, 4.988382, 4.984662, 4.979352, 4.972273, 
    4.963274, 4.952274, 4.9393, 4.924531, 4.908326, 4.89123, 4.873957, 
    4.857336, 4.842224, 4.829421, 4.819574, 4.813116, 4.810222, 4.810823, 
    4.814631,
  // totalHeight(22,7, 0-49)
    4.887733, 4.893962, 4.900485, 4.907114, 4.913703, 4.920143, 4.92636, 
    4.932308, 4.937963, 4.94332, 4.948382, 4.953161, 4.957674, 4.961939, 
    4.965983, 4.967781, 4.972977, 4.975623, 4.977752, 4.979605, 4.981266, 
    4.984348, 4.986871, 4.989161, 4.991158, 4.992808, 4.994019, 4.994727, 
    4.994781, 4.994075, 4.992127, 4.990852, 4.98828, 4.984199, 4.978396, 
    4.970678, 4.960901, 4.949014, 4.935112, 4.919465, 4.902544, 4.885012, 
    4.867685, 4.851458, 4.837206, 4.825689, 4.817468, 4.812854, 4.811893, 
    4.814398,
  // totalHeight(22,8, 0-49)
    4.88981, 4.895993, 4.902441, 4.908971, 4.915441, 4.921747, 4.927812, 
    4.933593, 4.939067, 4.944226, 4.949075, 4.953628, 4.957908, 4.96194, 
    4.965762, 4.967212, 4.971738, 4.974128, 4.976008, 4.977619, 4.979063, 
    4.982004, 4.98441, 4.986624, 4.988671, 4.990512, 4.992086, 4.993325, 
    4.994076, 4.994135, 4.992996, 4.992678, 4.991173, 4.988257, 4.983695, 
    4.977253, 4.968738, 4.958027, 4.945134, 4.930234, 4.913712, 4.896164, 
    4.878372, 4.86124, 4.845705, 4.832624, 4.822687, 4.816338, 4.813755, 
    4.814858,
  // totalHeight(22,9, 0-49)
    4.892284, 4.898389, 4.904727, 4.911123, 4.917439, 4.923574, 4.929457, 
    4.935043, 4.94031, 4.945249, 4.949864, 4.954177, 4.958208, 4.96199, 
    4.965567, 4.966765, 4.970487, 4.972616, 4.974267, 4.975658, 4.976905, 
    4.979655, 4.981893, 4.983966, 4.986002, 4.987977, 4.989863, 4.991588, 
    4.993001, 4.993782, 4.993412, 4.993945, 4.993408, 4.991569, 4.988178, 
    4.982973, 4.975715, 4.966225, 4.954433, 4.940427, 4.924498, 4.90716, 
    4.889142, 4.871335, 4.854712, 4.84022, 4.828661, 4.820616, 4.8164, 
    4.816047,
  // totalHeight(22,10, 0-49)
    4.895145, 4.901142, 4.907338, 4.913567, 4.919698, 4.925632, 4.931304, 
    4.93667, 4.941706, 4.946405, 4.950773, 4.95483, 4.958596, 4.96211, 
    4.965409, 4.96648, 4.969285, 4.971148, 4.972591, 4.973794, 4.974871, 
    4.977384, 4.979412, 4.981291, 4.983261, 4.985313, 4.987463, 4.989625, 
    4.991659, 4.993119, 4.993484, 4.99475, 4.995069, 4.994203, 4.991892, 
    4.987855, 4.981818, 4.973549, 4.96291, 4.949902, 4.93472, 4.917789, 
    4.899768, 4.881516, 4.864025, 4.8483, 4.835255, 4.825601, 4.819786, 
    4.817967,
  // totalHeight(22,11, 0-49)
    4.898359, 4.904222, 4.910252, 4.916286, 4.922204, 4.927913, 4.93335, 
    4.938472, 4.943258, 4.947702, 4.951809, 4.955594, 4.959082, 4.962301, 
    4.965283, 4.966367, 4.968176, 4.969769, 4.971031, 4.972083, 4.973031, 
    4.975266, 4.977045, 4.978685, 4.980544, 4.98263, 4.984991, 4.987542, 
    4.990149, 4.992247, 4.993314, 4.995196, 4.996253, 4.996246, 4.994911, 
    4.991952, 4.987071, 4.979993, 4.970516, 4.958566, 4.944244, 4.927882, 
    4.910058, 4.891582, 4.873441, 4.856687, 4.842321, 4.831179, 4.823837, 
    4.82058,
  // totalHeight(22,12, 0-49)
    4.901878, 4.907592, 4.913434, 4.919252, 4.924936, 4.930398, 4.935579, 
    4.940441, 4.944962, 4.949134, 4.952963, 4.956466, 4.959656, 4.962557, 
    4.965181, 4.966418, 4.967177, 4.968506, 4.96962, 4.970567, 4.97143, 
    4.973352, 4.974858, 4.976231, 4.977943, 4.980022, 4.98255, 4.985436, 
    4.988568, 4.991255, 4.992997, 4.995377, 4.997054, 4.99779, 4.997318, 
    4.995336, 4.991525, 4.98558, 4.977245, 4.966374, 4.952986, 4.937315, 
    4.919857, 4.901359, 4.882782, 4.865209, 4.849709, 4.837227, 4.828466, 
    4.823829,
  // totalHeight(22,13, 0-49)
    4.90565, 4.911202, 4.916841, 4.922431, 4.927863, 4.933063, 4.937972, 
    4.942556, 4.946795, 4.950685, 4.954226, 4.957429, 4.960305, 4.962861, 
    4.96509, 4.966601, 4.96628, 4.967366, 4.968375, 4.969272, 4.970106, 
    4.971691, 4.97291, 4.973999, 4.975545, 4.977583, 4.980232, 4.9834, 
    4.986999, 4.990225, 4.992621, 4.995386, 4.997564, 4.998925, 4.999202, 
    4.998087, 4.99525, 4.990359, 4.983118, 4.973319, 4.960899, 4.946009, 
    4.92905, 4.910706, 4.891897, 4.873711, 4.857275, 4.843622, 4.83357, 
    4.827637,
  // totalHeight(22,14, 0-49)
    4.909611, 4.915001, 4.920432, 4.925782, 4.930954, 4.935875, 4.940499, 
    4.944792, 4.948737, 4.952328, 4.955569, 4.958461, 4.961009, 4.963201, 
    4.965012, 4.966866, 4.965448, 4.966335, 4.967295, 4.968207, 4.969079, 
    4.970313, 4.971245, 4.97205, 4.973421, 4.975398, 4.978127, 4.981521, 
    4.985519, 4.989235, 4.992261, 4.995299, 4.997867, 4.999737, 5.000646, 
    5.000288, 4.998318, 4.994392, 4.988178, 4.979414, 4.96797, 4.953912, 
    4.937561, 4.919518, 4.900659, 4.882061, 4.864886, 4.850241, 4.839045, 
    4.831921,
  // totalHeight(22,15, 0-49)
    4.913706, 4.918937, 4.924161, 4.929266, 4.934164, 4.938797, 4.943122, 
    4.947111, 4.950749, 4.954034, 4.956963, 4.959537, 4.961747, 4.96357, 
    4.964959, 4.967154, 4.964622, 4.965373, 4.966358, 4.967362, 4.968349, 
    4.96923, 4.969894, 4.970437, 4.971638, 4.973541, 4.976313, 4.979875, 
    4.984203, 4.988347, 4.99198, 4.995186, 4.998031, 5.000298, 5.001725, 
    5.002008, 5.000802, 4.997742, 4.992472, 4.984691, 4.974206, 4.96101, 
    4.945339, 4.927721, 4.908974, 4.89015, 4.87243, 4.856977, 4.844789, 
    4.836594,
  // totalHeight(22,16, 0-49)
    4.917878, 4.922956, 4.927972, 4.932827, 4.937447, 4.94178, 4.945793, 
    4.949466, 4.952789, 4.95576, 4.958376, 4.960632, 4.962512, 4.963979, 
    4.964971, 4.967404, 4.963717, 4.964427, 4.965526, 4.966713, 4.967906, 
    4.968447, 4.96888, 4.969199, 4.970256, 4.972084, 4.974867, 4.978536, 
    4.983116, 4.987617, 4.991826, 4.995096, 4.998113, 5.000667, 5.002501, 
    5.003314, 5.00276, 5.000465, 4.996054, 4.989187, 4.979626, 4.967295, 
    4.952357, 4.935261, 4.916767, 4.897888, 4.879806, 4.863722, 4.850706, 
    4.841565,
  // totalHeight(22,17, 0-49)
    4.92207, 4.926999, 4.931807, 4.936404, 4.940733, 4.944755, 4.948444, 
    4.951794, 4.9548, 4.957461, 4.959776, 4.961733, 4.963308, 4.964456, 
    4.965109, 4.967572, 4.962652, 4.963425, 4.964743, 4.966219, 4.967717, 
    4.967952, 4.96821, 4.968366, 4.96932, 4.971087, 4.973859, 4.977577, 
    4.982324, 4.9871, 4.991838, 4.99507, 4.998154, 5.000888, 5.00302, 
    5.004251, 5.00424, 5.002608, 4.998962, 4.992938, 4.984252, 4.972774, 
    4.9586, 4.942105, 4.923982, 4.905201, 4.886931, 4.870391, 4.856705, 
    4.846749,
  // totalHeight(22,18, 0-49)
    4.926219, 4.930993, 4.935577, 4.939902, 4.943923, 4.94762, 4.950982, 
    4.954012, 4.956714, 4.95909, 4.961139, 4.96284, 4.964164, 4.96506, 
    4.965462, 4.967654, 4.961352, 4.962304, 4.963949, 4.965824, 4.967738, 
    4.967719, 4.967881, 4.967954, 4.96887, 4.970606, 4.973351, 4.977064, 
    4.981887, 4.986845, 4.99204, 4.995138, 4.998181, 5.000986, 5.003305, 
    5.004848, 5.005273, 5.004199, 5.001225, 4.995965, 4.988102, 4.977455, 
    4.964059, 4.948224, 4.930574, 4.912029, 4.893728, 4.876899, 4.862697, 
    4.852058,
  // totalHeight(22,19, 0-49)
    4.930254, 4.934838, 4.939164, 4.943184, 4.946876, 4.950236, 4.953277, 
    4.95601, 4.958449, 4.960598, 4.962448, 4.963972, 4.965132, 4.96587, 
    4.966131, 4.967701, 4.959782, 4.961017, 4.963089, 4.965472, 4.967917, 
    4.967721, 4.967884, 4.967977, 4.968936, 4.970692, 4.973415, 4.977076, 
    4.981885, 4.986914, 4.992465, 4.995318, 4.998209, 5.000971, 5.003365, 
    5.005108, 5.005862, 5.005246, 5.002851, 4.998276, 4.991178, 4.981333, 
    4.968722, 4.953592, 4.936501, 4.918311, 4.900126, 4.883163, 4.868595, 
    4.857404,
  // totalHeight(22,20, 0-49)
    4.935121, 4.940522, 4.945562, 4.95019, 4.954374, 4.958099, 4.961357, 
    4.964148, 4.966482, 4.968373, 4.969851, 4.970959, 4.971753, 4.972302, 
    4.972693, 30, 4.959976, 4.961293, 4.963098, 4.965001, 4.966878, 4.965349, 
    4.964415, 4.963618, 4.964009, 4.965533, 4.968349, 4.972388, 4.97783, 
    4.983681, 4.990357, 4.993667, 4.997002, 5.000195, 5.003012, 5.00518, 
    5.006382, 5.006256, 5.004407, 5.000442, 4.994011, 4.984875, 4.972975, 
    4.958509, 4.941978, 4.924188, 4.906198, 4.8892, 4.874375, 4.862727,
  // totalHeight(22,21, 0-49)
    4.939007, 4.944368, 4.949268, 4.953667, 4.957558, 4.960947, 4.963851, 
    4.966298, 4.968316, 4.969938, 4.971203, 4.972163, 4.972878, 4.973427, 
    4.973916, 30, 4.955731, 4.957488, 4.959795, 4.962227, 4.964609, 4.962763, 
    4.96166, 4.960739, 4.961128, 4.962759, 4.965786, 4.970114, 4.975934, 
    4.982237, 4.989596, 4.992975, 4.996485, 4.999949, 5.003128, 5.00574, 
    5.007459, 5.007914, 5.006705, 5.003426, 4.997713, 4.989299, 4.978093, 
    4.964244, 4.948203, 4.930723, 4.912822, 4.895671, 4.880454, 4.868197,
  // totalHeight(22,22, 0-49)
    4.942727, 4.948107, 4.952914, 4.957129, 4.960762, 4.96384, 4.966405, 
    4.968505, 4.970191, 4.971513, 4.972527, 4.973292, 4.973882, 4.974389, 
    4.974936, 30, 4.952352, 4.954473, 4.957218, 4.960129, 4.962974, 4.960836, 
    4.959574, 4.958531, 4.958904, 4.960607, 4.963778, 4.968307, 4.974384, 
    4.980988, 4.988835, 4.992147, 4.995678, 4.999262, 5.002652, 5.005566, 
    5.007674, 5.008605, 5.007951, 5.005296, 5.000262, 4.99256, 4.982064, 
    4.968881, 4.953407, 4.936348, 4.918674, 4.901524, 4.886073, 4.873363,
  // totalHeight(22,23, 0-49)
    4.946211, 4.951646, 4.956401, 4.960465, 4.963868, 4.966659, 4.968901, 
    4.970664, 4.972017, 4.973031, 4.973774, 4.974321, 4.974754, 4.975182, 
    4.975747, 30, 4.949856, 4.952229, 4.955276, 4.958517, 4.961682, 4.959258, 
    4.957822, 4.956636, 4.956953, 4.958671, 4.961921, 4.966574, 4.97282, 
    4.979625, 4.98781, 4.991016, 4.994521, 4.998165, 5.001703, 5.004858, 
    5.007296, 5.008648, 5.0085, 5.006428, 5.002038, 4.995022, 4.98522, 
    4.972703, 4.957818, 4.94122, 4.923836, 4.906774, 4.891189, 4.878129,
  // totalHeight(22,24, 0-49)
    4.949394, 4.954908, 4.959633, 4.963575, 4.966775, 4.969305, 4.971246, 
    4.972689, 4.973722, 4.97443, 4.9749, 4.975216, 4.975473, 4.975791, 
    4.976331, 30, 4.948518, 4.951012, 4.954212, 4.957628, 4.960968, 4.958356, 
    4.95681, 4.955535, 4.955814, 4.957535, 4.960822, 4.965538, 4.971878, 
    4.978793, 4.987182, 4.990316, 4.993803, 4.997482, 5.001118, 5.004433, 
    5.007102, 5.008749, 5.008963, 5.007317, 5.003409, 4.996915, 4.987658, 
    4.975676, 4.961286, 4.945103, 4.928017, 4.911108, 4.895511, 4.882263,
  // totalHeight(22,25, 0-49)
    4.952204, 4.957809, 4.962523, 4.966364, 4.969392, 4.971691, 4.973362, 
    4.97451, 4.975244, 4.975662, 4.975863, 4.975944, 4.97601, 4.976191, 
    4.976657, 30, 4.948055, 4.950538, 4.953739, 4.957167, 4.960527, 4.957858, 
    4.956294, 4.955017, 4.955307, 4.957049, 4.960361, 4.965107, 4.971481, 
    4.978438, 4.986895, 4.990032, 4.993546, 4.99728, 5.001002, 5.004436, 
    5.00726, 5.0091, 5.009548, 5.008173, 5.004572, 4.998418, 4.989519, 
    4.977905, 4.96387, 4.948008, 4.931185, 4.914455, 4.898934, 4.885649,
  // totalHeight(22,26, 0-49)
    4.95458, 4.960278, 4.964995, 4.96876, 4.971643, 4.973747, 4.975185, 
    4.976077, 4.97654, 4.97669, 4.976631, 4.976472, 4.976333, 4.976344, 
    4.976682, 30, 4.948453, 4.950796, 4.953845, 4.957116, 4.960338, 4.957754, 
    4.956271, 4.955087, 4.95545, 4.95724, 4.960577, 4.965328, 4.97169, 
    4.978623, 4.98702, 4.990255, 4.993862, 4.997688, 5.001496, 5.005016, 
    5.007926, 5.009855, 5.010394, 5.00912, 5.00563, 4.999599, 4.990843, 
    4.979391, 4.965537, 4.949868, 4.933245, 4.916705, 4.901348, 4.888179,
  // totalHeight(22,27, 0-49)
    4.95647, 4.962255, 4.966988, 4.970704, 4.973483, 4.975435, 4.976684, 
    4.977357, 4.977584, 4.977483, 4.977173, 4.976769, 4.976398, 4.976196, 
    4.976342, 30, 4.94983, 4.951895, 4.954633, 4.957582, 4.960505, 4.958111, 
    4.956778, 4.955749, 4.956214, 4.95806, 4.961405, 4.966125, 4.972418, 
    4.979264, 4.98748, 4.990894, 4.994651, 4.998594, 5.002487, 5.006057, 
    5.008984, 5.010896, 5.011392, 5.010053, 5.006485, 5.000376, 4.991556, 
    4.98007, 4.96623, 4.950636, 4.934154, 4.917815, 4.902705, 4.889807,
  // totalHeight(22,28, 0-49)
    4.957836, 4.963705, 4.968472, 4.972172, 4.974893, 4.976745, 4.977857, 
    4.978356, 4.978376, 4.978041, 4.977476, 4.976804, 4.976159, 4.975689, 
    4.975567, 30, 4.952566, 4.954219, 4.956491, 4.958948, 4.961411, 4.95925, 
    4.958077, 4.957208, 4.95776, 4.959622, 4.962923, 4.967553, 4.973707, 
    4.980392, 4.988312, 4.991958, 4.995893, 4.999952, 5.003895, 5.00745, 
    5.010296, 5.012068, 5.012367, 5.010787, 5.006949, 5.000559, 4.991478, 
    4.979781, 4.965812, 4.950198, 4.933821, 4.917719, 4.90296, 4.890495,
  // totalHeight(22,29, 0-49)
    4.95867, 4.964626, 4.969453, 4.973186, 4.975905, 4.977718, 4.978745, 
    4.979113, 4.978947, 4.978374, 4.97753, 4.976545, 4.975567, 4.974751, 
    4.974271, 30, 4.95646, 4.95757, 4.959221, 4.961021, 4.962852, 4.960859, 
    4.959756, 4.958962, 4.95951, 4.961305, 4.96448, 4.968947, 4.974889, 
    4.981332, 4.988841, 4.992712, 4.996807, 5.000953, 5.004909, 5.008403, 
    5.011117, 5.012687, 5.012722, 5.010827, 5.006638, 4.999887, 4.990465, 
    4.978487, 4.964337, 4.94868, 4.932421, 4.916602, 4.902275, 4.890357,
  // totalHeight(22,30, 0-49)
    4.958047, 4.963116, 4.967086, 4.970015, 4.972012, 4.973216, 4.973781, 
    4.973852, 4.973566, 4.973029, 4.972315, 4.97146, 4.970461, 4.969284, 
    4.96787, 4.971422, 4.957416, 4.958146, 4.959991, 4.962359, 4.964968, 
    4.964603, 4.964927, 4.965328, 4.966667, 4.968801, 4.971864, 4.975824, 
    4.980929, 4.98633, 4.992523, 4.995769, 4.999239, 5.002778, 5.006158, 
    5.009108, 5.011305, 5.01238, 5.011932, 5.009561, 5.00491, 4.997726, 
    4.987928, 4.975666, 4.961368, 4.945735, 4.929695, 4.914293, 4.900559, 
    4.889373,
  // totalHeight(22,31, 0-49)
    4.95789, 4.963067, 4.967144, 4.970172, 4.972244, 4.973488, 4.974046, 
    4.974065, 4.973676, 4.972998, 4.972118, 4.97109, 4.969933, 4.968622, 
    4.967101, 4.971066, 4.959039, 4.959276, 4.960526, 4.96225, 4.964221, 
    4.963971, 4.964255, 4.964615, 4.965906, 4.968037, 4.971161, 4.975234, 
    4.980437, 4.98588, 4.991862, 4.995546, 4.999402, 5.003253, 5.00686, 
    5.009934, 5.012142, 5.013105, 5.012422, 5.009698, 5.004597, 4.9969, 
    4.986571, 4.973823, 4.959142, 4.94329, 4.927226, 4.912013, 4.898664, 
    4.888015,
  // totalHeight(22,32, 0-49)
    4.957166, 4.962335, 4.966437, 4.969514, 4.971652, 4.972965, 4.973582, 
    4.97364, 4.973271, 4.972588, 4.971687, 4.970632, 4.969455, 4.968151, 
    4.96666, 4.970359, 4.96031, 4.960156, 4.960892, 4.962051, 4.963462, 
    4.963401, 4.963728, 4.964138, 4.96545, 4.967617, 4.970803, 4.974948, 
    4.980169, 4.985564, 4.991252, 4.995315, 4.999488, 5.003579, 5.007331, 
    5.010444, 5.012566, 5.013313, 5.012284, 5.009094, 5.003433, 4.995127, 
    4.984194, 4.970913, 4.955841, 4.939794, 4.923772, 4.908843, 4.895998, 
    4.886026,
  // totalHeight(22,33, 0-49)
    4.955983, 4.961055, 4.965122, 4.968218, 4.970413, 4.971811, 4.972531, 
    4.972694, 4.972424, 4.971832, 4.971011, 4.970033, 4.968942, 4.967745, 
    4.966402, 4.969375, 4.961257, 4.960827, 4.96114, 4.961818, 4.962752, 
    4.962927, 4.963367, 4.963902, 4.965289, 4.967519, 4.970751, 4.974916, 
    4.980073, 4.985337, 4.990673, 4.995048, 4.999469, 5.003721, 5.007534, 
    5.010592, 5.01253, 5.012957, 5.011473, 5.007711, 5.001394, 4.992397, 
    4.980807, 4.966975, 4.951529, 4.935343, 4.919448, 4.904913, 4.892695, 
    4.883534,
  // totalHeight(22,34, 0-49)
    4.954448, 4.95936, 4.963346, 4.966434, 4.968682, 4.970178, 4.971027, 
    4.971339, 4.971222, 4.970782, 4.970108, 4.969277, 4.968343, 4.967324, 
    4.966204, 4.968204, 4.961935, 4.961338, 4.961315, 4.96159, 4.962114, 
    4.962554, 4.963157, 4.963874, 4.965377, 4.967681, 4.970933, 4.975061, 
    4.980067, 4.985126, 4.99007, 4.994689, 4.999281, 5.003613, 5.007399, 
    5.010306, 5.01196, 5.011963, 5.009924, 5.005498, 4.998452, 4.988713, 
    4.976445, 4.962076, 4.946308, 4.930067, 4.914408, 4.900389, 4.888928, 
    4.880701,
  // totalHeight(22,35, 0-49)
    4.952672, 4.957375, 4.961246, 4.964301, 4.966592, 4.968191, 4.969186, 
    4.969673, 4.969746, 4.969497, 4.969015, 4.968374, 4.967635, 4.966836, 
    4.965979, 4.966949, 4.962429, 4.961751, 4.961463, 4.961401, 4.961579, 
    4.962293, 4.96309, 4.964033, 4.965674, 4.968048, 4.971286, 4.975313, 
    4.980082, 4.984866, 4.989388, 4.994173, 4.99885, 5.00317, 5.006832, 
    5.00949, 5.010759, 5.010242, 5.00756, 5.002398, 4.994569, 4.984073, 
    4.971148, 4.9563, 4.940302, 4.924123, 4.908833, 4.895466, 4.88489, 
    4.877709,
  // totalHeight(22,36, 0-49)
    4.950771, 4.955221, 4.958945, 4.961947, 4.96427, 4.965969, 4.967115, 
    4.96779, 4.968071, 4.968041, 4.967778, 4.967352, 4.96683, 4.966259, 
    4.965673, 4.965696, 4.962821, 4.962123, 4.961627, 4.961285, 4.961173, 
    4.96215, 4.963158, 4.96435, 4.96614, 4.968571, 4.97175, 4.975606, 
    4.980051, 4.984489, 4.988561, 4.993416, 4.99808, 5.002285, 5.005719, 
    5.008024, 5.008811, 5.007683, 5.004285, 4.998341, 4.98972, 4.978488, 
    4.96497, 4.949749, 4.933655, 4.917694, 4.902929, 4.890361, 4.880794, 
    4.874759,
  // totalHeight(22,37, 0-49)
    4.948856, 4.953017, 4.956562, 4.959488, 4.961827, 4.963615, 4.964911, 
    4.965777, 4.966276, 4.966475, 4.966443, 4.966245, 4.965945, 4.9656, 
    4.965266, 4.964514, 4.963181, 4.962499, 4.961835, 4.961262, 4.960908, 
    4.962128, 4.963348, 4.964801, 4.966734, 4.969196, 4.972267, 4.975879, 
    4.979912, 4.983932, 4.987516, 4.992332, 4.996866, 5.000842, 5.003934, 
    5.005777, 5.005983, 5.004169, 5.000006, 4.993264, 4.983874, 4.971982, 
    4.957987, 4.942545, 4.926535, 4.910977, 4.896918, 4.885301, 4.876864, 
    4.872054,
  // totalHeight(22,38, 0-49)
    4.947029, 4.95087, 4.954208, 4.957035, 4.959365, 4.961228, 4.962661, 
    4.96371, 4.964424, 4.964855, 4.965057, 4.965089, 4.965008, 4.964876, 
    4.964758, 4.963451, 4.963553, 4.962902, 4.962105, 4.961343, 4.960793, 
    4.962229, 4.963652, 4.965358, 4.967416, 4.969876, 4.972776, 4.976065, 
    4.979594, 4.983118, 4.98617, 4.990817, 4.995093, 4.99871, 5.00134, 
    5.002613, 5.00215, 4.999588, 4.994634, 4.987115, 4.977029, 4.964597, 
    4.950294, 4.934833, 4.919126, 4.904189, 4.891028, 4.880522, 4.873323, 
    4.869796,
  // totalHeight(22,39, 0-49)
    4.945388, 4.948878, 4.95198, 4.954679, 4.956977, 4.958889, 4.960439, 
    4.961655, 4.962572, 4.963227, 4.96366, 4.963917, 4.964046, 4.964107, 
    4.964168, 4.96253, 4.963966, 4.963343, 4.962438, 4.96153, 4.960828, 
    4.962446, 4.964049, 4.965991, 4.968144, 4.970555, 4.973221, 4.976102, 
    4.979031, 4.981975, 4.984433, 4.988768, 4.992643, 4.995764, 4.997804, 
    4.9984, 4.997189, 4.993839, 4.988104, 4.979869, 4.969203, 4.956405, 
    4.94201, 4.926777, 4.911627, 4.89755, 4.885493, 4.876248, 4.870383, 
    4.868177,
  // totalHeight(22,40, 0-49)
    4.944005, 4.947119, 4.949958, 4.952499, 4.954735, 4.956668, 4.958309, 
    4.959668, 4.960769, 4.96163, 4.962281, 4.962752, 4.96308, 4.963314, 
    4.963518, 4.961757, 4.964414, 4.963816, 4.962826, 4.961812, 4.960998, 
    4.962762, 4.964519, 4.966666, 4.968871, 4.971179, 4.973535, 4.975921, 
    4.978155, 4.980425, 4.982213, 4.986079, 4.989399, 4.99188, 4.993204, 
    4.993023, 4.991001, 4.986851, 4.980374, 4.971526, 4.960449, 4.947505, 
    4.933281, 4.918559, 4.904246, 4.891278, 4.880527, 4.87269, 4.868237, 
    4.867364,
  // totalHeight(22,41, 0-49)
    4.942934, 4.945651, 4.948199, 4.950552, 4.952695, 4.954617, 4.956311, 
    4.957786, 4.959041, 4.960086, 4.960935, 4.961604, 4.962116, 4.962505, 
    4.962822, 4.961109, 4.964873, 4.964289, 4.963243, 4.96216, 4.961271, 
    4.963148, 4.965024, 4.967335, 4.969543, 4.971682, 4.973652, 4.975451, 
    4.976894, 4.978395, 4.979421, 4.98265, 4.985257, 4.986954, 4.987439, 
    4.986394, 4.983522, 4.978585, 4.971448, 4.962138, 4.950858, 4.938031, 
    4.924275, 4.910371, 4.897185, 4.885581, 4.876331, 4.870027, 4.86704, 
    4.867486,
  // totalHeight(22,42, 0-49)
    4.942198, 4.944501, 4.946737, 4.948874, 4.950887, 4.952759, 4.954475, 
    4.956024, 4.957401, 4.9586, 4.959621, 4.960468, 4.961146, 4.961676, 
    4.962083, 4.960546, 4.965296, 4.964724, 4.963648, 4.962533, 4.961604, 
    4.963559, 4.96552, 4.967943, 4.970094, 4.971998, 4.973501, 4.974625, 
    4.975183, 4.975811, 4.975973, 4.978401, 4.980134, 4.980906, 4.980445, 
    4.978471, 4.974735, 4.969062, 4.961384, 4.951796, 4.940564, 4.928149, 
    4.91518, 4.90241, 4.890639, 4.880638, 4.873065, 4.868399, 4.866908, 
    4.868633,
  // totalHeight(22,43, 0-49)
    4.941798, 4.943673, 4.945574, 4.947466, 4.949317, 4.951102, 4.952796, 
    4.954382, 4.95584, 4.957156, 4.958319, 4.959318, 4.960145, 4.9608, 
    4.961287, 4.960012, 4.965619, 4.965061, 4.963984, 4.962872, 4.961929, 
    4.963934, 4.965942, 4.968421, 4.970454, 4.972047, 4.973005, 4.973367, 
    4.972955, 4.97261, 4.971803, 4.973268, 4.973981, 4.973707, 4.972209, 
    4.969264, 4.964683, 4.958358, 4.950296, 4.940651, 4.929743, 4.918052, 
    4.906193, 4.894865, 4.884781, 4.876598, 4.870849, 4.867894, 4.867904, 
    4.870842,
  // totalHeight(22,44, 0-49)
    4.941687, 4.943127, 4.944678, 4.9463, 4.947957, 4.949617, 4.95125, 
    4.952827, 4.954327, 4.955722, 4.956991, 4.958113, 4.959068, 4.959835, 
    4.960393, 4.959428, 4.965758, 4.965227, 4.96418, 4.963101, 4.962169, 
    4.964197, 4.966213, 4.968689, 4.970536, 4.971749, 4.972087, 4.97161, 
    4.970154, 4.968743, 4.966866, 4.967227, 4.966793, 4.965372, 4.962781, 
    4.958857, 4.953483, 4.946626, 4.938364, 4.928908, 4.918612, 4.907955, 
    4.897513, 4.88791, 4.87975, 4.87356, 4.869744, 4.868541, 4.870022, 
    4.874084,
  // totalHeight(22,45, 0-49)
    4.941793, 4.942795, 4.943985, 4.945317, 4.946753, 4.948253, 4.949785, 
    4.951314, 4.952811, 4.954244, 4.955584, 4.9568, 4.957859, 4.958724, 
    4.959352, 4.958708, 4.965632, 4.96514, 4.964149, 4.963128, 4.962224, 
    4.964252, 4.966239, 4.96865, 4.97025, 4.971015, 4.97067, 4.969294, 
    4.966736, 4.964185, 4.961152, 4.960292, 4.958618, 4.955986, 4.952279, 
    4.947404, 4.941326, 4.934086, 4.92583, 4.916817, 4.907412, 4.898078, 
    4.889328, 4.881688, 4.875639, 4.87157, 4.869749, 4.870298, 4.873192, 
    4.878266,
  // totalHeight(22,46, 0-49)
    4.942007, 4.942574, 4.943394, 4.944422, 4.945613, 4.946927, 4.948323, 
    4.949766, 4.951222, 4.952654, 4.954029, 4.955307, 4.956448, 4.957397, 
    4.958094, 4.957758, 4.965144, 4.964711, 4.963798, 4.962851, 4.961987, 
    4.963995, 4.965917, 4.968205, 4.969499, 4.96976, 4.968681, 4.966363, 
    4.962676, 4.958935, 4.954689, 4.952533, 4.949564, 4.9457, 4.940897, 
    4.935141, 4.928477, 4.921025, 4.91299, 4.904661, 4.896404, 4.888639, 
    4.881803, 4.876304, 4.87249, 4.870608, 4.870795, 4.873055, 4.877275, 
    4.88323,
  // totalHeight(22,47, 0-49)
    4.942184, 4.942324, 4.942777, 4.943493, 4.944427, 4.94553, 4.946764, 
    4.948091, 4.949472, 4.950871, 4.952249, 4.95356, 4.954759, 4.955781, 
    4.956546, 4.956481, 4.964205, 4.963849, 4.963029, 4.962167, 4.961345, 
    4.963313, 4.965137, 4.967248, 4.968189, 4.967905, 4.966066, 4.96279, 
    4.957972, 4.953028, 4.947546, 4.944068, 4.939801, 4.934735, 4.928899, 
    4.922368, 4.915265, 4.907782, 4.900171, 4.892743, 4.885846, 4.879838, 
    4.875064, 4.87181, 4.870286, 4.870596, 4.872749, 4.876638, 4.882066, 
    4.888757,
  // totalHeight(22,48, 0-49)
    4.942157, 4.941879, 4.941971, 4.942379, 4.943048, 4.943933, 4.94499, 
    4.94618, 4.947465, 4.948805, 4.95016, 4.951481, 4.952719, 4.953801, 
    4.954633, 4.95479, 4.962732, 4.962471, 4.961751, 4.960971, 4.960187, 
    4.962099, 4.963796, 4.965682, 4.966233, 4.965381, 4.962782, 4.958564, 
    4.952653, 4.946531, 4.939835, 4.935065, 4.929556, 4.923367, 4.916611, 
    4.909441, 4.902061, 4.894722, 4.887719, 4.881363, 4.875974, 4.871838, 
    4.869196, 4.86821, 4.868954, 4.871396, 4.875418, 4.880815, 4.887309, 
    4.894578,
  // totalHeight(22,49, 0-49)
    4.942302, 4.941273, 4.940712, 4.94055, 4.940726, 4.94118, 4.941866, 
    4.942734, 4.943739, 4.944835, 4.945973, 4.947086, 4.948108, 4.94893, 
    4.949424, 4.949001, 4.964243, 4.962885, 4.960816, 4.958843, 4.957083, 
    4.960893, 4.964464, 4.968607, 4.970275, 4.969415, 4.9654, 4.958524, 
    4.948629, 4.938767, 4.928291, 4.922237, 4.915466, 4.908151, 4.900531, 
    4.892879, 4.885505, 4.878732, 4.872895, 4.868293, 4.865188, 4.863756, 
    4.864096, 4.866197, 4.869948, 4.875145, 4.881518, 4.888731, 4.896425, 
    4.904231,
  // totalHeight(23,0, 0-49)
    4.895426, 4.901486, 4.90759, 4.913628, 4.919533, 4.92527, 4.930825, 
    4.936199, 4.941404, 4.946454, 4.951359, 4.956124, 4.960742, 4.965197, 
    4.969453, 4.973246, 4.977482, 4.980842, 4.983828, 4.986425, 4.988595, 
    4.990544, 4.991959, 4.992893, 4.993297, 4.993151, 4.992422, 4.991085, 
    4.989092, 4.986431, 4.982956, 4.978846, 4.973688, 4.967337, 4.959653, 
    4.950525, 4.939891, 4.927777, 4.914315, 4.899775, 4.884562, 4.869212, 
    4.85435, 4.840641, 4.828725, 4.819151, 4.812321, 4.808452, 4.807563, 
    4.809484,
  // totalHeight(23,1, 0-49)
    4.896116, 4.90232, 4.908538, 4.914664, 4.920634, 4.92641, 4.931978, 
    4.937342, 4.942514, 4.947505, 4.952327, 4.956984, 4.961471, 4.965774, 
    4.969862, 4.97324, 4.977746, 4.980855, 4.983581, 4.985966, 4.987989, 
    4.990112, 4.991745, 4.993001, 4.993792, 4.994096, 4.993859, 4.993059, 
    4.991638, 4.989619, 4.986797, 4.983615, 4.979371, 4.973888, 4.966999, 
    4.958545, 4.948429, 4.936629, 4.923249, 4.908527, 4.892865, 4.876808, 
    4.861016, 4.846209, 4.8331, 4.822316, 4.814339, 4.809461, 4.807758, 
    4.809104,
  // totalHeight(23,2, 0-49)
    4.896848, 4.903163, 4.909467, 4.915654, 4.921661, 4.927448, 4.933006, 
    4.938334, 4.943444, 4.948349, 4.953061, 4.957585, 4.961919, 4.966052, 
    4.96996, 4.972911, 4.977615, 4.980476, 4.982946, 4.985118, 4.986993, 
    4.989272, 4.991097, 4.992633, 4.993772, 4.994483, 4.9947, 4.994403, 
    4.993524, 4.99211, 4.989905, 4.987619, 4.98428, 4.979692, 4.973659, 
    4.965992, 4.956553, 4.945277, 4.932223, 4.917595, 4.901763, 4.885261, 
    4.868759, 4.853016, 4.838797, 4.826807, 4.81761, 4.81158, 4.808866, 
    4.809398,
  // totalHeight(23,3, 0-49)
    4.897707, 4.904102, 4.910461, 4.91668, 4.922695, 4.928468, 4.933987, 
    4.939251, 4.944274, 4.949068, 4.953646, 4.958017, 4.962181, 4.966132, 
    4.969855, 4.972373, 4.977182, 4.979805, 4.98203, 4.983992, 4.985715, 
    4.988125, 4.990106, 4.991872, 4.993307, 4.994374, 4.994997, 4.99516, 
    4.994784, 4.993926, 4.992285, 4.990835, 4.988363, 4.984661, 4.979513, 
    4.972706, 4.964067, 4.953493, 4.940991, 4.926718, 4.910996, 4.894328, 
    4.877372, 4.860893, 4.845701, 4.832562, 4.822122, 4.814842, 4.810956, 
    4.810467,
  // totalHeight(23,4, 0-49)
    4.898767, 4.905207, 4.911588, 4.917809, 4.923801, 4.929531, 4.934984, 
    4.940162, 4.945074, 4.949735, 4.954161, 4.958361, 4.962342, 4.966105, 
    4.969644, 4.971735, 4.976532, 4.978934, 4.980926, 4.982686, 4.984258, 
    4.986763, 4.988861, 4.990802, 4.992469, 4.993831, 4.994809, 4.995383, 
    4.99547, 4.995112, 4.993973, 4.993282, 4.991616, 4.988761, 4.984494, 
    4.978585, 4.970834, 4.9611, 4.949344, 4.935659, 4.920317, 4.903763, 
    4.886617, 4.869635, 4.853644, 4.839461, 4.827805, 4.819223, 4.814049, 
    4.812364,
  // totalHeight(23,5, 0-49)
    4.900073, 4.906525, 4.912896, 4.919085, 4.925028, 4.930689, 4.93605, 
    4.941118, 4.945899, 4.950413, 4.95467, 4.958691, 4.962481, 4.966052, 
    4.969409, 4.971094, 4.975749, 4.977942, 4.979719, 4.981287, 4.982709, 
    4.985273, 4.987438, 4.989486, 4.991323, 4.992917, 4.994195, 4.995135, 
    4.995642, 4.995732, 4.995035, 4.995014, 4.994076, 4.992012, 4.988597, 
    4.983593, 4.976781, 4.967987, 4.957124, 4.94423, 4.929503, 4.913324, 
    4.896254, 4.879013, 4.862425, 4.847337, 4.834532, 4.824646, 4.818106, 
    4.815096,
  // totalHeight(23,6, 0-49)
    4.901654, 4.908082, 4.914409, 4.920537, 4.926403, 4.931969, 4.937221, 
    4.94216, 4.946796, 4.951147, 4.95523, 4.959061, 4.962658, 4.966038, 
    4.969217, 4.970532, 4.974907, 4.976904, 4.978485, 4.979873, 4.981148, 
    4.983724, 4.985905, 4.987993, 4.989932, 4.991693, 4.993219, 4.994479, 
    4.995372, 4.995861, 4.995553, 4.996108, 4.995815, 4.994474, 4.991864, 
    4.987747, 4.98189, 4.974093, 4.964232, 4.952282, 4.938368, 4.922791, 
    4.906042, 4.888782, 4.87181, 4.855984, 4.842136, 4.830983, 4.823049, 
    4.818624,
  // totalHeight(23,7, 0-49)
    4.903516, 4.909886, 4.916139, 4.922179, 4.927942, 4.933392, 4.938515, 
    4.943311, 4.947791, 4.951973, 4.955874, 4.959517, 4.96292, 4.966109, 
    4.96911, 4.97011, 4.974067, 4.975875, 4.977278, 4.9785, 4.979634, 
    4.982173, 4.984315, 4.986372, 4.988348, 4.990219, 4.991941, 4.99348, 
    4.994731, 4.995581, 4.995622, 4.996662, 4.996929, 4.996234, 4.994371, 
    4.991102, 4.986189, 4.979417, 4.970619, 4.959719, 4.946767, 4.931982, 
    4.915766, 4.898709, 4.881564, 4.86518, 4.85042, 4.838073, 4.82876, 4.82288,
  // totalHeight(23,8, 0-49)
    4.905653, 4.911932, 4.918082, 4.924006, 4.929646, 4.934963, 4.939943, 
    4.944586, 4.948904, 4.952912, 4.956631, 4.960085, 4.963297, 4.966295, 
    4.969112, 4.969871, 4.973276, 4.974898, 4.97614, 4.977212, 4.978214, 
    4.980665, 4.982713, 4.984673, 4.986623, 4.988544, 4.990419, 4.992204, 
    4.99379, 4.994974, 4.995334, 4.996774, 4.997522, 4.997402, 4.996218, 
    4.993746, 4.989747, 4.98399, 4.976279, 4.966488, 4.954601, 4.940746, 
    4.925236, 4.908576, 4.891455, 4.874695, 4.859173, 4.845736, 4.835096, 
    4.827761,
  // totalHeight(23,9, 0-49)
    4.908045, 4.914205, 4.920225, 4.926012, 4.931508, 4.936678, 4.941504, 
    4.945988, 4.95014, 4.953975, 4.957514, 4.960781, 4.963801, 4.966605, 
    4.969224, 4.969835, 4.972563, 4.973999, 4.975098, 4.976038, 4.976922, 
    4.979229, 4.981129, 4.982932, 4.984797, 4.986721, 4.988709, 4.99071, 
    4.992615, 4.994116, 4.994787, 4.996551, 4.997704, 4.998085, 4.997517, 
    4.995781, 4.992645, 4.987872, 4.981241, 4.972581, 4.961812, 4.948979, 
    4.934303, 4.918199, 4.901276, 4.884313, 4.868188, 4.853786, 4.841904, 
    4.833155,
  // totalHeight(23,10, 0-49)
    4.910669, 4.916684, 4.922551, 4.928182, 4.93352, 4.938529, 4.943195, 
    4.947515, 4.951498, 4.955161, 4.958521, 4.961602, 4.96443, 4.967033, 
    4.969435, 4.969999, 4.971944, 4.973189, 4.97416, 4.974993, 4.975775, 
    4.977887, 4.979592, 4.981181, 4.982915, 4.984797, 4.986864, 4.989058, 
    4.991269, 4.993081, 4.994066, 4.996086, 4.997576, 4.998394, 4.998374, 
    4.997312, 4.994981, 4.991141, 4.985553, 4.978009, 4.968371, 4.956611, 
    4.942855, 4.927424, 4.910847, 4.893844, 4.877275, 4.862051, 4.849038, 
    4.838949,
  // totalHeight(23,11, 0-49)
    4.9135, 4.919349, 4.925044, 4.930502, 4.935669, 4.94051, 4.945008, 
    4.94916, 4.952974, 4.956462, 4.959645, 4.96254, 4.965172, 4.967559, 
    4.969719, 4.970341, 4.971409, 4.972464, 4.973328, 4.974075, 4.974782, 
    4.976649, 4.978117, 4.979452, 4.981015, 4.982821, 4.984939, 4.9873, 
    4.989808, 4.991928, 4.993247, 4.995461, 4.997231, 4.998425, 4.998889, 
    4.998437, 4.996847, 4.993878, 4.989277, 4.98281, 4.974285, 4.963607, 
    4.950817, 4.936144, 4.92003, 4.903127, 4.886267, 4.870369, 4.856357, 
    4.845033,
  // totalHeight(23,12, 0-49)
    4.916521, 4.922186, 4.927694, 4.932967, 4.937951, 4.942612, 4.946934, 
    4.950913, 4.954554, 4.957866, 4.960867, 4.963572, 4.965996, 4.968154, 
    4.970044, 4.970819, 4.970935, 4.971805, 4.972583, 4.973278, 4.97394, 
    4.975521, 4.976722, 4.97777, 4.979136, 4.98084, 4.982984, 4.985491, 
    4.988282, 4.990713, 4.99239, 4.994746, 4.996741, 4.998255, 4.999147, 
    4.999241, 4.998323, 4.996156, 4.992476, 4.987025, 4.97957, 4.969954, 
    4.958146, 4.944283, 4.928721, 4.912042, 4.895033, 4.878615, 4.863748, 
    4.851315,
  // totalHeight(23,13, 0-49)
    4.919718, 4.925189, 4.930497, 4.935571, 4.940359, 4.944829, 4.948966, 
    4.952762, 4.956221, 4.95935, 4.962162, 4.964666, 4.966873, 4.968783, 
    4.970378, 4.971375, 4.97047, 4.971176, 4.971901, 4.972583, 4.97324, 
    4.9745, 4.975414, 4.976161, 4.977314, 4.978903, 4.981051, 4.983681, 
    4.98674, 4.989478, 4.991546, 4.993996, 4.996167, 4.997951, 4.999214, 
    4.999793, 4.999481, 4.998042, 4.995209, 4.990702, 4.984257, 4.975666, 
    4.964827, 4.951798, 4.936854, 4.920501, 4.903476, 4.886686, 4.871117, 
    4.857717,
  // totalHeight(23,14, 0-49)
    4.92309, 4.928356, 4.933453, 4.938313, 4.942891, 4.947155, 4.95109, 
    4.954689, 4.957953, 4.960886, 4.963496, 4.96579, 4.967766, 4.969412, 
    4.970696, 4.97194, 4.96995, 4.970529, 4.971247, 4.971963, 4.972665, 
    4.973577, 4.974202, 4.97465, 4.975592, 4.977057, 4.979191, 4.981923, 
    4.985222, 4.988264, 4.990751, 4.99325, 4.995551, 4.997555, 4.999138, 
    5.000143, 5.000372, 4.999589, 4.997525, 4.993887, 4.988383, 4.980763, 
    4.970865, 4.958676, 4.944394, 4.928452, 4.91153, 4.894514, 4.878398, 
    4.864184,
  // totalHeight(23,15, 0-49)
    4.926639, 4.931692, 4.936564, 4.941194, 4.945542, 4.949579, 4.95329, 
    4.956672, 4.959722, 4.962442, 4.964838, 4.966904, 4.968638, 4.970015, 
    4.970989, 4.972441, 4.969296, 4.969801, 4.970569, 4.97138, 4.972188, 
    4.972746, 4.973093, 4.973263, 4.974007, 4.975351, 4.977458, 4.980263, 
    4.983772, 4.9871, 4.99003, 4.992534, 4.99492, 4.997099, 4.99895, 
    5.000324, 5.001028, 5.000831, 4.999461, 4.996616, 4.99198, 4.985271, 
    4.976275, 4.96492, 4.95133, 4.93587, 4.919161, 4.902054, 4.885547, 
    4.870674,
  // totalHeight(23,16, 0-49)
    4.93037, 4.935199, 4.939828, 4.944206, 4.948298, 4.952079, 4.95554, 
    4.958678, 4.961491, 4.96398, 4.966144, 4.967977, 4.969463, 4.970573, 
    4.971258, 4.972813, 4.968417, 4.968924, 4.969812, 4.970793, 4.971777, 
    4.971989, 4.972089, 4.97202, 4.972597, 4.973833, 4.975907, 4.978754, 
    4.982432, 4.986019, 4.989403, 4.991866, 4.994292, 4.996596, 4.998665, 
    5.000351, 5.00147, 5.001792, 5.001044, 4.998916, 4.995078, 4.989218, 
    4.981081, 4.970545, 4.957668, 4.942747, 4.926349, 4.909281, 4.892532, 
    4.877156,
  // totalHeight(23,17, 0-49)
    4.934283, 4.938868, 4.943231, 4.947325, 4.951125, 4.954617, 4.957797, 
    4.960662, 4.963215, 4.965456, 4.967381, 4.968978, 4.970225, 4.971089, 
    4.971526, 4.973015, 4.967241, 4.967832, 4.968923, 4.970154, 4.971397, 
    4.971285, 4.971189, 4.970938, 4.971395, 4.972552, 4.974586, 4.97745, 
    4.981249, 4.985054, 4.988883, 4.991256, 4.99367, 4.99605, 4.998283, 
    5.000228, 5.001703, 5.002481, 5.002286, 5.000806, 4.997698, 4.992626, 
    4.985308, 4.975571, 4.96342, 4.94909, 4.933088, 4.91618, 4.89933, 4.883603,
  // totalHeight(23,18, 0-49)
    4.938361, 4.942673, 4.946726, 4.950492, 4.953959, 4.957124, 4.95999, 
    4.962561, 4.964844, 4.966834, 4.968524, 4.969899, 4.970932, 4.971589, 
    4.971833, 4.973045, 4.96572, 4.966478, 4.967849, 4.969416, 4.971005, 
    4.970614, 4.970387, 4.970029, 4.97043, 4.971549, 4.973553, 4.976407, 
    4.980273, 4.98424, 4.988482, 4.990712, 4.993061, 4.995459, 4.9978, 
    4.999946, 5.001716, 5.002888, 5.003185, 5.00229, 4.99985, 4.995514, 
    4.988973, 4.980016, 4.968597, 4.9549, 4.939373, 4.922735, 4.905919, 
    4.889985,
  // totalHeight(23,19, 0-49)
    4.942561, 4.94654, 4.950226, 4.953609, 4.956694, 4.959494, 4.962023, 
    4.964293, 4.96631, 4.96807, 4.969558, 4.970748, 4.971611, 4.972114, 
    4.972234, 4.972956, 4.963853, 4.964847, 4.966568, 4.968548, 4.970571, 
    4.969965, 4.969689, 4.969313, 4.969736, 4.970868, 4.972862, 4.97569, 
    4.979569, 4.98363, 4.988221, 4.990247, 4.992464, 4.994816, 4.9972, 
    4.999482, 5.001488, 5.002994, 5.003723, 5.003355, 5.001528, 4.99788, 
    4.992079, 4.983882, 4.973204, 4.960176, 4.945191, 4.928922, 4.912266, 
    4.896266,
  // totalHeight(23,20, 0-49)
    4.947812, 4.952392, 4.956592, 4.960402, 4.963821, 4.966853, 4.969504, 
    4.971782, 4.973697, 4.975266, 4.976511, 4.977463, 4.978164, 4.978666, 
    4.97904, 30, 4.962282, 4.963513, 4.965213, 4.966989, 4.9687, 4.967034, 
    4.965853, 4.964697, 4.964581, 4.965442, 4.967443, 4.970533, 4.974926, 
    4.979701, 4.98531, 4.987769, 4.990425, 4.993213, 4.996024, 4.998729, 
    5.001162, 5.003111, 5.004313, 5.004456, 5.003191, 5.000156, 4.995014, 
    4.987504, 4.977509, 4.965121, 4.950686, 4.934827, 4.918398, 4.902422,
  // totalHeight(23,21, 0-49)
    4.952321, 4.956649, 4.960524, 4.963956, 4.966967, 4.969578, 4.971817, 
    4.973706, 4.975272, 4.97654, 4.977539, 4.978305, 4.978885, 4.979341, 
    4.979759, 30, 4.957336, 4.958926, 4.96105, 4.963284, 4.965437, 4.96349, 
    4.962173, 4.960936, 4.960859, 4.961868, 4.964108, 4.967514, 4.972302, 
    4.977538, 4.983817, 4.986392, 4.989252, 4.992331, 4.995506, 4.998638, 
    5.001549, 5.004018, 5.005775, 5.006501, 5.005841, 5.003427, 4.99891, 
    4.992016, 4.982603, 4.970729, 4.956704, 4.941106, 4.924758, 4.90866,
  // totalHeight(23,22, 0-49)
    4.956862, 4.960968, 4.964542, 4.967612, 4.970216, 4.972399, 4.974205, 
    4.975675, 4.97685, 4.977767, 4.978467, 4.978996, 4.979407, 4.979776, 
    4.98021, 30, 4.953183, 4.955079, 4.957577, 4.960221, 4.962775, 4.960561, 
    4.959106, 4.957771, 4.957701, 4.958802, 4.961205, 4.96483, 4.969896, 
    4.975457, 4.982234, 4.984813, 4.987763, 4.991016, 4.994449, 4.997913, 
    5.001224, 5.004153, 5.00642, 5.0077, 5.007632, 5.005837, 5.001956, 
    4.995699, 4.986902, 4.975594, 4.962046, 4.946799, 4.930641, 4.914544,
  // totalHeight(23,23, 0-49)
    4.961319, 4.96523, 4.968522, 4.971242, 4.973449, 4.975204, 4.976571, 
    4.977608, 4.978371, 4.97891, 4.979281, 4.979536, 4.979744, 4.979992, 
    4.980406, 30, 4.949828, 4.951932, 4.954688, 4.957613, 4.960438, 4.957965, 
    4.956351, 4.954892, 4.954782, 4.955913, 4.958411, 4.962177, 4.967437, 
    4.973226, 4.980362, 4.982919, 4.985924, 4.989314, 4.992963, 4.996723, 
    5.000404, 5.00377, 5.006535, 5.008361, 5.008878, 5.007699, 5.004451, 
    4.998827, 4.990645, 4.979904, 4.966846, 4.951975, 4.936047, 4.920007,
  // totalHeight(23,24, 0-49)
    4.965569, 4.969304, 4.972334, 4.974724, 4.976551, 4.977893, 4.978831, 
    4.979438, 4.979786, 4.97994, 4.979965, 4.979927, 4.979905, 4.98, 4.98035, 
    30, 4.947584, 4.949786, 4.952665, 4.955732, 4.958699, 4.956051, 4.954333, 
    4.952793, 4.952653, 4.953795, 4.956342, 4.960189, 4.965566, 4.971498, 
    4.97887, 4.981437, 4.984508, 4.988023, 4.991858, 4.995862, 4.999844, 
    5.003561, 5.006723, 5.008988, 5.009978, 5.009296, 5.006564, 5.001464, 
    4.993795, 4.983542, 4.970922, 4.956411, 4.940742, 4.924834,
  // totalHeight(23,25, 0-49)
    4.969476, 4.973059, 4.975853, 4.977944, 4.97942, 4.980377, 4.980908, 
    4.981107, 4.981056, 4.98083, 4.980508, 4.980166, 4.979897, 4.979808, 
    4.980052, 30, 4.946215, 4.948393, 4.951257, 4.954316, 4.95728, 4.954575, 
    4.95283, 4.951283, 4.951154, 4.952318, 4.9549, 4.958794, 4.96423, 
    4.970243, 4.97773, 4.980377, 4.983562, 4.987227, 4.991247, 4.995472, 
    4.999707, 5.003707, 5.007178, 5.009773, 5.011113, 5.010795, 5.008437, 
    5.003716, 4.996426, 4.986541, 4.974265, 4.960062, 4.944643, 4.928911,
  // totalHeight(23,26, 0-49)
    4.972922, 4.976376, 4.97897, 4.980797, 4.981965, 4.982578, 4.982746, 
    4.982569, 4.982144, 4.981558, 4.980897, 4.980248, 4.979712, 4.979408, 
    4.979493, 30, 4.945743, 4.947777, 4.950482, 4.953379, 4.956195, 4.95355, 
    4.951866, 4.950394, 4.950324, 4.951531, 4.954144, 4.95806, 4.963513, 
    4.969546, 4.977036, 4.979848, 4.983212, 4.987065, 4.991282, 4.995709, 
    5.000151, 5.00436, 5.008039, 5.010841, 5.012385, 5.012269, 5.010112, 
    5.005596, 4.998515, 4.988846, 4.976793, 4.962817, 4.947624, 4.932106,
  // totalHeight(23,27, 0-49)
    4.975794, 4.979151, 4.981586, 4.983203, 4.984118, 4.984444, 4.9843, 
    4.983793, 4.983029, 4.982104, 4.981112, 4.980152, 4.979331, 4.978775, 
    4.978641, 30, 4.946302, 4.948066, 4.950467, 4.953045, 4.955564, 4.953069, 
    4.9515, 4.950153, 4.950165, 4.951417, 4.954041, 4.957945, 4.963362, 
    4.969354, 4.976735, 4.979789, 4.983385, 4.987454, 4.991872, 4.996479, 
    5.001076, 5.005418, 5.009205, 5.012092, 5.013698, 5.013628, 5.011506, 
    5.007021, 4.999983, 4.990378, 4.978427, 4.964598, 4.9496, 4.934321,
  // totalHeight(23,28, 0-49)
    4.978009, 4.981311, 4.983644, 4.985114, 4.985842, 4.985948, 4.985551, 
    4.984766, 4.983699, 4.982455, 4.981137, 4.979851, 4.978716, 4.977863, 
    4.977447, 30, 4.948286, 4.949656, 4.951609, 4.953715, 4.955791, 4.953478, 
    4.952028, 4.950802, 4.950869, 4.952122, 4.9547, 4.958529, 4.963839, 
    4.969721, 4.97689, 4.98023, 4.984081, 4.988367, 4.992958, 4.997692, 
    5.002371, 5.006748, 5.010526, 5.01336, 5.014878, 5.014691, 5.012437, 
    5.007819, 5.000664, 4.990985, 4.979025, 4.965273, 4.950454, 4.935455,
  // totalHeight(23,29, 0-49)
    4.979519, 4.98282, 4.985117, 4.98652, 4.987142, 4.987102, 4.986516, 
    4.985497, 4.984156, 4.982601, 4.980945, 4.979306, 4.977814, 4.976609, 
    4.975844, 30, 4.951502, 4.952365, 4.95373, 4.955213, 4.956685, 4.954491, 
    4.953069, 4.951875, 4.951902, 4.953065, 4.955513, 4.959191, 4.964319, 
    4.970014, 4.976858, 4.980478, 4.984567, 4.989044, 4.993778, 4.998605, 
    5.003326, 5.007692, 5.011411, 5.01414, 5.015511, 5.015141, 5.012679, 
    5.007847, 5.000496, 4.990666, 4.978632, 4.964911, 4.95025, 4.93554,
  // totalHeight(23,30, 0-49)
    4.979384, 4.981814, 4.983278, 4.983901, 4.98382, 4.983175, 4.9821, 
    4.980711, 4.979107, 4.977366, 4.975537, 4.973642, 4.971686, 4.969653, 
    4.967526, 4.968501, 4.95388, 4.953983, 4.955086, 4.956669, 4.958492, 
    4.957497, 4.95718, 4.956963, 4.957675, 4.959179, 4.961603, 4.964932, 
    4.969421, 4.974288, 4.980054, 4.983217, 4.986848, 4.990884, 4.995209, 
    4.999662, 5.004045, 5.008105, 5.011535, 5.013987, 5.015082, 5.014435, 
    5.011695, 5.006598, 4.999016, 4.98902, 4.976917, 4.96326, 4.948817, 
    4.934488,
  // totalHeight(23,31, 0-49)
    4.979453, 4.981999, 4.983564, 4.984265, 4.984229, 4.983586, 4.982464, 
    4.980983, 4.979244, 4.977332, 4.97531, 4.973215, 4.971061, 4.968839, 
    4.966521, 4.968116, 4.955175, 4.954739, 4.955228, 4.956167, 4.957366, 
    4.956451, 4.956088, 4.955835, 4.956506, 4.958014, 4.960509, 4.963962, 
    4.96857, 4.97352, 4.979156, 4.9828, 4.986884, 4.991324, 4.995992, 
    5.000715, 5.005282, 5.009428, 5.012842, 5.01517, 5.016033, 5.015054, 
    5.011901, 5.006335, 4.99827, 4.987822, 4.975352, 4.961461, 4.94695, 
    4.932743,
  // totalHeight(23,32, 0-49)
    4.978727, 4.981336, 4.98298, 4.983766, 4.983811, 4.983236, 4.982162, 
    4.980702, 4.978957, 4.977013, 4.974936, 4.972773, 4.970546, 4.968249, 
    4.965855, 4.967472, 4.956299, 4.9554, 4.955333, 4.955686, 4.956318, 
    4.955542, 4.955204, 4.95499, 4.955684, 4.95724, 4.959817, 4.963375, 
    4.968049, 4.97302, 4.978463, 4.982544, 4.987028, 4.991814, 4.996756, 
    5.001674, 5.006341, 5.010485, 5.013781, 5.015877, 5.016394, 5.014968, 
    5.011288, 5.00515, 4.996514, 4.985552, 4.97268, 4.958555, 4.944016, 
    4.929998,
  // totalHeight(23,33, 0-49)
    4.977302, 4.979942, 4.981656, 4.982538, 4.982697, 4.982244, 4.981289, 
    4.979935, 4.97828, 4.976404, 4.974379, 4.972252, 4.970052, 4.967782, 
    4.965415, 4.966619, 4.957237, 4.955972, 4.955427, 4.955264, 4.955398, 
    4.954807, 4.954551, 4.954451, 4.955221, 4.956857, 4.959517, 4.963147, 
    4.967824, 4.972751, 4.977959, 4.982429, 4.987256, 4.992321, 4.997468, 
    5.002501, 5.007183, 5.011227, 5.014306, 5.01606, 5.016119, 5.014136, 
    5.009826, 5.003026, 4.99375, 4.982231, 4.968952, 4.954619, 4.940107, 
    4.926363,
  // totalHeight(23,34, 0-49)
    4.975289, 4.977936, 4.979716, 4.98071, 4.981011, 4.98072, 4.979937, 
    4.978752, 4.977258, 4.975528, 4.97363, 4.971616, 4.969521, 4.967354, 
    4.965097, 4.965625, 4.958004, 4.956473, 4.955529, 4.954925, 4.954628, 
    4.954253, 4.954134, 4.954203, 4.955094, 4.956829, 4.959558, 4.963218, 
    4.967833, 4.972657, 4.977599, 4.982405, 4.987512, 4.992789, 4.998067, 
    5.003136, 5.007743, 5.011593, 5.01435, 5.015658, 5.015156, 5.012516, 
    5.007489, 4.99996, 4.990002, 4.977917, 4.964249, 4.94976, 4.935356, 
    4.921988,
  // totalHeight(23,35, 0-49)
    4.972805, 4.975446, 4.977287, 4.978399, 4.978864, 4.978765, 4.978192, 
    4.977223, 4.97594, 4.97441, 4.972696, 4.970852, 4.968914, 4.966905, 
    4.964818, 4.964561, 4.958642, 4.956938, 4.955672, 4.954696, 4.954036, 
    4.953892, 4.953948, 4.954236, 4.955279, 4.957119, 4.959894, 4.963537, 
    4.96802, 4.972685, 4.977338, 4.982416, 4.987737, 4.993151, 4.998478, 
    5.003494, 5.007935, 5.011493, 5.013832, 5.014596, 5.013438, 5.010059, 
    5.004251, 4.995952, 4.985302, 4.972674, 4.958676, 4.944117, 4.929926, 
    4.917049,
  // totalHeight(23,36, 0-49)
    4.969972, 4.972589, 4.974487, 4.975722, 4.97636, 4.976475, 4.976136, 
    4.975414, 4.974378, 4.973086, 4.971597, 4.969959, 4.968216, 4.966397, 
    4.964516, 4.963494, 4.959198, 4.957397, 4.955878, 4.954597, 4.953636, 
    4.953732, 4.95399, 4.954529, 4.955745, 4.957692, 4.960482, 4.964052, 
    4.968329, 4.972781, 4.977126, 4.9824, 4.987854, 4.993322, 4.99861, 
    5.00348, 5.007657, 5.010827, 5.01265, 5.01278, 5.01089, 5.006711, 
    5.000083, 4.991011, 4.979698, 4.966591, 4.952356, 4.937846, 4.924, 
    4.911744,
  // totalHeight(23,37, 0-49)
    4.966919, 4.969494, 4.971436, 4.972788, 4.973604, 4.973938, 4.973849, 
    4.973393, 4.972626, 4.971597, 4.970358, 4.968953, 4.967428, 4.965818, 
    4.964155, 4.96248, 4.959714, 4.957877, 4.956165, 4.954644, 4.953441, 
    4.953775, 4.954249, 4.955064, 4.95646, 4.9585, 4.961268, 4.964707, 
    4.968708, 4.972888, 4.976903, 4.982288, 4.987783, 4.99321, 4.998359, 
    5.002985, 5.006799, 5.009483, 5.010701, 5.010118, 5.007432, 5.002418, 
    4.994967, 4.985151, 4.973249, 4.959768, 4.945435, 4.931123, 4.917774, 
    4.906282,
  // totalHeight(23,38, 0-49)
    4.963768, 4.966279, 4.968248, 4.969707, 4.970693, 4.971244, 4.971407, 
    4.971223, 4.970736, 4.969985, 4.969013, 4.967857, 4.966562, 4.96517, 
    4.963725, 4.96156, 4.96023, 4.958398, 4.956545, 4.954842, 4.953458, 
    4.95402, 4.954714, 4.955815, 4.95739, 4.959505, 4.962207, 4.965453, 
    4.969102, 4.972951, 4.976608, 4.982003, 4.987434, 4.992712, 4.997617, 
    5.001892, 5.005239, 5.007343, 5.007872, 5.006511, 5.002993, 4.997136, 
    4.988894, 4.978408, 4.96603, 4.952328, 4.938067, 4.924137, 4.911459, 
    4.90088,
  // totalHeight(23,39, 0-49)
    4.960637, 4.963058, 4.965035, 4.96658, 4.967719, 4.968476, 4.968884, 
    4.968968, 4.968763, 4.968296, 4.967598, 4.966702, 4.965645, 4.964471, 
    4.963233, 4.960762, 4.96077, 4.958971, 4.957023, 4.955193, 4.953681, 
    4.954453, 4.955369, 4.956755, 4.958495, 4.960657, 4.963246, 4.966229, 
    4.969455, 4.972909, 4.976169, 4.981458, 4.986709, 4.99172, 4.996265, 
    5.000077, 5.002857, 5.00429, 5.004058, 5.001873, 4.997508, 4.990834, 
    4.981874, 4.970839, 4.958142, 4.944409, 4.930429, 4.917086, 4.905265, 
    4.895751,
  // totalHeight(23,40, 0-49)
    4.95763, 4.959937, 4.961891, 4.963499, 4.964767, 4.965711, 4.966346, 
    4.966689, 4.966758, 4.96657, 4.966147, 4.965512, 4.964697, 4.963742, 
    4.962697, 4.960098, 4.961344, 4.959596, 4.957597, 4.95569, 4.954103, 
    4.95507, 4.956193, 4.957851, 4.959733, 4.961905, 4.964325, 4.966981, 
    4.969707, 4.972701, 4.975508, 4.980567, 4.98551, 4.990129, 4.99419, 
    4.997423, 4.999531, 5.000209, 4.99916, 4.996129, 4.990932, 4.983507, 
    4.973942, 4.962516, 4.949704, 4.936168, 4.922704, 4.910172, 4.8994, 
    4.891098,
  // totalHeight(23,41, 0-49)
    4.95484, 4.957002, 4.958905, 4.960543, 4.961915, 4.963018, 4.963856, 
    4.964436, 4.964763, 4.964844, 4.96469, 4.964315, 4.963742, 4.963002, 
    4.962139, 4.959574, 4.961953, 4.96027, 4.958256, 4.956322, 4.954705, 
    4.955848, 4.957162, 4.959065, 4.961057, 4.963192, 4.965388, 4.967646, 
    4.9698, 4.972257, 4.974547, 4.979238, 4.983736, 4.987826, 4.991275, 
    4.993814, 4.995153, 4.995003, 4.993098, 4.989223, 4.983247, 4.975173, 
    4.965159, 4.953546, 4.940858, 4.927775, 4.915082, 4.903592, 4.89406, 
    4.887104,
  // totalHeight(23,42, 0-49)
    4.952335, 4.954322, 4.956143, 4.957779, 4.959219, 4.960448, 4.961461, 
    4.962251, 4.962814, 4.963148, 4.963252, 4.963131, 4.962798, 4.962269, 
    4.961581, 4.959179, 4.962581, 4.960975, 4.958985, 4.95707, 4.955463, 
    4.956761, 4.958241, 4.960354, 4.962413, 4.964461, 4.966369, 4.96816, 
    4.96967, 4.971512, 4.973205, 4.977383, 4.981291, 4.984713, 4.987421, 
    4.989151, 4.989631, 4.988597, 4.985819, 4.981133, 4.974466, 4.965889, 
    4.955624, 4.944065, 4.931768, 4.919414, 4.907753, 4.897533, 4.889417, 
    4.883925,
  // totalHeight(23,43, 0-49)
    4.950162, 4.951948, 4.953654, 4.955253, 4.956722, 4.958042, 4.959195, 
    4.960165, 4.960937, 4.9615, 4.961845, 4.961969, 4.961868, 4.961549, 
    4.961031, 4.958889, 4.963201, 4.961686, 4.959754, 4.957897, 4.956337, 
    4.957767, 4.959386, 4.961664, 4.963741, 4.965644, 4.967198, 4.968454, 
    4.96925, 4.970394, 4.971401, 4.97492, 4.97809, 4.980704, 4.982542, 
    4.983356, 4.982902, 4.980946, 4.977309, 4.971876, 4.964646, 4.955748, 
    4.945463, 4.934228, 4.922611, 4.91127, 4.900899, 4.892162, 4.885618, 
    4.881681,
  // totalHeight(23,44, 0-49)
    4.948341, 4.9499, 4.951458, 4.952984, 4.954449, 4.955821, 4.957075, 
    4.958187, 4.959137, 4.959904, 4.96047, 4.960821, 4.960945, 4.960835, 
    4.960487, 4.958665, 4.963771, 4.962362, 4.960526, 4.958759, 4.957273, 
    4.958815, 4.960539, 4.962932, 4.96497, 4.966668, 4.967808, 4.968459, 
    4.968475, 4.968838, 4.96906, 4.971774, 4.974064, 4.975734, 4.976582, 
    4.976389, 4.974941, 4.972054, 4.967598, 4.961523, 4.953889, 4.944887, 
    4.934844, 4.92422, 4.913573, 4.903521, 4.894681, 4.887616, 4.882772, 
    4.88045,
  // totalHeight(23,45, 0-49)
    4.946861, 4.948171, 4.949554, 4.950976, 4.952395, 4.95378, 4.955097, 
    4.956316, 4.957407, 4.958346, 4.959108, 4.95967, 4.960007, 4.960099, 
    4.959925, 4.958453, 4.964239, 4.962955, 4.961242, 4.959595, 4.958201, 
    4.959833, 4.961634, 4.964084, 4.966026, 4.967455, 4.968119, 4.968105, 
    4.967281, 4.966781, 4.966122, 4.967893, 4.969166, 4.96977, 4.969526, 
    4.968252, 4.96578, 4.961977, 4.956776, 4.950191, 4.942346, 4.933481, 
    4.923957, 4.914234, 4.904842, 4.896333, 4.889235, 4.883993, 4.880938, 
    4.880261,
  // totalHeight(23,46, 0-49)
    4.945683, 4.946728, 4.947913, 4.949197, 4.950539, 4.951898, 4.953238, 
    4.954524, 4.955721, 4.9568, 4.957727, 4.958476, 4.959012, 4.959301, 
    4.959304, 4.958188, 4.964537, 4.963399, 4.961836, 4.96033, 4.959041, 
    4.960747, 4.962584, 4.965035, 4.966822, 4.967922, 4.968055, 4.967322, 
    4.965609, 4.964171, 4.962538, 4.963241, 4.963384, 4.962819, 4.961406, 
    4.959006, 4.955505, 4.950835, 4.944994, 4.938061, 4.930218, 4.921744, 
    4.913013, 4.904469, 4.896591, 4.889844, 4.884655, 4.881347, 4.88013, 
    4.881088,
  // totalHeight(23,47, 0-49)
    4.944736, 4.945503, 4.946472, 4.947594, 4.948827, 4.950127, 4.951453, 
    4.952766, 4.954033, 4.955215, 4.956281, 4.957191, 4.957909, 4.958385, 
    4.958569, 4.957788, 4.964588, 4.96362, 4.962227, 4.960876, 4.959701, 
    4.961462, 4.963302, 4.965695, 4.96727, 4.967989, 4.967543, 4.96605, 
    4.96341, 4.960971, 4.958283, 4.957822, 4.956746, 4.954939, 4.952308, 
    4.948769, 4.944271, 4.938815, 4.932464, 4.925364, 4.917743, 4.909908, 
    4.902228, 4.895111, 4.888963, 4.884154, 4.880991, 4.879674, 4.8803, 
    4.882845,
  // totalHeight(23,48, 0-49)
    4.943918, 4.9444, 4.945139, 4.946082, 4.947184, 4.948393, 4.949674, 
    4.950984, 4.952284, 4.953536, 4.954707, 4.955752, 4.956629, 4.957283, 
    4.957647, 4.957171, 4.964309, 4.96353, 4.962326, 4.961139, 4.960081, 
    4.961879, 4.963689, 4.965969, 4.967283, 4.967573, 4.966515, 4.964235, 
    4.960649, 4.957168, 4.953364, 4.951672, 4.949322, 4.946239, 4.942382, 
    4.93773, 4.932302, 4.926166, 4.919459, 4.91238, 4.905197, 4.898226, 
    4.891818, 4.886326, 4.882068, 4.87931, 4.878233, 4.878918, 4.881347, 
    4.885399,
  // totalHeight(23,49, 0-49)
    4.943139, 4.943075, 4.943346, 4.94389, 4.944658, 4.945593, 4.946653, 
    4.94779, 4.948959, 4.950121, 4.951228, 4.952226, 4.953055, 4.953636, 
    4.953867, 4.95286, 4.96727, 4.965607, 4.963223, 4.960995, 4.959105, 
    4.962934, 4.966742, 4.971398, 4.97398, 4.974425, 4.972114, 4.967323, 
    4.959898, 4.952757, 4.94517, 4.942115, 4.938286, 4.93369, 4.928385, 
    4.922455, 4.916029, 4.909282, 4.902445, 4.895787, 4.889615, 4.884236, 
    4.879951, 4.877014, 4.875607, 4.87583, 4.877696, 4.881118, 4.885932, 
    4.8919,
  // totalHeight(24,0, 0-49)
    4.910848, 4.916671, 4.922301, 4.927701, 4.932858, 4.937772, 4.942453, 
    4.946915, 4.951171, 4.955228, 4.959091, 4.962752, 4.9662, 4.969418, 
    4.972382, 4.974842, 4.97764, 4.97967, 4.981387, 4.98284, 4.984052, 
    4.985279, 4.986291, 4.987188, 4.987974, 4.988667, 4.989259, 4.989744, 
    4.990077, 4.99023, 4.990046, 4.989658, 4.988633, 4.986763, 4.983824, 
    4.979576, 4.973786, 4.966261, 4.95687, 4.945582, 4.932493, 4.917852, 
    4.902067, 4.8857, 4.869432, 4.854009, 4.840175, 4.8286, 4.81981, 4.81415,
  // totalHeight(24,1, 0-49)
    4.911695, 4.917596, 4.923278, 4.928706, 4.933865, 4.938758, 4.943394, 
    4.94779, 4.951956, 4.955903, 4.959635, 4.963151, 4.96644, 4.969491, 
    4.972285, 4.974345, 4.977362, 4.979176, 4.980673, 4.981947, 4.983039, 
    4.984436, 4.985643, 4.986808, 4.987906, 4.988943, 4.989892, 4.990752, 
    4.991471, 4.992055, 4.9923, 4.992604, 4.992283, 4.991125, 4.988891, 
    4.985327, 4.980186, 4.973246, 4.964348, 4.95343, 4.940554, 4.92594, 
    4.909973, 4.89321, 4.876342, 4.860144, 4.845407, 4.832861, 4.823102, 
    4.816533,
  // totalHeight(24,2, 0-49)
    4.912669, 4.91862, 4.924327, 4.929756, 4.934893, 4.93974, 4.944309, 
    4.948617, 4.952674, 4.956494, 4.960084, 4.963445, 4.966572, 4.969456, 
    4.972089, 4.973764, 4.97696, 4.978581, 4.979879, 4.980993, 4.981977, 
    4.983537, 4.984918, 4.986313, 4.987674, 4.988997, 4.990244, 4.99141, 
    4.992443, 4.993364, 4.993931, 4.994814, 4.995092, 4.994552, 4.992957, 
    4.990049, 4.985571, 4.979286, 4.97101, 4.96065, 4.948229, 4.933926, 
    4.918087, 4.901238, 4.884052, 4.867312, 4.851837, 4.8384, 4.827665, 
    4.820106,
  // totalHeight(24,3, 0-49)
    4.91381, 4.919782, 4.925487, 4.93089, 4.935981, 4.940762, 4.945244, 
    4.949446, 4.953381, 4.957063, 4.960503, 4.963704, 4.966669, 4.969393, 
    4.971877, 4.973185, 4.976495, 4.977949, 4.979077, 4.98005, 4.980939, 
    4.982646, 4.984173, 4.98575, 4.987319, 4.988866, 4.990348, 4.991757, 
    4.993032, 4.994204, 4.994997, 4.996337, 4.997099, 4.997078, 4.996046, 
    4.993749, 4.98993, 4.984341, 4.976785, 4.967137, 4.955381, 4.941644, 
    4.92622, 4.909581, 4.892362, 4.875326, 4.859296, 4.845084, 4.833405, 
    4.824807,
  // totalHeight(24,4, 0-49)
    4.915136, 4.921102, 4.926778, 4.932133, 4.937155, 4.941853, 4.946233, 
    4.950315, 4.954117, 4.957655, 4.960942, 4.963984, 4.966791, 4.969364, 
    4.971712, 4.972683, 4.976027, 4.977337, 4.978322, 4.979175, 4.979979, 
    4.981809, 4.983449, 4.985155, 4.986871, 4.988581, 4.990238, 4.991829, 
    4.993289, 4.994633, 4.995562, 4.997245, 4.998381, 4.99878, 4.998229, 
    4.996487, 4.993301, 4.988431, 4.98166, 4.972841, 4.961918, 4.948961, 
    4.934201, 4.918041, 4.901056, 4.883966, 4.867583, 4.852731, 4.840173, 
    4.830526,
  // totalHeight(24,5, 0-49)
    4.916652, 4.922581, 4.928205, 4.933492, 4.938432, 4.943027, 4.947294, 
    4.951252, 4.954916, 4.958307, 4.961441, 4.964331, 4.966985, 4.969419, 
    4.971646, 4.972317, 4.975591, 4.976784, 4.977652, 4.978406, 4.979137, 
    4.981061, 4.982773, 4.984549, 4.986351, 4.988163, 4.989937, 4.99166, 
    4.993255, 4.994709, 4.995702, 4.997621, 4.999029, 4.999756, 4.999607, 
    4.99836, 4.995777, 4.99162, 4.985671, 4.977759, 4.967791, 4.95578, 
    4.941885, 4.926431, 4.909919, 4.893005, 4.876468, 4.861129, 4.847784, 
    4.837109,
  // totalHeight(24,6, 0-49)
    4.918346, 4.924214, 4.929765, 4.934965, 4.939806, 4.944293, 4.948441, 
    4.952268, 4.955794, 4.959041, 4.962029, 4.96477, 4.967284, 4.969589, 
    4.971706, 4.972129, 4.975222, 4.976313, 4.97709, 4.977765, 4.978433, 
    4.980412, 4.982152, 4.983939, 4.985767, 4.98762, 4.989464, 4.991274, 
    4.992972, 4.994491, 4.995498, 4.997561, 4.999152, 5.000124, 5.000306, 
    4.999494, 4.997471, 4.994012, 4.988893, 4.98193, 4.972991, 4.96204, 
    4.949162, 4.934595, 4.918754, 4.902222, 4.885718, 4.870051, 4.856028, 
    4.844377,
  // totalHeight(24,7, 0-49)
    4.920202, 4.925986, 4.931444, 4.936544, 4.941278, 4.945648, 4.949674, 
    4.953372, 4.956764, 4.959872, 4.962719, 4.965323, 4.967707, 4.969892, 
    4.971903, 4.972137, 4.97493, 4.975934, 4.976643, 4.977257, 4.977875, 
    4.979867, 4.981587, 4.983323, 4.985119, 4.986961, 4.988832, 4.990698, 
    4.992476, 4.994034, 4.995025, 4.997155, 4.998858, 5.000006, 5.000455, 
    5.000026, 4.99852, 4.995724, 4.991423, 4.985418, 4.977546, 4.96772, 
    4.955954, 4.942404, 4.92739, 4.911408, 4.89511, 4.879266, 4.864686, 
    4.852138,
  // totalHeight(24,8, 0-49)
    4.922203, 4.927882, 4.933229, 4.938216, 4.942835, 4.947088, 4.95099, 
    4.954564, 4.957827, 4.960806, 4.963521, 4.965996, 4.968257, 4.970326, 
    4.972233, 4.972349, 4.97472, 4.975642, 4.976302, 4.976875, 4.977454, 
    4.979413, 4.981066, 4.982692, 4.984403, 4.986189, 4.988052, 4.989952, 
    4.991802, 4.993388, 4.994358, 4.996493, 4.998249, 4.999518, 5.000184, 
    5.000089, 4.999055, 4.996887, 4.993373, 4.988306, 4.981501, 4.972822, 
    4.962221, 4.949767, 4.935689, 4.92039, 4.904442, 4.888564, 4.873551, 
    4.860202,
  // totalHeight(24,9, 0-49)
    4.924329, 4.929885, 4.935111, 4.939977, 4.944474, 4.948607, 4.95239, 
    4.955841, 4.958982, 4.961837, 4.964429, 4.966784, 4.968927, 4.970881, 
    4.972672, 4.972748, 4.974584, 4.975426, 4.976051, 4.9766, 4.977153, 
    4.97903, 4.980568, 4.982034, 4.983612, 4.985303, 4.987132, 4.989051, 
    4.990974, 4.992595, 4.993559, 4.995654, 4.997419, 4.998772, 4.999612, 
    4.999809, 4.999207, 4.997621, 4.994853, 4.990687, 4.98492, 4.977376, 
    4.967946, 4.956625, 4.943548, 4.929025, 4.913544, 4.897759, 4.88244, 
    4.868397,
  // totalHeight(24,10, 0-49)
    4.926576, 4.931991, 4.937082, 4.941818, 4.946189, 4.950202, 4.953865, 
    4.957198, 4.960221, 4.962958, 4.965433, 4.967671, 4.969696, 4.971531, 
    4.973192, 4.97331, 4.974496, 4.975257, 4.975863, 4.976406, 4.976948, 
    4.978693, 4.980071, 4.981329, 4.982737, 4.984304, 4.98608, 4.98801, 
    4.990017, 4.99169, 4.992681, 4.994704, 4.996451, 4.997856, 4.998842, 
    4.999298, 4.999086, 4.998041, 4.995966, 4.992651, 4.98787, 4.981419, 
    4.973136, 4.962947, 4.9509, 4.937212, 4.922284, 4.906702, 4.891196, 
    4.876576,
  // totalHeight(24,11, 0-49)
    4.928943, 4.934204, 4.939147, 4.943745, 4.947984, 4.95187, 4.955413, 
    4.958628, 4.961534, 4.964156, 4.966515, 4.968637, 4.97054, 4.972244, 
    4.973755, 4.973986, 4.97442, 4.975101, 4.975702, 4.976256, 4.976806, 
    4.978368, 4.97955, 4.980563, 4.981774, 4.983195, 4.984904, 4.986845, 
    4.988947, 4.990697, 4.991765, 4.993696, 4.995408, 4.996849, 4.997957, 
    4.998643, 4.998786, 4.998235, 4.996804, 4.994276, 4.990419, 4.985002, 
    4.977817, 4.968729, 4.957708, 4.944883, 4.930571, 4.91528, 4.899696, 
    4.884621,
  // totalHeight(24,12, 0-49)
    4.931442, 4.936534, 4.941318, 4.945765, 4.949864, 4.953617, 4.957031, 
    4.960122, 4.962908, 4.965411, 4.967651, 4.969649, 4.971423, 4.972981, 
    4.974318, 4.974725, 4.974307, 4.974916, 4.975528, 4.976114, 4.976694, 
    4.978027, 4.978982, 4.979725, 4.98072, 4.981984, 4.983621, 4.985569, 
    4.98778, 4.989639, 4.990843, 4.992671, 4.994336, 4.995801, 4.997019, 
    4.997913, 4.998381, 4.998281, 4.997436, 4.995634, 4.992631, 4.988174, 
    4.982021, 4.973984, 4.963962, 4.952005, 4.938346, 4.923423, 4.907864, 
    4.892451,
  // totalHeight(24,13, 0-49)
    4.934093, 4.939003, 4.943612, 4.947893, 4.951836, 4.955441, 4.958715, 
    4.961672, 4.964326, 4.966701, 4.968812, 4.970676, 4.972308, 4.973703, 
    4.974848, 4.975464, 4.974095, 4.974648, 4.975296, 4.975943, 4.976576, 
    4.977641, 4.978346, 4.978808, 4.97958, 4.980684, 4.982246, 4.984205, 
    4.986533, 4.988531, 4.989935, 4.991654, 4.993267, 4.994752, 4.996068, 
    4.997155, 4.997918, 4.99823, 4.997921, 4.996779, 4.994556, 4.990984, 
    4.985788, 4.978738, 4.969673, 4.958571, 4.94559, 4.931089, 4.915645, 
    4.900013,
  // totalHeight(24,14, 0-49)
    4.936921, 4.94163, 4.946046, 4.950143, 4.953909, 4.957345, 4.96046, 
    4.963262, 4.96577, 4.968, 4.969966, 4.971681, 4.973152, 4.974371, 
    4.975314, 4.976134, 4.973717, 4.97424, 4.974955, 4.975695, 4.976418, 
    4.977182, 4.977629, 4.977811, 4.978366, 4.979317, 4.980805, 4.982772, 
    4.985224, 4.987384, 4.989049, 4.990658, 4.992219, 4.993719, 4.995128, 
    4.996392, 4.997429, 4.998117, 4.998294, 4.997752, 4.996239, 4.993473, 
    4.989157, 4.983024, 4.974865, 4.964593, 4.952296, 4.938266, 4.923021, 
    4.907284,
  // totalHeight(24,15, 0-49)
    4.939954, 4.944445, 4.948641, 4.952525, 4.956085, 4.959326, 4.962252, 
    4.964876, 4.967212, 4.969275, 4.971076, 4.972627, 4.973923, 4.974956, 
    4.975694, 4.976676, 4.973099, 4.973635, 4.974455, 4.975329, 4.976182, 
    4.976626, 4.976819, 4.976738, 4.977095, 4.977906, 4.979325, 4.981301, 
    4.983872, 4.986211, 4.988193, 4.98969, 4.991199, 4.992713, 4.994207, 
    4.995636, 4.996924, 4.997959, 4.998579, 4.99858, 4.99771, 4.995675, 
    4.992167, 4.986881, 4.979572, 4.970099, 4.958487, 4.944963, 4.929991, 
    4.914255,
  // totalHeight(24,16, 0-49)
    4.943211, 4.947452, 4.951399, 4.955036, 4.958356, 4.961365, 4.964069, 
    4.966485, 4.968622, 4.970495, 4.972114, 4.973482, 4.974594, 4.975438, 
    4.975983, 4.977036, 4.972176, 4.972776, 4.97375, 4.974805, 4.975837, 
    4.975954, 4.975911, 4.9756, 4.975791, 4.976484, 4.977843, 4.979822, 
    4.982503, 4.985028, 4.98737, 4.988751, 4.990204, 4.991729, 4.993303, 
    4.994886, 4.996407, 4.997757, 4.998783, 4.999278, 4.99899, 4.997621, 
    4.994846, 4.990343, 4.983829, 4.97512, 4.964186, 4.9512, 4.936568, 
    4.920935,
  // totalHeight(24,17, 0-49)
    4.946694, 4.950654, 4.95431, 4.957654, 4.960692, 4.963429, 4.965877, 
    4.968051, 4.969965, 4.971627, 4.973047, 4.974223, 4.975149, 4.97581, 
    4.976184, 4.977188, 4.970901, 4.971617, 4.972795, 4.974083, 4.975348, 
    4.975148, 4.974903, 4.974407, 4.974476, 4.975085, 4.976398, 4.978378, 
    4.981153, 4.983857, 4.986584, 4.987842, 4.989233, 4.990761, 4.992407, 
    4.994132, 4.995866, 4.997506, 4.998901, 4.999847, 5.000089, 4.999326, 
    4.997222, 4.993437, 4.987666, 4.979686, 4.969424, 4.956998, 4.942767, 
    4.927331,
  // totalHeight(24,18, 0-49)
    4.950392, 4.954015, 4.957329, 4.960334, 4.963038, 4.965462, 4.96762, 
    4.969528, 4.9712, 4.972644, 4.973861, 4.974846, 4.975591, 4.976085, 
    4.976321, 4.97714, 4.969261, 4.970144, 4.971568, 4.973141, 4.974692, 
    4.974195, 4.973797, 4.973176, 4.973178, 4.973746, 4.975035, 4.977013, 
    4.97986, 4.982726, 4.985838, 4.986964, 4.988281, 4.9898, 4.991502, 
    4.99335, 4.99528, 4.997187, 4.998922, 5.000279, 5.001005, 5.000793, 
    4.999304, 4.996184, 4.991109, 4.983826, 4.974225, 4.962378, 4.948599, 
    4.933446,
  // totalHeight(24,19, 0-49)
    4.954257, 4.957479, 4.960381, 4.962982, 4.965306, 4.967378, 4.969222, 
    4.970854, 4.972284, 4.973517, 4.974545, 4.975358, 4.975943, 4.976294, 
    4.976423, 4.976936, 4.967296, 4.968376, 4.970076, 4.971971, 4.973859, 
    4.973104, 4.972607, 4.971929, 4.971931, 4.972509, 4.973804, 4.975785, 
    4.978683, 4.981678, 4.985153, 4.986128, 4.987349, 4.988836, 4.990572, 
    4.992523, 4.994625, 4.996772, 4.998816, 5.000549, 5.001719, 5.002016, 
    5.001093, 4.99859, 4.994166, 4.98755, 4.978599, 4.967349, 4.954068, 
    4.939276,
  // totalHeight(24,20, 0-49)
    4.959174, 4.962858, 4.966164, 4.969108, 4.971708, 4.973982, 4.975949, 
    4.977625, 4.979029, 4.980179, 4.981099, 4.981818, 4.982371, 4.982801, 
    4.983164, 30, 4.964798, 4.966055, 4.967796, 4.969609, 4.971327, 4.969703, 
    4.968443, 4.967083, 4.966592, 4.9669, 4.968161, 4.970348, 4.973696, 
    4.977341, 4.981765, 4.983172, 4.984841, 4.986776, 4.988951, 4.991327, 
    4.993841, 4.996396, 4.998845, 5.000997, 5.002602, 5.003364, 5.002938, 
    5.000969, 4.997112, 4.991087, 4.982724, 4.972033, 4.959246, 4.944842,
  // totalHeight(24,21, 0-49)
    4.963408, 4.966722, 4.969628, 4.972158, 4.974346, 4.976221, 4.977811, 
    4.979146, 4.980244, 4.981132, 4.981833, 4.982378, 4.982804, 4.983163, 
    4.983527, 30, 4.959586, 4.9611, 4.963162, 4.96533, 4.967396, 4.965482, 
    4.964082, 4.96265, 4.96222, 4.962704, 4.964239, 4.966779, 4.970561, 
    4.974705, 4.979818, 4.98141, 4.983339, 4.985602, 4.98816, 4.990963, 
    4.993931, 4.996956, 4.999882, 5.002509, 5.004585, 5.00581, 5.005842, 
    5.004326, 5.000915, 4.995324, 4.987371, 4.97705, 4.964567, 4.950371,
  // totalHeight(24,22, 0-49)
    4.967702, 4.970664, 4.973182, 4.975305, 4.977076, 4.978538, 4.979732, 
    4.980693, 4.981451, 4.982034, 4.982473, 4.982803, 4.983067, 4.983329, 
    4.983677, 30, 4.955086, 4.956829, 4.959173, 4.961654, 4.964025, 4.961829, 
    4.960271, 4.958739, 4.958321, 4.95891, 4.960636, 4.963431, 4.967537, 
    4.97206, 4.977712, 4.979404, 4.981507, 4.984018, 4.986888, 4.990057, 
    4.993435, 4.9969, 5.000288, 5.003388, 5.00594, 5.007639, 5.008145, 
    5.007098, 5.004148, 4.999008, 4.99149, 4.981569, 4.969436, 4.955513,
  // totalHeight(24,23, 0-49)
    4.971951, 4.974577, 4.976721, 4.978443, 4.979802, 4.980852, 4.98164, 
    4.982214, 4.98261, 4.982863, 4.983012, 4.983098, 4.983173, 4.983312, 
    4.983619, 30, 4.951283, 4.953178, 4.955709, 4.958392, 4.960952, 4.958478, 
    4.956745, 4.95508, 4.954624, 4.955256, 4.957099, 4.960074, 4.964422, 
    4.969233, 4.975299, 4.977072, 4.979327, 4.982063, 4.985225, 4.988744, 
    4.992522, 4.996426, 5.000281, 5.003865, 5.006908, 5.009098, 5.010088, 
    5.009516, 5.007031, 5.002338, 4.995245, 4.985715, 4.973922, 4.960277,
  // totalHeight(24,24, 0-49)
    4.976042, 4.978349, 4.980137, 4.981477, 4.982438, 4.983085, 4.983476, 
    4.983662, 4.983689, 4.983603, 4.983446, 4.983268, 4.98313, 4.983118, 
    4.983349, 30, 4.948518, 4.95047, 4.953073, 4.955839, 4.958478, 4.955807, 
    4.953943, 4.952183, 4.951692, 4.952342, 4.954256, 4.957346, 4.961858, 
    4.966876, 4.973243, 4.975129, 4.977551, 4.980509, 4.98394, 4.987772, 
    4.991901, 4.996183, 5.000436, 5.004429, 5.007885, 5.010486, 5.011881, 
    5.011705, 5.009609, 5.005295, 4.998567, 4.989384, 4.97791, 4.964542,
  // totalHeight(24,25, 0-49)
    4.979859, 4.981875, 4.983335, 4.984321, 4.984909, 4.985174, 4.985183, 
    4.984993, 4.984659, 4.984231, 4.983762, 4.983307, 4.982939, 4.982748, 
    4.982862, 30, 4.94658, 4.948485, 4.951038, 4.953754, 4.956346, 4.953585, 
    4.951666, 4.949878, 4.949385, 4.95006, 4.952026, 4.955197, 4.959819, 
    4.964978, 4.971531, 4.973589, 4.976222, 4.979423, 4.983128, 4.987259, 
    4.991705, 4.996318, 5.000906, 5.005232, 5.009016, 5.011939, 5.013646, 
    5.013772, 5.011967, 5.007938, 5.00149, 4.992584, 4.981378, 4.968261,
  // totalHeight(24,26, 0-49)
    4.983298, 4.98506, 4.986228, 4.986894, 4.987146, 4.987062, 4.986718, 
    4.986174, 4.985493, 4.984731, 4.983946, 4.983204, 4.982584, 4.982186, 
    4.982136, 30, 4.945513, 4.947264, 4.949642, 4.952173, 4.954591, 4.951852, 
    4.949958, 4.948216, 4.947764, 4.948481, 4.95049, 4.953713, 4.958396, 
    4.963634, 4.970265, 4.972566, 4.975461, 4.978936, 4.982924, 4.987339, 
    4.992069, 4.996956, 5.001805, 5.006377, 5.010392, 5.013525, 5.015426, 
    5.015734, 5.014105, 5.01025, 5.003979, 4.99526, 4.984254, 4.97135,
  // totalHeight(24,27, 0-49)
    4.986259, 4.987812, 4.988739, 4.989136, 4.989098, 4.988709, 4.988045, 
    4.987175, 4.986165, 4.985077, 4.983976, 4.982936, 4.982043, 4.9814, 
    4.981136, 30, 4.94546, 4.946948, 4.949024, 4.951235, 4.95335, 4.950716, 
    4.948902, 4.947252, 4.946861, 4.947614, 4.949643, 4.952878, 4.957563, 
    4.962814, 4.969408, 4.972008, 4.975201, 4.978966, 4.983234, 4.987912, 
    4.99288, 4.997982, 5.003019, 5.007753, 5.011899, 5.015141, 5.017131, 
    5.017511, 5.015946, 5.012156, 5.005963, 4.997341, 4.986464, 4.973726,
  // totalHeight(24,28, 0-49)
    4.988665, 4.990068, 4.990814, 4.991004, 4.990735, 4.990089, 4.989146, 
    4.98798, 4.986658, 4.985248, 4.983824, 4.982468, 4.981272, 4.980346, 
    4.979819, 30, 4.946815, 4.947936, 4.949587, 4.951346, 4.953032, 4.950542, 
    4.948813, 4.947252, 4.946893, 4.947637, 4.949623, 4.952797, 4.957403, 
    4.962586, 4.969032, 4.971952, 4.975448, 4.97949, 4.984002, 4.98889, 
    4.994031, 4.999268, 5.004402, 5.0092, 5.013378, 5.016623, 5.018593, 
    5.018941, 5.017337, 5.013512, 5.007304, 4.998701, 4.987891, 4.975283,
  // totalHeight(24,29, 0-49)
    4.990462, 4.991789, 4.992432, 4.992489, 4.992052, 4.991203, 4.990024, 
    4.988585, 4.986959, 4.985222, 4.983455, 4.981752, 4.980217, 4.978965, 
    4.978124, 30, 4.949393, 4.950053, 4.951162, 4.952341, 4.953464, 4.951066, 
    4.949343, 4.947788, 4.947369, 4.948007, 4.949859, 4.952889, 4.957327, 
    4.96235, 4.968523, 4.971735, 4.9755, 4.97978, 4.984496, 4.989554, 
    4.994829, 5.000166, 5.005371, 5.010205, 5.014393, 5.01762, 5.019548, 
    5.019832, 5.018151, 5.014245, 5.007967, 4.999325, 4.988527, 4.976,
  // totalHeight(24,30, 0-49)
    4.990738, 4.99121, 4.991029, 4.990311, 4.989165, 4.987687, 4.985961, 
    4.984056, 4.982023, 4.979897, 4.977703, 4.975448, 4.973134, 4.970758, 
    4.968334, 4.967433, 4.952801, 4.952506, 4.95306, 4.954014, 4.955168, 
    4.953628, 4.952737, 4.951961, 4.952108, 4.953052, 4.954916, 4.957685, 
    4.961609, 4.965942, 4.971194, 4.974047, 4.977447, 4.981374, 4.985769, 
    4.990544, 4.995582, 5.000725, 5.005774, 5.010484, 5.014568, 5.017704, 
    5.019542, 5.019734, 5.017958, 5.013961, 5.007609, 4.998928, 4.988154, 
    4.975735,
  // totalHeight(24,31, 0-49)
    4.991224, 4.991782, 4.991659, 4.990963, 4.989799, 4.988257, 4.986423, 
    4.984369, 4.982151, 4.979816, 4.977396, 4.974913, 4.972373, 4.969775, 
    4.967119, 4.966956, 4.953699, 4.952859, 4.952815, 4.953157, 4.953729, 
    4.952262, 4.951339, 4.950546, 4.950665, 4.951616, 4.953545, 4.956422, 
    4.960444, 4.964846, 4.969977, 4.973281, 4.977116, 4.981448, 4.986209, 
    4.991305, 4.996608, 5.001957, 5.007145, 5.011923, 5.016, 5.01905, 
    5.020725, 5.020681, 5.018607, 5.014267, 5.007555, 4.998531, 4.987468, 
    4.97485,
  // totalHeight(24,32, 0-49)
    4.990952, 4.991582, 4.991526, 4.990881, 4.989748, 4.988213, 4.986357, 
    4.984251, 4.981956, 4.979523, 4.976988, 4.974381, 4.971712, 4.968981, 
    4.966177, 4.966247, 4.954534, 4.953211, 4.952619, 4.952398, 4.952437, 
    4.951101, 4.950212, 4.94947, 4.949618, 4.950622, 4.952628, 4.955601, 
    4.959674, 4.964085, 4.969033, 4.97274, 4.976955, 4.98163, 4.986691, 
    4.992035, 4.99753, 5.003008, 5.008257, 5.013021, 5.017007, 5.019885, 
    5.02131, 5.020944, 5.018488, 5.013731, 5.006595, 4.997181, 4.985804, 
    4.972989,
  // totalHeight(24,33, 0-49)
    4.989976, 4.990683, 4.990708, 4.990148, 4.98909, 4.987619, 4.985811, 
    4.983734, 4.981448, 4.979006, 4.976447, 4.973802, 4.971087, 4.968307, 
    4.965442, 4.965351, 4.955271, 4.953551, 4.952481, 4.951764, 4.95134, 
    4.950182, 4.949387, 4.948767, 4.949002, 4.950088, 4.952173, 4.955213, 
    4.959281, 4.96364, 4.968359, 4.972418, 4.976954, 4.981907, 4.987197, 
    4.992716, 4.998327, 5.003853, 5.00908, 5.013745, 5.017552, 5.020169, 
    5.021256, 5.020481, 5.017564, 5.012319, 5.004707, 4.994871, 4.983172, 
    4.970181,
  // totalHeight(24,34, 0-49)
    4.988362, 4.989154, 4.989285, 4.98884, 4.9879, 4.986543, 4.984841, 
    4.982858, 4.980649, 4.978268, 4.975753, 4.973141, 4.970451, 4.967691, 
    4.964846, 4.964324, 4.955907, 4.953883, 4.95241, 4.951271, 4.950449, 
    4.949511, 4.948865, 4.948426, 4.948793, 4.949985, 4.952144, 4.955214, 
    4.959218, 4.96347, 4.967926, 4.972286, 4.977082, 4.982247, 4.987697, 
    4.993318, 4.998965, 5.004459, 5.009578, 5.014056, 5.017594, 5.019861, 
    5.020521, 5.019255, 5.015803, 5.010012, 5.001885, 4.991614, 4.979609, 
    4.96648,
  // totalHeight(24,35, 0-49)
    4.986187, 4.987076, 4.987331, 4.987029, 4.986242, 4.985043, 4.983495, 
    4.981658, 4.979582, 4.977318, 4.974906, 4.972382, 4.969771, 4.967087, 
    4.964324, 4.963235, 4.956457, 4.954219, 4.952422, 4.950934, 4.949782, 
    4.94909, 4.948639, 4.948434, 4.94897, 4.950284, 4.952501, 4.955562, 
    4.959439, 4.963533, 4.967704, 4.972306, 4.977299, 4.98261, 4.988148, 
    4.993796, 4.9994, 5.004778, 5.009702, 5.013903, 5.017081, 5.018907, 
    5.019053, 5.017218, 5.013171, 5.006792, 4.998133, 4.987436, 4.975163, 
    4.961967,
  // totalHeight(24,36, 0-49)
    4.983537, 4.98453, 4.984925, 4.98479, 4.984187, 4.983179, 4.981824, 
    4.980174, 4.978276, 4.976174, 4.973908, 4.971516, 4.969026, 4.966462, 
    4.963827, 4.962144, 4.956951, 4.95458, 4.952532, 4.950767, 4.949354, 
    4.948923, 4.9487, 4.948773, 4.949505, 4.950946, 4.953201, 4.956208, 
    4.959899, 4.963787, 4.967659, 4.972442, 4.977566, 4.982953, 4.988503, 
    4.994096, 4.999576, 5.004749, 5.009388, 5.013221, 5.015947, 5.017244, 
    5.016798, 5.014329, 5.009636, 5.002648, 4.993464, 4.982381, 4.969909, 
    4.956739,
  // totalHeight(24,37, 0-49)
    4.980508, 4.981606, 4.982151, 4.982196, 4.981798, 4.981007, 4.979875, 
    4.978444, 4.976758, 4.974855, 4.972772, 4.970547, 4.968214, 4.965799, 
    4.963324, 4.9611, 4.957419, 4.954983, 4.952751, 4.950772, 4.949162, 
    4.949, 4.949028, 4.949411, 4.950358, 4.951927, 4.954195, 4.957103, 
    4.96055, 4.96419, 4.967753, 4.97265, 4.977834, 4.983218, 4.988704, 
    4.99416, 4.999428, 5.004307, 5.008569, 5.01194, 5.014123, 5.014809, 
    5.013699, 5.010541, 5.005176, 4.997579, 4.987903, 4.976503, 4.963933, 
    4.950914,
  // totalHeight(24,38, 0-49)
    4.977201, 4.978397, 4.979091, 4.979325, 4.979144, 4.978589, 4.977698, 
    4.976512, 4.975065, 4.97339, 4.971519, 4.969489, 4.967337, 4.965096, 
    4.962796, 4.960145, 4.957889, 4.955441, 4.953079, 4.950952, 4.949204, 
    4.949308, 4.949604, 4.950312, 4.951482, 4.953172, 4.955426, 4.958192, 
    4.96134, 4.964695, 4.967939, 4.972879, 4.978047, 4.983353, 4.988689, 
    4.993921, 4.998884, 5.003378, 5.007168, 5.009984, 5.011538, 5.011535, 
    5.0097, 5.005819, 4.999774, 4.991597, 4.981497, 4.96988, 4.957343, 
    4.944621,
  // totalHeight(24,39, 0-49)
    4.973715, 4.974999, 4.975837, 4.976258, 4.976297, 4.975984, 4.975348, 
    4.974423, 4.973234, 4.971807, 4.970172, 4.968362, 4.966412, 4.964359, 
    4.962245, 4.959305, 4.958379, 4.955961, 4.953523, 4.9513, 4.949468, 
    4.949832, 4.950396, 4.951439, 4.95283, 4.954629, 4.956837, 4.959415, 
    4.962219, 4.965253, 4.968168, 4.973073, 4.978147, 4.983289, 4.988388, 
    4.993306, 4.997871, 5.001883, 5.005105, 5.007277, 5.00812, 5.007362, 
    5.004759, 5.000136, 4.993432, 4.984732, 4.974305, 4.962605, 4.950256, 
    4.938003,
  // totalHeight(24,40, 0-49)
    4.970154, 4.971507, 4.972474, 4.973073, 4.973326, 4.973255, 4.972881, 
    4.972223, 4.971304, 4.970143, 4.968762, 4.967189, 4.965458, 4.963606, 
    4.96168, 4.958601, 4.958908, 4.956546, 4.954076, 4.951808, 4.949941, 
    4.950551, 4.951377, 4.952746, 4.95435, 4.956237, 4.958365, 4.960715, 
    4.96313, 4.96581, 4.968381, 4.973172, 4.978065, 4.982956, 4.987728, 
    4.992238, 4.996309, 4.999742, 5.002305, 5.003745, 5.003803, 5.002235, 
    4.998837, 4.993484, 4.986167, 4.977036, 4.966411, 4.954787, 4.942811, 
    4.931215,
  // totalHeight(24,41, 0-49)
    4.966611, 4.968009, 4.969085, 4.969845, 4.970301, 4.970465, 4.970348, 
    4.969962, 4.969318, 4.968431, 4.967318, 4.965998, 4.964501, 4.962861, 
    4.961126, 4.958048, 4.959484, 4.957199, 4.954734, 4.952466, 4.950603, 
    4.951441, 4.952514, 4.954194, 4.955987, 4.957934, 4.959948, 4.96203, 
    4.964015, 4.966311, 4.968513, 4.973105, 4.977732, 4.982281, 4.98663, 
    4.990634, 4.994115, 4.996872, 4.998685, 4.999315, 4.998528, 4.996117, 
    4.99192, 4.985871, 4.978022, 4.96858, 4.957916, 4.946559, 4.935153, 
    4.924411,
  // totalHeight(24,42, 0-49)
    4.963175, 4.964589, 4.965748, 4.966649, 4.96729, 4.967675, 4.967805, 
    4.967684, 4.967317, 4.966709, 4.96587, 4.964814, 4.963562, 4.962146, 
    4.960603, 4.957645, 4.960103, 4.957912, 4.955489, 4.953257, 4.951434, 
    4.952474, 4.953773, 4.955733, 4.957686, 4.959659, 4.961521, 4.963294, 
    4.964817, 4.966691, 4.968498, 4.972802, 4.977069, 4.98118, 4.985012, 
    4.988411, 4.991204, 4.993195, 4.994174, 4.993927, 4.992252, 4.988981, 
    4.984013, 4.977334, 4.969066, 4.959468, 4.948955, 4.938068, 4.927447, 
    4.917754,
  // totalHeight(24,43, 0-49)
    4.959915, 4.961318, 4.962533, 4.963548, 4.964352, 4.964938, 4.965301, 
    4.965435, 4.965337, 4.965007, 4.964446, 4.963661, 4.962666, 4.96148, 
    4.960136, 4.957391, 4.960761, 4.95868, 4.956325, 4.954162, 4.952404, 
    4.953622, 4.955115, 4.957315, 4.959389, 4.961347, 4.963018, 4.964441, 
    4.965469, 4.966885, 4.968258, 4.972181, 4.975993, 4.979571, 4.982786, 
    4.985485, 4.987495, 4.988636, 4.988711, 4.987537, 4.984951, 4.980837, 
    4.97515, 4.967946, 4.959401, 4.94983, 4.939674, 4.929479, 4.919853, 
    4.911402,
  // totalHeight(24,44, 0-49)
    4.956895, 4.958255, 4.959497, 4.960596, 4.961537, 4.962301, 4.962876, 
    4.963249, 4.963411, 4.963352, 4.963067, 4.962556, 4.961821, 4.960875, 
    4.959737, 4.957268, 4.961443, 4.959482, 4.957224, 4.955157, 4.953481, 
    4.954848, 4.956501, 4.958893, 4.961037, 4.962934, 4.964368, 4.965406, 
    4.965909, 4.966825, 4.967713, 4.971162, 4.974424, 4.97737, 4.979871, 
    4.981776, 4.98292, 4.983132, 4.98225, 4.98012, 4.976628, 4.971716, 
    4.965401, 4.957804, 4.949159, 4.93982, 4.930246, 4.920966, 4.912542, 
    4.905505,
  // totalHeight(24,45, 0-49)
    4.954153, 4.955442, 4.956679, 4.957835, 4.958883, 4.959798, 4.960562, 
    4.961154, 4.961558, 4.961758, 4.961742, 4.961503, 4.961034, 4.960333, 
    4.959406, 4.957256, 4.962121, 4.960298, 4.958159, 4.956203, 4.954621, 
    4.95611, 4.957882, 4.960408, 4.962569, 4.964353, 4.96551, 4.966124, 
    4.966069, 4.96644, 4.966787, 4.969665, 4.972278, 4.974496, 4.976191, 
    4.977215, 4.977416, 4.976646, 4.974771, 4.971683, 4.967322, 4.961689, 
    4.95487, 4.947047, 4.938503, 4.929619, 4.920855, 4.912706, 4.905671, 
    4.900196,
  // totalHeight(24,46, 0-49)
    4.951709, 4.952902, 4.954107, 4.955286, 4.956411, 4.957448, 4.958375, 
    4.959161, 4.959786, 4.960229, 4.960472, 4.960496, 4.96029, 4.959839, 
    4.959132, 4.957314, 4.962758, 4.961088, 4.95909, 4.957263, 4.955777, 
    4.957358, 4.959206, 4.961804, 4.963924, 4.965539, 4.966373, 4.966525, 
    4.965885, 4.965662, 4.965401, 4.967614, 4.969483, 4.970881, 4.971683, 
    4.97175, 4.970951, 4.969162, 4.966289, 4.962273, 4.957111, 4.950871, 
    4.943702, 4.935844, 4.927619, 4.919419, 4.911686, 4.904869, 4.899387, 
    4.895587,
  // totalHeight(24,47, 0-49)
    4.949562, 4.950633, 4.951778, 4.952954, 4.954126, 4.955256, 4.956315, 
    4.957269, 4.95809, 4.958755, 4.959237, 4.959513, 4.959562, 4.959362, 
    4.958882, 4.957393, 4.963307, 4.961806, 4.959966, 4.958274, 4.956888, 
    4.958531, 4.960414, 4.963019, 4.965039, 4.966431, 4.966897, 4.96655, 
    4.965296, 4.964425, 4.963489, 4.964943, 4.965979, 4.966473, 4.966308, 
    4.965361, 4.963523, 4.960705, 4.956856, 4.951973, 4.946115, 4.939414, 
    4.932077, 4.924395, 4.916712, 4.90942, 4.902925, 4.897609, 4.893805, 
    4.891757,
  // totalHeight(24,48, 0-49)
    4.94768, 4.948614, 4.949677, 4.950824, 4.952013, 4.953206, 4.954365, 
    4.955455, 4.956445, 4.957305, 4.958005, 4.958517, 4.958811, 4.958855, 
    4.958607, 4.95743, 4.963704, 4.962394, 4.960724, 4.959174, 4.957884, 
    4.959568, 4.961443, 4.963991, 4.965849, 4.966964, 4.967022, 4.966144, 
    4.964246, 4.962679, 4.960994, 4.961605, 4.961727, 4.961245, 4.960056, 
    4.958057, 4.95517, 4.951344, 4.946577, 4.940922, 4.934504, 4.927511, 
    4.920208, 4.912917, 4.905994, 4.899813, 4.894729, 4.891049, 4.889009, 
    4.888746,
  // totalHeight(24,49, 0-49)
    4.945692, 4.946275, 4.947063, 4.948007, 4.949056, 4.950163, 4.951286, 
    4.952384, 4.953416, 4.954346, 4.955135, 4.95574, 4.956119, 4.956212, 
    4.955952, 4.954215, 4.967573, 4.965439, 4.962609, 4.960008, 4.957872, 
    4.961558, 4.965416, 4.970356, 4.973582, 4.975026, 4.974078, 4.971011, 
    4.965668, 4.960866, 4.955824, 4.955507, 4.954542, 4.952848, 4.950368, 
    4.947054, 4.942887, 4.937885, 4.932127, 4.925748, 4.918957, 4.912019, 
    4.905252, 4.899001, 4.89361, 4.88939, 4.886611, 4.885452, 4.886003, 
    4.888259,
  // totalHeight(25,0, 0-49)
    4.925933, 4.931124, 4.936015, 4.940607, 4.944907, 4.948923, 4.952667, 
    4.956147, 4.959369, 4.962331, 4.965029, 4.967461, 4.969619, 4.971503, 
    4.973116, 4.974247, 4.975694, 4.976534, 4.977195, 4.977763, 4.978303, 
    4.97908, 4.979904, 4.98088, 4.98202, 4.983343, 4.984835, 4.986478, 
    4.988221, 4.990023, 4.991735, 4.993485, 4.994883, 4.995748, 4.995881, 
    4.995065, 4.993076, 4.989686, 4.984684, 4.977894, 4.969201, 4.95857, 
    4.946083, 4.931956, 4.916556, 4.9004, 4.884132, 4.868479, 4.854189, 
    4.841959,
  // totalHeight(25,1, 0-49)
    4.927026, 4.932236, 4.937124, 4.941692, 4.945944, 4.949895, 4.953556, 
    4.956938, 4.960046, 4.962883, 4.965448, 4.967741, 4.96976, 4.971508, 
    4.972995, 4.97379, 4.975451, 4.976137, 4.976635, 4.977072, 4.977521, 
    4.978458, 4.979441, 4.980615, 4.981967, 4.983503, 4.985191, 4.98702, 
    4.988934, 4.99092, 4.992792, 4.994941, 4.996752, 4.998055, 4.998661, 
    4.998352, 4.996904, 4.994087, 4.98968, 4.983487, 4.975367, 4.965255, 
    4.953193, 4.939358, 4.924083, 4.907857, 4.891315, 4.875189, 4.860251, 
    4.847242,
  // totalHeight(25,2, 0-49)
    4.928236, 4.933441, 4.938304, 4.942826, 4.947015, 4.950887, 4.954455, 
    4.95773, 4.960721, 4.963433, 4.965869, 4.968032, 4.969925, 4.971556, 
    4.972939, 4.973425, 4.975278, 4.975841, 4.976205, 4.97653, 4.976901, 
    4.977989, 4.979106, 4.980435, 4.981947, 4.983635, 4.985459, 4.987404, 
    4.989417, 4.991495, 4.993425, 4.995854, 4.997965, 4.999597, 5.000571, 
    5.000686, 4.999723, 4.997451, 4.993648, 4.988107, 4.980661, 4.97122, 
    4.959781, 4.946479, 4.931597, 4.91558, 4.899025, 4.882655, 4.867242, 
    4.853558,
  // totalHeight(25,3, 0-49)
    4.929566, 4.934745, 4.939562, 4.944022, 4.948135, 4.951917, 4.955383, 
    4.958548, 4.961421, 4.964013, 4.966328, 4.968372, 4.970154, 4.971688, 
    4.972991, 4.973203, 4.975204, 4.975671, 4.975931, 4.976166, 4.976469, 
    4.977692, 4.978915, 4.980353, 4.981971, 4.983752, 4.985653, 4.987656, 
    4.989704, 4.991798, 4.993697, 4.996298, 4.998598, 5.000453, 5.001705, 
    5.00216, 5.001616, 4.99985, 4.996643, 4.991779, 4.985082, 4.976425, 
    4.965772, 4.953203, 4.938946, 4.923386, 4.907069, 4.890676, 4.874971, 
    4.860731,
  // totalHeight(25,4, 0-49)
    4.931008, 4.93614, 4.940896, 4.945281, 4.949308, 4.952993, 4.956354, 
    4.959407, 4.962167, 4.964643, 4.966847, 4.968788, 4.970478, 4.971931, 
    4.973177, 4.973155, 4.975237, 4.975637, 4.975821, 4.975992, 4.976242, 
    4.977576, 4.978874, 4.98037, 4.982038, 4.983856, 4.98578, 4.987794, 
    4.98983, 4.991879, 4.993676, 4.996348, 4.998741, 5.000727, 5.002164, 
    5.002882, 5.002693, 5.001389, 4.998754, 4.994576, 4.988664, 4.980871, 
    4.971121, 4.959445, 4.946002, 4.931112, 4.915251, 4.899047, 4.883229, 
    4.868569,
  // totalHeight(25,5, 0-49)
    4.932553, 4.937619, 4.942299, 4.9466, 4.950532, 4.954118, 4.957373, 
    4.960318, 4.962967, 4.965339, 4.967442, 4.969292, 4.970905, 4.9723, 
    4.973505, 4.973295, 4.975376, 4.975733, 4.975873, 4.975999, 4.976211, 
    4.977631, 4.978968, 4.980473, 4.982137, 4.983939, 4.985843, 4.987827, 
    4.98982, 4.991777, 4.993423, 4.996082, 4.998482, 5.000516, 5.002064, 
    5.002976, 5.003079, 5.002186, 5.000093, 4.996589, 4.991478, 4.984593, 
    4.975825, 4.965151, 4.952667, 4.938615, 4.923396, 4.907567, 4.891808, 
    4.876867,
  // totalHeight(25,6, 0-49)
    4.934185, 4.93917, 4.943763, 4.94797, 4.951805, 4.955288, 4.95844, 
    4.961281, 4.963829, 4.966102, 4.968116, 4.96989, 4.97144, 4.97279, 
    4.973968, 4.973625, 4.975606, 4.975941, 4.976063, 4.97617, 4.976358, 
    4.977833, 4.979174, 4.980636, 4.982246, 4.983988, 4.985836, 4.987762, 
    4.989691, 4.991532, 4.992995, 4.995569, 4.997908, 4.999924, 5.001517, 
    5.00256, 5.002903, 5.002374, 5.000784, 4.997931, 4.993614, 4.987652, 
    4.979905, 4.970301, 4.958872, 4.945784, 4.931354, 4.916058, 4.900511, 
    4.885429,
  // totalHeight(25,7, 0-49)
    4.935893, 4.940784, 4.94528, 4.949388, 4.953124, 4.956505, 4.959556, 
    4.962297, 4.964751, 4.966934, 4.968871, 4.970577, 4.972075, 4.973391, 
    4.974547, 4.974128, 4.975905, 4.976233, 4.976362, 4.976471, 4.976653, 
    4.97815, 4.979456, 4.980828, 4.98234, 4.983981, 4.985743, 4.987593, 
    4.989452, 4.991168, 4.992439, 4.994873, 4.997096, 4.999042, 5.000629, 
    5.001756, 5.002291, 5.002082, 5.000955, 4.998718, 4.995172, 4.990123, 
    4.983405, 4.974901, 4.964583, 4.952542, 4.939005, 4.924366, 4.909166, 
    4.894073,
  // totalHeight(25,8, 0-49)
    4.937671, 4.942457, 4.946848, 4.950853, 4.954486, 4.957766, 4.960718, 
    4.963364, 4.965728, 4.96783, 4.969694, 4.971343, 4.972795, 4.974077, 
    4.975214, 4.97478, 4.976242, 4.976571, 4.97673, 4.976866, 4.977058, 
    4.97854, 4.979775, 4.981012, 4.982388, 4.983896, 4.985551, 4.987316, 
    4.98911, 4.990705, 4.991796, 4.994046, 4.996115, 4.997952, 4.999499, 
    5.00067, 5.001359, 5.001431, 5.000728, 4.999069, 4.996257, 4.992092, 
    4.986383, 4.978979, 4.969792, 4.958836, 4.946263, 4.932373, 4.91763, 
    4.902642,
  // totalHeight(25,9, 0-49)
    4.939522, 4.944192, 4.948471, 4.952366, 4.955894, 4.959072, 4.961926, 
    4.964479, 4.966755, 4.96878, 4.970574, 4.972166, 4.973575, 4.974823, 
    4.975928, 4.975544, 4.976576, 4.976916, 4.977123, 4.977306, 4.977529, 
    4.978956, 4.980087, 4.981149, 4.982355, 4.983707, 4.985243, 4.986919, 
    4.988662, 4.990154, 4.991093, 4.993133, 4.995021, 4.996726, 4.998206, 
    4.999397, 5.00021, 5.000529, 5.000213, 4.999092, 4.996973, 4.993648, 
    4.988911, 4.982576, 4.974506, 4.964649, 4.953072, 4.939991, 4.92579, 
    4.911009,
  // totalHeight(25,10, 0-49)
    4.941456, 4.945998, 4.950157, 4.953936, 4.957352, 4.960425, 4.963178, 
    4.965636, 4.967824, 4.96977, 4.971497, 4.973028, 4.974387, 4.975594, 
    4.976652, 4.976379, 4.976869, 4.977222, 4.977496, 4.977747, 4.978018, 
    4.979352, 4.980344, 4.981201, 4.982213, 4.983394, 4.984804, 4.986394, 
    4.988105, 4.989521, 4.990354, 4.992166, 4.993861, 4.99542, 4.99682, 
    4.998015, 4.998931, 4.999473, 4.999509, 4.998883, 4.997409, 4.994874, 
    4.991057, 4.985744, 4.978755, 4.969977, 4.959402, 4.947165, 4.933567, 
    4.919079,
  // totalHeight(25,11, 0-49)
    4.943488, 4.947892, 4.951918, 4.955572, 4.958869, 4.961828, 4.964473, 
    4.96683, 4.968925, 4.970785, 4.972435, 4.973901, 4.975202, 4.976351, 
    4.977344, 4.977236, 4.977071, 4.977445, 4.9778, 4.978139, 4.978481, 
    4.979679, 4.980506, 4.981133, 4.981936, 4.982936, 4.984219, 4.985733, 
    4.98743, 4.988805, 4.98959, 4.991169, 4.992666, 4.994079, 4.995396, 
    4.996587, 4.997594, 4.998336, 4.998695, 4.998528, 4.99765, 4.995848, 
    4.992891, 4.988542, 4.982579, 4.97484, 4.96525, 4.953867, 4.940912, 
    4.926785,
  // totalHeight(25,12, 0-49)
    4.94564, 4.949892, 4.953773, 4.957288, 4.960452, 4.963284, 4.965809, 
    4.968053, 4.970044, 4.971808, 4.973372, 4.974759, 4.975985, 4.977059, 
    4.97797, 4.978063, 4.977129, 4.977533, 4.97799, 4.978438, 4.978873, 
    4.979895, 4.980533, 4.980914, 4.981503, 4.982321, 4.983479, 4.984927, 
    4.986634, 4.988007, 4.988809, 4.990157, 4.991462, 4.992733, 4.993971, 
    4.995159, 4.996251, 4.997179, 4.997838, 4.998092, 4.997764, 4.996637, 
    4.994474, 4.991019, 4.986021, 4.979267, 4.970627, 4.960088, 4.947798, 
    4.934089,
  // totalHeight(25,13, 0-49)
    4.947933, 4.952016, 4.955732, 4.959089, 4.962103, 4.964792, 4.967181, 
    4.969296, 4.971166, 4.972819, 4.97428, 4.975571, 4.976707, 4.977689, 
    4.978497, 4.978809, 4.976994, 4.977444, 4.978021, 4.978601, 4.979153, 
    4.979963, 4.980396, 4.980526, 4.980901, 4.981544, 4.982584, 4.983975, 
    4.985711, 4.987123, 4.988012, 4.989138, 4.990263, 4.991405, 4.992577, 
    4.993766, 4.994943, 4.996046, 4.996986, 4.997628, 4.997803, 4.997297, 
    4.995863, 4.99323, 4.989122, 4.983292, 4.975555, 4.965837, 4.95422, 
    4.94097,
  // totalHeight(25,14, 0-49)
    4.950387, 4.954278, 4.957808, 4.960986, 4.963825, 4.966348, 4.968579, 
    4.970545, 4.972275, 4.973796, 4.975134, 4.976312, 4.977338, 4.97821, 
    4.978907, 4.979425, 4.97661, 4.97713, 4.977851, 4.978589, 4.979284, 
    4.979852, 4.980071, 4.979954, 4.980126, 4.980606, 4.981539, 4.982883, 
    4.984664, 4.98615, 4.987199, 4.988118, 4.989079, 4.990109, 4.991226, 
    4.99243, 4.993695, 4.994971, 4.996171, 4.997174, 4.99781, 4.99787, 
    4.997099, 4.995217, 4.991927, 4.98695, 4.980062, 4.971135, 4.960188, 
    4.947428,
  // totalHeight(25,15, 0-49)
    4.953012, 4.956685, 4.960002, 4.96297, 4.965608, 4.967937, 4.969985, 
    4.971778, 4.973346, 4.974717, 4.975914, 4.976958, 4.977856, 4.978607, 
    4.979187, 4.979874, 4.975935, 4.976555, 4.977448, 4.97837, 4.979236, 
    4.979536, 4.979541, 4.979192, 4.97918, 4.979517, 4.980358, 4.981665, 
    4.983503, 4.985093, 4.986369, 4.987097, 4.987914, 4.988852, 4.989933, 
    4.991162, 4.992521, 4.993965, 4.995416, 4.996754, 4.997815, 4.998388, 
    4.998218, 4.997016, 4.99447, 4.990279, 4.98418, 4.976004, 4.965717, 
    4.95347,
  // totalHeight(25,16, 0-49)
    4.955808, 4.959229, 4.9623, 4.965026, 4.967431, 4.969538, 4.971376, 
    4.972972, 4.974357, 4.975558, 4.976596, 4.97749, 4.978249, 4.978869, 
    4.979337, 4.980128, 4.974936, 4.975688, 4.976779, 4.977916, 4.978982, 
    4.978996, 4.978796, 4.978239, 4.978075, 4.978295, 4.979061, 4.980342, 
    4.982244, 4.983959, 4.98552, 4.986079, 4.986772, 4.987638, 4.9887, 
    4.989968, 4.99143, 4.993042, 4.994732, 4.996383, 4.997833, 4.998872, 
    4.999245, 4.998656, 4.996783, 4.993306, 4.987936, 4.98047, 4.970826, 
    4.959108,
  // totalHeight(25,17, 0-49)
    4.958763, 4.961892, 4.964672, 4.96712, 4.969258, 4.971113, 4.972718, 
    4.974096, 4.975282, 4.976298, 4.977165, 4.9779, 4.978511, 4.979, 
    4.979367, 4.980179, 4.9736, 4.974513, 4.975829, 4.977204, 4.978499, 
    4.97822, 4.977831, 4.977103, 4.976825, 4.976961, 4.977675, 4.978942, 
    4.980911, 4.982769, 4.984655, 4.985065, 4.985654, 4.986466, 4.987527, 
    4.988847, 4.990417, 4.992199, 4.994118, 4.99606, 4.997868, 4.99933, 
    5.000191, 5.000153, 4.998885, 4.996056, 4.991358, 4.984556, 4.975537, 
    4.964358,
  // totalHeight(25,18, 0-49)
    4.961843, 4.964629, 4.967072, 4.969197, 4.971034, 4.972611, 4.973962, 
    4.975113, 4.976092, 4.976921, 4.977616, 4.97819, 4.978654, 4.979015, 
    4.979291, 4.980046, 4.971954, 4.973047, 4.974599, 4.976233, 4.977781, 
    4.977211, 4.976659, 4.975799, 4.975451, 4.975545, 4.976236, 4.977504, 
    4.979541, 4.981548, 4.983785, 4.984062, 4.984563, 4.985336, 4.986408, 
    4.98779, 4.989474, 4.991421, 4.993559, 4.995777, 4.997911, 4.999756, 
    5.001056, 5.001511, 5.000786, 4.998543, 4.99446, 4.988282, 4.979865, 
    4.969234,
  // totalHeight(25,19, 0-49)
    4.965, 4.967378, 4.969427, 4.971184, 4.972685, 4.973964, 4.975053, 
    4.975977, 4.976758, 4.977411, 4.977946, 4.978371, 4.978695, 4.978937, 
    4.979131, 4.97977, 4.970062, 4.97134, 4.973125, 4.975019, 4.976834, 
    4.975983, 4.975299, 4.974353, 4.973983, 4.974082, 4.974786, 4.976074, 
    4.978185, 4.980337, 4.982932, 4.983087, 4.983509, 4.98425, 4.985336, 
    4.986781, 4.988577, 4.990685, 4.993031, 4.995503, 4.99794, 5.000132, 
    5.001826, 5.002723, 5.002485, 5.000772, 4.997253, 4.991659, 4.983825, 
    4.973745,
  // totalHeight(25,20, 0-49)
    4.96907, 4.971853, 4.97428, 4.976379, 4.978179, 4.979703, 4.980981, 
    4.982036, 4.982894, 4.983582, 4.984131, 4.98457, 4.984934, 4.985262, 
    4.9856, 30, 4.967362, 4.968657, 4.970433, 4.97227, 4.973977, 4.972389, 
    4.971055, 4.969516, 4.968708, 4.968553, 4.969211, 4.970665, 4.973172, 
    4.975917, 4.979388, 4.979959, 4.980811, 4.981984, 4.98349, 4.985337, 
    4.98751, 4.989974, 4.992662, 4.995465, 4.99823, 5.000757, 5.002801, 
    5.00407, 5.004237, 5.002963, 4.999919, 4.994827, 4.987511, 4.977941,
  // totalHeight(25,21, 0-49)
    4.972409, 4.974806, 4.976856, 4.978595, 4.980055, 4.981269, 4.982268, 
    4.983077, 4.983721, 4.984225, 4.984614, 4.984921, 4.985179, 4.985434, 
    4.985746, 30, 4.962254, 4.963721, 4.965726, 4.967824, 4.969792, 4.9679, 
    4.966414, 4.964807, 4.964072, 4.964111, 4.965068, 4.966903, 4.969873, 
    4.97314, 4.977301, 4.978094, 4.979231, 4.980741, 4.982622, 4.984862, 
    4.987442, 4.990312, 4.993392, 4.996568, 4.999682, 5.002536, 5.004883, 
    5.006442, 5.00689, 5.005895, 5.003135, 4.998338, 4.991322, 4.982051,
  // totalHeight(25,22, 0-49)
    4.97575, 4.977777, 4.979461, 4.980845, 4.981971, 4.982874, 4.983584, 
    4.984133, 4.984543, 4.984839, 4.985049, 4.985203, 4.985339, 4.98551, 
    4.985789, 30, 4.957802, 4.959422, 4.961627, 4.96395, 4.966136, 4.963939, 
    4.962275, 4.960557, 4.959836, 4.959994, 4.961162, 4.963283, 4.966613, 
    4.970295, 4.975018, 4.975973, 4.977332, 4.97912, 4.981323, 4.983923, 
    4.986884, 4.990145, 4.993617, 4.997175, 5.000654, 5.003854, 5.006526, 
    5.008392, 5.009137, 5.008434, 5.005967, 5.001472, 4.994767, 4.985815,
  // totalHeight(25,23, 0-49)
    4.97903, 4.9807, 4.98203, 4.983072, 4.98387, 4.984463, 4.984885, 
    4.985168, 4.985334, 4.985412, 4.985426, 4.985411, 4.985411, 4.985483, 
    4.985715, 30, 4.953951, 4.955665, 4.95799, 4.960441, 4.962743, 4.960247, 
    4.958386, 4.956528, 4.955769, 4.955982, 4.957291, 4.959627, 4.96324, 
    4.967253, 4.972426, 4.973531, 4.9751, 4.977151, 4.979666, 4.982618, 
    4.98596, 4.98962, 4.993496, 4.997456, 5.001327, 5.004899, 5.007923, 
    5.010116, 5.011169, 5.010761, 5.00858, 5.00437, 4.997954, 4.989296,
  // totalHeight(25,24, 0-49)
    4.982182, 4.983513, 4.984507, 4.985221, 4.985703, 4.985996, 4.986135, 
    4.98615, 4.98607, 4.985919, 4.985728, 4.985533, 4.98538, 4.985335, 
    4.985494, 30, 4.951048, 4.95278, 4.955128, 4.957605, 4.959929, 4.957211, 
    4.9552, 4.953234, 4.952438, 4.952682, 4.954084, 4.956569, 4.960389, 
    4.964658, 4.970174, 4.971457, 4.973247, 4.975561, 4.978374, 4.98165, 
    4.985334, 4.989345, 4.993575, 4.997882, 5.002086, 5.005975, 5.009296, 
    5.011769, 5.013084, 5.012925, 5.010993, 5.007029, 5.000869, 4.992476,
  // totalHeight(25,25, 0-49)
    4.985147, 4.986164, 4.986844, 4.98725, 4.987433, 4.987438, 4.9873, 
    4.987053, 4.986725, 4.986343, 4.985937, 4.985548, 4.985225, 4.98504, 
    4.985095, 30, 4.948891, 4.950555, 4.952825, 4.955217, 4.957455, 4.95462, 
    4.952531, 4.950522, 4.949719, 4.949996, 4.95147, 4.954067, 4.958037, 
    4.962492, 4.968243, 4.969755, 4.971803, 4.974401, 4.977515, 4.981103, 
    4.985105, 4.989431, 4.993968, 4.998568, 5.003051, 5.007197, 5.010757, 
    5.013449, 5.014969, 5.015006, 5.013266, 5.009499, 5.003544, 4.99537,
  // totalHeight(25,26, 0-49)
    4.987865, 4.9886, 4.988998, 4.98912, 4.989028, 4.98876, 4.988358, 
    4.987854, 4.987276, 4.986655, 4.986023, 4.985425, 4.98491, 4.984558, 
    4.98447, 30, 4.947531, 4.949038, 4.951124, 4.95332, 4.955368, 4.952527, 
    4.950438, 4.948456, 4.947687, 4.948007, 4.94954, 4.952215, 4.956279, 
    4.960855, 4.966729, 4.968522, 4.970867, 4.97377, 4.97719, 4.98108, 
    4.985371, 4.989972, 4.994764, 4.999599, 5.004291, 5.008625, 5.01235, 
    5.015193, 5.01685, 5.017016, 5.015405, 5.011773, 5.005966, 4.997958,
  // totalHeight(25,27, 0-49)
    4.990288, 4.990781, 4.990932, 4.990807, 4.990461, 4.989943, 4.989286, 
    4.988528, 4.987698, 4.986828, 4.985954, 4.985124, 4.984395, 4.983844, 
    4.983571, 30, 4.947104, 4.948366, 4.950164, 4.952053, 4.953806, 4.951047, 
    4.949018, 4.947112, 4.946393, 4.946748, 4.948308, 4.951011, 4.9551, 
    4.959718, 4.965595, 4.967705, 4.970366, 4.973579, 4.977294, 4.981462, 
    4.986007, 4.990837, 4.995832, 5.000842, 5.005686, 5.010149, 5.013985, 
    5.016919, 5.018657, 5.018899, 5.017364, 5.013811, 5.008099, 5.000204,
  // totalHeight(25,28, 0-49)
    4.992364, 4.99267, 4.992622, 4.992288, 4.991722, 4.990971, 4.990073, 
    4.989061, 4.987968, 4.986831, 4.985691, 4.984602, 4.983626, 4.982843, 
    4.982348, 30, 4.947995, 4.94893, 4.950346, 4.951824, 4.953187, 4.950557, 
    4.948601, 4.946773, 4.946075, 4.946415, 4.947931, 4.950579, 4.954597, 
    4.959157, 4.964909, 4.967333, 4.970298, 4.97379, 4.977762, 4.982154, 
    4.986895, 4.991891, 4.997024, 5.002145, 5.00708, 5.011614, 5.015508, 
    5.018489, 5.020265, 5.020542, 5.019038, 5.015524, 5.009858, 5.002028,
  // totalHeight(25,29, 0-49)
    4.99406, 4.994244, 4.994057, 4.993563, 4.992815, 4.991854, 4.990718, 
    4.989445, 4.98807, 4.986638, 4.985197, 4.983812, 4.982553, 4.981504, 
    4.980756, 30, 4.950003, 4.95055, 4.951498, 4.952468, 4.953333, 4.950801, 
    4.948859, 4.947036, 4.946271, 4.946498, 4.947872, 4.950364, 4.954204, 
    4.958596, 4.964083, 4.966768, 4.969983, 4.973703, 4.97788, 4.982456, 
    4.98736, 4.992499, 4.997761, 5.002997, 5.008034, 5.012661, 5.016634, 
    5.019682, 5.021515, 5.021831, 5.020354, 5.016856, 5.011202, 5.003389,
  // totalHeight(25,30, 0-49)
    4.994519, 4.993861, 4.992861, 4.991597, 4.990131, 4.988516, 4.986785, 
    4.984964, 4.983063, 4.981089, 4.979038, 4.976903, 4.974685, 4.97239, 
    4.970056, 4.968032, 4.954024, 4.95362, 4.953893, 4.954456, 4.955149, 
    4.953227, 4.951905, 4.950692, 4.950378, 4.950848, 4.952226, 4.954489, 
    4.957869, 4.961644, 4.966294, 4.968657, 4.97154, 4.974941, 4.978828, 
    4.983158, 4.987868, 4.99287, 4.998047, 5.00325, 5.008296, 5.012966, 
    5.017006, 5.020132, 5.02204, 5.022424, 5.021001, 5.017544, 5.01192, 
    5.004138,
  // totalHeight(25,31, 0-49)
    4.995345, 4.994719, 4.99372, 4.992418, 4.990875, 4.98914, 4.98725, 
    4.985236, 4.983119, 4.98091, 4.978617, 4.976248, 4.9738, 4.97128, 
    4.968707, 4.967444, 4.954495, 4.953582, 4.953315, 4.953332, 4.953514, 
    4.951689, 4.950369, 4.949167, 4.948839, 4.949316, 4.950732, 4.953062, 
    4.956487, 4.960275, 4.964766, 4.967505, 4.970757, 4.974515, 4.978742, 
    4.983388, 4.988389, 4.993653, 4.999059, 5.004455, 5.009655, 5.014433, 
    5.018531, 5.02166, 5.023511, 5.023779, 5.022181, 5.018497, 5.012614, 
    5.004563,
  // totalHeight(25,32, 0-49)
    4.995613, 4.995025, 4.99404, 4.992726, 4.991141, 4.989335, 4.987347, 
    4.985208, 4.982944, 4.980573, 4.978112, 4.975571, 4.972955, 4.970267, 
    4.967512, 4.966613, 4.954969, 4.953597, 4.952828, 4.952345, 4.952063, 
    4.950393, 4.949138, 4.948009, 4.947721, 4.948237, 4.949703, 4.952083, 
    4.955504, 4.959243, 4.96351, 4.966569, 4.97013, 4.97418, 4.978678, 
    4.983575, 4.988803, 4.994267, 4.999846, 5.005381, 5.010685, 5.015527, 
    5.019639, 5.022727, 5.024477, 5.024584, 5.022766, 5.018817, 5.01264, 
    5.00429,
  // totalHeight(25,33, 0-49)
    4.995334, 4.994799, 4.993851, 4.992554, 4.990967, 4.989133, 4.987097, 
    4.984889, 4.982537, 4.980067, 4.977499, 4.97485, 4.972124, 4.969328, 
    4.966456, 4.965581, 4.955402, 4.953644, 4.952435, 4.951514, 4.95083, 
    4.949367, 4.948236, 4.947248, 4.947051, 4.947638, 4.949155, 4.951556, 
    4.954919, 4.958547, 4.962534, 4.96586, 4.96967, 4.973946, 4.978648, 
    4.983727, 4.989114, 4.994714, 5.000402, 5.006021, 5.011372, 5.016219, 
    5.020291, 5.023284, 5.024884, 5.024779, 5.022697, 5.01844, 5.011938, 
    5.003271,
  // totalHeight(25,34, 0-49)
    4.994516, 4.994058, 4.993176, 4.991931, 4.990377, 4.98856, 4.986521, 
    4.984294, 4.981909, 4.979394, 4.976773, 4.974064, 4.971285, 4.968438, 
    4.965515, 4.964412, 4.955777, 4.953714, 4.952136, 4.950844, 4.949824, 
    4.94861, 4.947661, 4.946874, 4.946813, 4.947495, 4.949058, 4.95145, 
    4.954698, 4.95816, 4.961833, 4.965373, 4.969373, 4.97381, 4.978651, 
    4.983845, 4.989325, 4.994994, 5.000727, 5.006361, 5.011694, 5.016483, 
    5.020451, 5.02329, 5.024677, 5.024305, 5.02191, 5.017309, 5.010454, 
    5.001464,
  // totalHeight(25,35, 0-49)
    4.993182, 4.992826, 4.992038, 4.990879, 4.989397, 4.987638, 4.985642, 
    4.983441, 4.98107, 4.978556, 4.975928, 4.97321, 4.970424, 4.967576, 
    4.96466, 4.963175, 4.9561, 4.953816, 4.951942, 4.95035, 4.949063, 
    4.948124, 4.947401, 4.946869, 4.946983, 4.94778, 4.949381, 4.95173, 
    4.954807, 4.958058, 4.961395, 4.965098, 4.969231, 4.97377, 4.978685, 
    4.983928, 4.989433, 4.995101, 5.000806, 5.006383, 5.011625, 5.016284, 
    5.020075, 5.022686, 5.023796, 5.023099, 5.02034, 5.015363, 5.008144, 
    4.998838,
  // totalHeight(25,36, 0-49)
    4.99136, 4.991127, 4.990465, 4.989424, 4.988052, 4.986389, 4.984475, 
    4.982344, 4.980028, 4.97756, 4.974968, 4.972284, 4.969531, 4.966724, 
    4.963866, 4.961936, 4.956396, 4.953965, 4.951863, 4.950037, 4.948545, 
    4.947903, 4.94744, 4.947205, 4.947526, 4.948452, 4.950078, 4.95235, 
    4.955209, 4.958213, 4.961207, 4.965024, 4.969234, 4.973816, 4.978744, 
    4.983969, 4.989426, 4.995021, 5.000623, 5.006064, 5.011133, 5.01558, 
    5.019113, 5.02142, 5.022179, 5.021094, 5.017928, 5.012548, 5.004965, 
    4.995371,
  // totalHeight(25,37, 0-49)
    4.989093, 4.989005, 4.988489, 4.987594, 4.986362, 4.984831, 4.983038, 
    4.981017, 4.9788, 4.976418, 4.973905, 4.97129, 4.968606, 4.965876, 
    4.963112, 4.960749, 4.956685, 4.954175, 4.951907, 4.949906, 4.948266, 
    4.947929, 4.947752, 4.947848, 4.9484, 4.949461, 4.951101, 4.953265, 
    4.955864, 4.958595, 4.961247, 4.96513, 4.969367, 4.973936, 4.978812, 
    4.983953, 4.989293, 4.994737, 5.000153, 5.005373, 5.010181, 5.014324, 
    5.01751, 5.019426, 5.01976, 5.018228, 5.014614, 5.008818, 5.000887, 
    4.991054,
  // totalHeight(25,38, 0-49)
    4.986433, 4.986499, 4.986148, 4.985423, 4.98436, 4.982993, 4.981357, 
    4.979482, 4.977402, 4.975144, 4.972745, 4.970237, 4.967655, 4.965031, 
    4.962386, 4.959657, 4.956991, 4.954454, 4.952072, 4.949954, 4.948216, 
    4.948183, 4.948303, 4.948752, 4.949552, 4.950753, 4.952391, 4.954421, 
    4.956728, 4.959168, 4.961491, 4.965396, 4.969607, 4.974107, 4.978873, 
    4.983865, 4.989013, 4.994225, 4.999371, 5.004277, 5.008728, 5.012469, 
    5.015213, 5.016651, 5.016483, 5.014445, 5.010352, 5.00414, 4.995898, 
    4.985897,
  // totalHeight(25,39, 0-49)
    4.98344, 4.983667, 4.983495, 4.982955, 4.982084, 4.980909, 4.979459, 
    4.977764, 4.975853, 4.973757, 4.971507, 4.969138, 4.966689, 4.964193, 
    4.961687, 4.95869, 4.957332, 4.954806, 4.952355, 4.950166, 4.948378, 
    4.948637, 4.949059, 4.949871, 4.950925, 4.952264, 4.953889, 4.955763, 
    4.957753, 4.959896, 4.961904, 4.965787, 4.969928, 4.974308, 4.978906, 
    4.983677, 4.988561, 4.99346, 4.998243, 5.002738, 5.006731, 5.009968, 
    5.01217, 5.013039, 5.012294, 5.0097, 5.00511, 4.998499, 4.990002, 4.97993,
  // totalHeight(25,40, 0-49)
    4.980185, 4.980569, 4.980579, 4.980239, 4.979576, 4.978613, 4.977376, 
    4.975892, 4.974182, 4.972278, 4.970209, 4.96801, 4.96572, 4.963377, 
    4.961021, 4.957868, 4.957716, 4.955232, 4.952751, 4.950531, 4.948729, 
    4.949263, 4.949982, 4.951154, 4.952459, 4.953933, 4.955529, 4.957229, 
    4.95889, 4.960732, 4.962445, 4.966266, 4.970292, 4.974501, 4.978872, 
    4.983361, 4.987904, 4.992404, 4.996732, 5.000714, 5.004144, 5.006771, 
    5.008329, 5.008542, 5.007154, 5.003967, 4.998874, 4.9919, 4.983227, 
    4.973203,
  // totalHeight(25,41, 0-49)
    4.976741, 4.977275, 4.977466, 4.97733, 4.976886, 4.976152, 4.975149, 
    4.973896, 4.972416, 4.970734, 4.968876, 4.966875, 4.964769, 4.962596, 
    4.960401, 4.957204, 4.958153, 4.95573, 4.953249, 4.951032, 4.949247, 
    4.950036, 4.951032, 4.952551, 4.954097, 4.955692, 4.957246, 4.958759, 
    4.960083, 4.96163, 4.963066, 4.966787, 4.970655, 4.974645, 4.978733, 
    4.982875, 4.987002, 4.991017, 4.994792, 4.998161, 5.000918, 5.00283, 
    5.003649, 5.003125, 5.001037, 4.997231, 4.991654, 4.984376, 4.975628, 
    4.965791,
  // totalHeight(25,42, 0-49)
    4.973186, 4.973859, 4.974224, 4.97429, 4.974071, 4.973577, 4.972821, 
    4.971821, 4.970592, 4.969154, 4.967532, 4.965755, 4.963854, 4.96187, 
    4.959843, 4.956702, 4.958642, 4.956295, 4.953839, 4.951653, 4.949909, 
    4.950922, 4.952172, 4.954015, 4.955778, 4.957478, 4.958976, 4.96029, 
    4.961278, 4.962534, 4.963706, 4.967291, 4.970962, 4.974685, 4.978436, 
    4.982165, 4.985803, 4.989247, 4.992375, 4.995026, 4.997008, 4.998106, 
    4.998096, 4.996766, 4.993938, 4.989511, 4.983484, 4.975986, 4.967286, 
    4.957791,
  // totalHeight(25,43, 0-49)
    4.969604, 4.970394, 4.970921, 4.971184, 4.971187, 4.970936, 4.970438, 
    4.969702, 4.968741, 4.967569, 4.966205, 4.964672, 4.962998, 4.961216, 
    4.959366, 4.956364, 4.959184, 4.95692, 4.954512, 4.952376, 4.950689, 
    4.951897, 4.953369, 4.955495, 4.957449, 4.959227, 4.960651, 4.961758, 
    4.962413, 4.963387, 4.964305, 4.967716, 4.971148, 4.97456, 4.977921, 
    4.981175, 4.984247, 4.987039, 4.989427, 4.991263, 4.992372, 4.992564, 
    4.99165, 4.989461, 4.985876, 4.980847, 4.974436, 4.966821, 4.958312, 
    4.949332,
  // totalHeight(25,44, 0-49)
    4.966064, 4.966953, 4.967626, 4.968073, 4.968293, 4.968284, 4.968047, 
    4.967584, 4.966902, 4.966008, 4.964917, 4.963645, 4.962215, 4.960651, 
    4.958984, 4.956183, 4.95977, 4.9576, 4.955254, 4.953185, 4.951562, 
    4.952929, 4.954587, 4.956951, 4.959055, 4.960881, 4.962212, 4.963103, 
    4.963431, 4.964125, 4.96479, 4.967986, 4.971137, 4.974195, 4.977112, 
    4.979828, 4.982265, 4.984324, 4.98589, 4.986822, 4.986973, 4.986184, 
    4.984309, 4.981235, 4.976897, 4.971315, 4.964608, 4.957005, 4.948846, 
    4.940559,
  // totalHeight(25,45, 0-49)
    4.962638, 4.963603, 4.964401, 4.965019, 4.965446, 4.965672, 4.965693, 
    4.965505, 4.965105, 4.964497, 4.96369, 4.962691, 4.961516, 4.960183, 
    4.958711, 4.95615, 4.96039, 4.958319, 4.956052, 4.954056, 4.952502, 
    4.953992, 4.955791, 4.95834, 4.960548, 4.962384, 4.963598, 4.964264, 
    4.96427, 4.96468, 4.965085, 4.968025, 4.97085, 4.973502, 4.975922, 
    4.978043, 4.97978, 4.981034, 4.9817, 4.981656, 4.98078, 4.978958, 
    4.976094, 4.972135, 4.967084, 4.961026, 4.954139, 4.946698, 4.939058, 
    4.931637,
  // totalHeight(25,46, 0-49)
    4.959384, 4.960401, 4.961304, 4.962074, 4.962692, 4.963142, 4.963412, 
    4.963494, 4.963376, 4.963057, 4.962538, 4.961819, 4.96091, 4.959814, 
    4.958544, 4.956244, 4.961024, 4.959065, 4.956888, 4.954971, 4.95348, 
    4.955057, 4.95695, 4.959622, 4.961882, 4.963686, 4.964756, 4.965185, 
    4.964869, 4.964985, 4.965108, 4.967745, 4.970198, 4.972394, 4.974265, 
    4.975734, 4.97671, 4.977099, 4.976804, 4.975729, 4.973786, 4.970906, 
    4.967056, 4.962245, 4.956552, 4.950125, 4.9432, 4.936079, 4.92913, 
    4.922746,
  // totalHeight(25,47, 0-49)
    4.95635, 4.957393, 4.95838, 4.959281, 4.960072, 4.960729, 4.961237, 
    4.961576, 4.961733, 4.961699, 4.961466, 4.961028, 4.960386, 4.959536, 
    4.958477, 4.956443, 4.961648, 4.959813, 4.957735, 4.955901, 4.954465, 
    4.956092, 4.958033, 4.960762, 4.963014, 4.964739, 4.965635, 4.965809, 
    4.965172, 4.964973, 4.964783, 4.967062, 4.969089, 4.970776, 4.972046, 
    4.972809, 4.972975, 4.972452, 4.971157, 4.969021, 4.966, 4.962074, 
    4.957274, 4.951685, 4.945455, 4.938794, 4.931985, 4.925356, 4.919264, 
    4.914069,
  // totalHeight(25,48, 0-49)
    4.953563, 4.954612, 4.955658, 4.956668, 4.957611, 4.958456, 4.959181, 
    4.959764, 4.960183, 4.96042, 4.960465, 4.960305, 4.959929, 4.959326, 
    4.958488, 4.956709, 4.96223, 4.960528, 4.958559, 4.956808, 4.955421, 
    4.957064, 4.959004, 4.961722, 4.963907, 4.965501, 4.966192, 4.966093, 
    4.965123, 4.964581, 4.964033, 4.965894, 4.967434, 4.968557, 4.969174, 
    4.969187, 4.968502, 4.967037, 4.964726, 4.961534, 4.957456, 4.952534, 
    4.946867, 4.940608, 4.933976, 4.927238, 4.920715, 4.914744, 4.909664, 
    4.90578,
  // totalHeight(25,49, 0-49)
    4.95051, 4.9514, 4.952364, 4.953356, 4.954337, 4.95527, 4.956123, 
    4.956862, 4.957456, 4.957881, 4.95811, 4.958118, 4.957881, 4.957365, 
    4.956535, 4.954092, 4.966395, 4.963832, 4.960638, 4.957756, 4.955451, 
    4.959006, 4.962871, 4.96796, 4.971593, 4.973686, 4.973638, 4.971708, 
    4.96775, 4.964478, 4.961112, 4.962604, 4.963628, 4.964084, 4.963889, 
    4.962953, 4.961198, 4.958563, 4.95502, 4.950583, 4.945317, 4.939349, 
    4.932869, 4.926122, 4.919407, 4.91305, 4.907397, 4.902774, 4.899466, 
    4.897687,
  // totalHeight(26,0, 0-49)
    4.94, 4.944391, 4.94844, 4.952157, 4.95555, 4.958627, 4.961393, 4.963849, 
    4.965998, 4.96784, 4.969378, 4.970623, 4.97159, 4.972304, 4.9728, 
    4.972906, 4.973375, 4.973431, 4.973461, 4.973564, 4.973804, 4.974427, 
    4.975248, 4.976345, 4.977716, 4.979355, 4.981232, 4.983315, 4.985551, 
    4.987894, 4.990223, 4.992686, 4.994967, 4.996955, 4.998531, 4.999562, 
    4.999901, 4.999391, 4.997859, 4.995126, 4.991014, 4.985359, 4.978026, 
    4.968945, 4.958121, 4.945682, 4.931883, 4.917126, 4.901945, 4.886976,
  // totalHeight(26,1, 0-49)
    4.941255, 4.945621, 4.949628, 4.95329, 4.956614, 4.959611, 4.962287, 
    4.96465, 4.966698, 4.96844, 4.96988, 4.971029, 4.971907, 4.972544, 
    4.972975, 4.97282, 4.973508, 4.973464, 4.973378, 4.973377, 4.973534, 
    4.974285, 4.975206, 4.976415, 4.977892, 4.979619, 4.981553, 4.983666, 
    4.985904, 4.988244, 4.990533, 4.993175, 4.995648, 4.997859, 4.999695, 
    5.00104, 5.001753, 5.001679, 5.000646, 4.998471, 4.994966, 4.989946, 
    4.983253, 4.97478, 4.964502, 4.952498, 4.938988, 4.924335, 4.909052, 
    4.893767,
  // totalHeight(26,2, 0-49)
    4.942569, 4.946893, 4.950846, 4.954443, 4.957692, 4.960606, 4.963196, 
    4.965467, 4.967426, 4.969079, 4.970437, 4.971511, 4.972326, 4.97291, 
    4.973302, 4.972916, 4.973806, 4.973686, 4.973504, 4.973412, 4.973489, 
    4.974351, 4.975346, 4.976624, 4.978158, 4.979918, 4.981861, 4.983953, 
    4.986146, 4.988422, 4.990607, 4.993344, 4.995931, 4.998283, 5.000306, 
    5.001887, 5.002901, 5.0032, 5.002613, 5.00096, 4.998045, 4.993671, 
    4.987662, 4.979883, 4.970272, 4.958864, 4.945834, 4.931497, 4.916326, 
    4.900925,
  // totalHeight(26,3, 0-49)
    4.943935, 4.948204, 4.952092, 4.955615, 4.958785, 4.961618, 4.964122, 
    4.966311, 4.968189, 4.969768, 4.97106, 4.97208, 4.972853, 4.973409, 
    4.973786, 4.973205, 4.974256, 4.974084, 4.97383, 4.973662, 4.973668, 
    4.974619, 4.975657, 4.976962, 4.978502, 4.98025, 4.982156, 4.984193, 
    4.986302, 4.988472, 4.990499, 4.99326, 4.995889, 4.99831, 5.000443, 
    5.002193, 5.003439, 5.004045, 5.003849, 5.002671, 5.000317, 4.996583, 
    4.991277, 4.984245, 4.975389, 4.964705, 4.952313, 4.938476, 4.923614, 
    4.908288,
  // totalHeight(26,4, 0-49)
    4.945349, 4.949549, 4.953363, 4.956806, 4.959896, 4.962646, 4.96507, 
    4.967181, 4.96899, 4.970509, 4.97175, 4.972735, 4.973485, 4.974032, 
    4.974418, 4.973681, 4.974834, 4.974633, 4.974329, 4.974107, 4.97405, 
    4.975069, 4.976121, 4.977407, 4.978909, 4.980601, 4.982437, 4.984389, 
    4.986394, 4.988424, 4.990258, 4.992982, 4.995586, 4.998013, 5.000195, 
    5.002046, 5.003461, 5.004312, 5.004447, 5.003695, 5.001862, 4.998744, 
    4.994145, 4.987888, 4.979846, 4.969979, 4.958351, 4.945166, 4.930783, 
    4.915707,
  // totalHeight(26,5, 0-49)
    4.946802, 4.950924, 4.954657, 4.958016, 4.961022, 4.96369, 4.966037, 
    4.968078, 4.969824, 4.971294, 4.9725, 4.973464, 4.974208, 4.974766, 
    4.975174, 4.974328, 4.975505, 4.975296, 4.974972, 4.974713, 4.974607, 
    4.97567, 4.976707, 4.977932, 4.979356, 4.980954, 4.982691, 4.984538, 
    4.986431, 4.988306, 4.989924, 4.992555, 4.995082, 4.997459, 4.999632, 
    5.001528, 5.003053, 5.004092, 5.004505, 5.004128, 5.002773, 5.000243, 
    4.996334, 4.99086, 4.983668, 4.974679, 4.963905, 4.951492, 4.937729, 
    4.923054,
  // totalHeight(26,6, 0-49)
    4.948296, 4.952331, 4.955975, 4.959248, 4.962167, 4.964754, 4.967025, 
    4.969, 4.97069, 4.972117, 4.973296, 4.974251, 4.975002, 4.975583, 
    4.976024, 4.975116, 4.97623, 4.976032, 4.975711, 4.975441, 4.975303, 
    4.976385, 4.977377, 4.978502, 4.979811, 4.981283, 4.982903, 4.984636, 
    4.986417, 4.988131, 4.989528, 4.992019, 4.994424, 4.996704, 4.998821, 
    5.000714, 5.002299, 5.003477, 5.004117, 5.004066, 5.00315, 5.001173, 
    4.997931, 4.99323, 4.986898, 4.978821, 4.968964, 4.957409, 4.944374, 
    4.930231,
  // totalHeight(26,7, 0-49)
    4.949835, 4.953774, 4.957324, 4.960505, 4.963335, 4.965837, 4.968033, 
    4.96994, 4.971579, 4.972966, 4.974124, 4.975074, 4.97584, 4.976448, 
    4.976927, 4.976012, 4.976964, 4.976792, 4.976501, 4.976244, 4.976095, 
    4.977169, 4.97809, 4.97908, 4.980241, 4.981565, 4.983052, 4.984669, 
    4.986344, 4.987903, 4.98909, 4.991405, 4.993648, 4.995795, 4.997818, 
    4.999667, 5.001273, 5.002547, 5.003373, 5.003607, 5.003088, 5.001628, 
    4.999024, 4.995079, 4.989602, 4.982448, 4.97354, 4.962898, 4.950672, 
    4.93716,
  // totalHeight(26,8, 0-49)
    4.951429, 4.955265, 4.958713, 4.961794, 4.96453, 4.966943, 4.969059, 
    4.970898, 4.97248, 4.97383, 4.974967, 4.975914, 4.976696, 4.977333, 
    4.977845, 4.976974, 4.97766, 4.977527, 4.977291, 4.977073, 4.976935, 
    4.977974, 4.978799, 4.979623, 4.980614, 4.98177, 4.983119, 4.98462, 
    4.986207, 4.987626, 4.988623, 4.99073, 4.992783, 4.994769, 4.996668, 
    4.998445, 5.000041, 5.001379, 5.002355, 5.002841, 5.002684, 5.001705, 
    4.99971, 4.99649, 4.991849, 4.985611, 4.97766, 4.967961, 4.956597, 
    4.943792,
  // totalHeight(26,9, 0-49)
    4.953088, 4.956812, 4.96015, 4.963123, 4.965757, 4.968074, 4.970102, 
    4.971866, 4.973389, 4.974695, 4.975805, 4.976745, 4.977537, 4.978196, 
    4.978734, 4.97796, 4.97827, 4.978189, 4.978033, 4.97788, 4.97778, 
    4.978755, 4.97946, 4.980095, 4.980895, 4.981874, 4.98308, 4.984471, 
    4.985987, 4.987292, 4.988131, 4.990008, 4.991851, 4.993655, 4.995411, 
    4.997094, 4.998659, 5.000037, 5.00114, 5.001849, 5.002026, 5.001497, 
    5.000074, 4.99755, 4.993714, 4.988372, 4.981369, 4.972619, 4.962144, 
    4.950095,
  // totalHeight(26,10, 0-49)
    4.954827, 4.958428, 4.961646, 4.964502, 4.967022, 4.969234, 4.971165, 
    4.972841, 4.974293, 4.975544, 4.97662, 4.977544, 4.978334, 4.979006, 
    4.979555, 4.97893, 4.97875, 4.978733, 4.978679, 4.978618, 4.978583, 
    4.979466, 4.980032, 4.980456, 4.981056, 4.981851, 4.982915, 4.984207, 
    4.985671, 4.986889, 4.987614, 4.989247, 4.990867, 4.992477, 4.99408, 
    4.995658, 4.997178, 4.998582, 4.999794, 5.000707, 5.001192, 5.001086, 
    5.000204, 4.998339, 4.995272, 4.990792, 4.98471, 4.976898, 4.967317, 
    4.956054,
  // totalHeight(26,11, 0-49)
    4.956657, 4.960123, 4.963208, 4.965933, 4.968327, 4.970419, 4.972239, 
    4.973818, 4.975185, 4.976367, 4.977395, 4.978288, 4.979064, 4.97973, 
    4.980277, 4.979839, 4.979058, 4.979119, 4.979188, 4.979247, 4.979304, 
    4.980065, 4.980476, 4.980678, 4.981071, 4.981682, 4.982608, 4.983808, 
    4.985242, 4.986406, 4.987069, 4.98845, 4.989841, 4.991255, 4.992701, 
    4.994172, 4.995643, 4.997068, 4.998378, 4.99948, 5.000252, 5.000543, 
    5.00017, 4.998927, 4.996589, 4.992929, 4.987732, 4.98083, 4.972133, 
    4.961664,
  // totalHeight(26,12, 0-49)
    4.958586, 4.961901, 4.964838, 4.967417, 4.96967, 4.971628, 4.973322, 
    4.974786, 4.976053, 4.977152, 4.978113, 4.978957, 4.9797, 4.980344, 
    4.98087, 4.980648, 4.979154, 4.979307, 4.979526, 4.97973, 4.979906, 
    4.980518, 4.980759, 4.980734, 4.980921, 4.981354, 4.982149, 4.983266, 
    4.984689, 4.985831, 4.986491, 4.987618, 4.988783, 4.990006, 4.9913, 
    4.992667, 4.994092, 4.995536, 4.996943, 4.998224, 4.99927, 4.999934, 
    5.000038, 4.999378, 4.997725, 4.994837, 4.990478, 4.984446, 4.976607, 
    4.966925,
  // totalHeight(26,13, 0-49)
    4.960617, 4.963764, 4.966533, 4.968949, 4.971044, 4.97285, 4.974402, 
    4.975734, 4.976882, 4.97788, 4.978757, 4.979533, 4.980224, 4.980828, 
    4.981322, 4.981328, 4.979001, 4.979272, 4.979662, 4.980037, 4.98036, 
    4.980793, 4.980856, 4.980605, 4.980595, 4.980857, 4.981531, 4.982577, 
    4.984003, 4.985156, 4.985874, 4.986757, 4.987704, 4.988744, 4.989898, 
    4.991172, 4.992559, 4.994028, 4.99553, 4.996988, 4.998293, 4.999307, 
    4.999858, 4.999741, 4.998724, 4.996556, 4.992984, 4.987775, 4.980757, 
    4.971845,
  // totalHeight(26,14, 0-49)
    4.962743, 4.965701, 4.968283, 4.970517, 4.972435, 4.974072, 4.975463, 
    4.976647, 4.977662, 4.978541, 4.979313, 4.980003, 4.980623, 4.981172, 
    4.981625, 4.981853, 4.978575, 4.978984, 4.97957, 4.980143, 4.980638, 
    4.980866, 4.980747, 4.980277, 4.980084, 4.980192, 4.980755, 4.98174, 
    4.983183, 4.984377, 4.985216, 4.985863, 4.986608, 4.987482, 4.988513, 
    4.989711, 4.991073, 4.992577, 4.994179, 4.995807, 4.99736, 4.998702, 
    4.999669, 5.000055, 4.999626, 4.998124, 4.995279, 4.99084, 4.984598, 
    4.976427,
  // totalHeight(26,15, 0-49)
    4.96495, 4.967693, 4.970068, 4.972099, 4.973822, 4.975271, 4.976488, 
    4.977509, 4.978373, 4.979118, 4.979771, 4.980357, 4.980891, 4.98137, 
    4.981779, 4.982203, 4.977856, 4.978431, 4.979234, 4.980026, 4.980718, 
    4.98072, 4.98042, 4.979746, 4.97939, 4.979363, 4.979831, 4.980763, 
    4.982235, 4.983498, 4.984517, 4.984947, 4.985507, 4.986237, 4.987163, 
    4.988302, 4.989655, 4.991206, 4.992913, 4.99471, 4.996499, 4.998151, 
    4.999502, 5.000349, 5.000455, 4.999561, 4.997384, 4.993657, 4.98814, 
    4.980677,
  // totalHeight(26,16, 0-49)
    4.967216, 4.969719, 4.971859, 4.973665, 4.975173, 4.97642, 4.977448, 
    4.978295, 4.979, 4.979597, 4.98012, 4.98059, 4.981026, 4.981429, 4.98179, 
    4.98237, 4.976842, 4.977604, 4.978645, 4.979676, 4.980588, 4.980343, 
    4.979868, 4.979012, 4.978518, 4.978383, 4.978773, 4.979663, 4.981173, 
    4.982527, 4.983779, 4.984013, 4.984412, 4.98502, 4.985863, 4.986963, 
    4.988326, 4.989933, 4.991749, 4.993711, 4.995725, 4.997665, 4.999369, 
    5.000635, 5.001229, 5.000884, 4.999315, 4.996238, 4.991397, 4.984601,
  // totalHeight(26,17, 0-49)
    4.969512, 4.97174, 4.973618, 4.975176, 4.976452, 4.977484, 4.978314, 
    4.97898, 4.979518, 4.979966, 4.980352, 4.980701, 4.981031, 4.981352, 
    4.981671, 4.982362, 4.975548, 4.976512, 4.977801, 4.979086, 4.980233, 
    4.979731, 4.979088, 4.978076, 4.977477, 4.977263, 4.977597, 4.978462, 
    4.980017, 4.981482, 4.98301, 4.983071, 4.983333, 4.983841, 4.984626, 
    4.985706, 4.987091, 4.988766, 4.990695, 4.99282, 4.995048, 4.997253, 
    4.999278, 5.000922, 5.001952, 5.002101, 5.001079, 4.998593, 4.994374, 
    4.988206,
  // totalHeight(26,18, 0-49)
    4.971802, 4.973717, 4.975297, 4.976582, 4.977609, 4.978417, 4.979047, 
    4.979535, 4.979914, 4.980217, 4.98047, 4.980698, 4.980921, 4.981159, 
    4.981435, 4.982197, 4.974019, 4.975191, 4.976727, 4.978267, 4.979657, 
    4.978886, 4.978089, 4.97695, 4.976281, 4.976023, 4.97633, 4.977189, 
    4.978799, 4.980386, 4.982221, 4.982135, 4.982282, 4.982712, 4.983455, 
    4.984532, 4.985951, 4.9877, 4.989746, 4.992026, 4.994454, 4.996904, 
    4.999218, 5.001203, 5.002622, 5.003211, 5.00268, 5.00073, 4.99708, 
    4.991498,
  // totalHeight(26,19, 0-49)
    4.974044, 4.975593, 4.976839, 4.977823, 4.978588, 4.979169, 4.979604, 
    4.979926, 4.980161, 4.980335, 4.98047, 4.980588, 4.98071, 4.980864, 
    4.981096, 4.981905, 4.972337, 4.973706, 4.975469, 4.977249, 4.978876, 
    4.977831, 4.976893, 4.975658, 4.974956, 4.974691, 4.975004, 4.975879, 
    4.977556, 4.979274, 4.981433, 4.981222, 4.981273, 4.981641, 4.982354, 
    4.983438, 4.984897, 4.986722, 4.98888, 4.991309, 4.993922, 4.996593, 
    4.999171, 5.001457, 5.003224, 5.004207, 5.004115, 5.00265, 4.999523, 
    4.994492,
  // totalHeight(26,20, 0-49)
    4.977043, 4.979004, 4.980653, 4.982024, 4.983145, 4.984046, 4.984755, 
    4.985302, 4.985719, 4.986032, 4.986275, 4.986479, 4.986677, 4.986904, 
    4.987205, 30, 4.969875, 4.971127, 4.972816, 4.974531, 4.976083, 4.974407, 
    4.972915, 4.971169, 4.97008, 4.969584, 4.969836, 4.970838, 4.972848, 
    4.975082, 4.978014, 4.978158, 4.978577, 4.979314, 4.980385, 4.981804, 
    4.983576, 4.985689, 4.988112, 4.990792, 4.993645, 4.996556, 4.999379, 
    5.001928, 5.003983, 5.005283, 5.005549, 5.004485, 5.001798, 4.997241,
  // totalHeight(26,21, 0-49)
    4.97925, 4.980883, 4.98223, 4.983332, 4.984216, 4.984912, 4.985448, 
    4.985849, 4.986141, 4.98635, 4.9865, 4.986621, 4.986745, 4.986916, 
    4.987184, 30, 4.965111, 4.966493, 4.968369, 4.970301, 4.97207, 4.970103, 
    4.968467, 4.966664, 4.965661, 4.965364, 4.965918, 4.967295, 4.969753, 
    4.972483, 4.976055, 4.976404, 4.977072, 4.978096, 4.979475, 4.981217, 
    4.983313, 4.985742, 4.988464, 4.991421, 4.994527, 4.997666, 5.000692, 
    5.003428, 5.005657, 5.007132, 5.007581, 5.006714, 5.004252, 4.999951,
  // totalHeight(26,22, 0-49)
    4.981404, 4.982722, 4.983783, 4.984627, 4.985284, 4.985783, 4.986148, 
    4.986403, 4.986568, 4.986663, 4.986715, 4.986749, 4.986797, 4.986908, 
    4.98714, 30, 4.96099, 4.962482, 4.964514, 4.966624, 4.968567, 4.966304, 
    4.964496, 4.962591, 4.961608, 4.961434, 4.962199, 4.963859, 4.966667, 
    4.969792, 4.973887, 4.974385, 4.975251, 4.976512, 4.978163, 4.980196, 
    4.982597, 4.985335, 4.988364, 4.991613, 4.994995, 4.998389, 5.00165, 
    5.004604, 5.007035, 5.008707, 5.009351, 5.008693, 5.006459, 5.002415,
  // totalHeight(26,23, 0-49)
    4.983479, 4.984495, 4.985284, 4.985883, 4.986323, 4.986632, 4.986832, 
    4.98694, 4.986977, 4.986959, 4.986909, 4.98685, 4.986816, 4.986859, 
    4.987047, 30, 4.957404, 4.958957, 4.961073, 4.96328, 4.965307, 4.962757, 
    4.96076, 4.958724, 4.957712, 4.957599, 4.958509, 4.960382, 4.963464, 
    4.966908, 4.971419, 4.972058, 4.973106, 4.974591, 4.9765, 4.978821, 
    4.981529, 4.984586, 4.987936, 4.991505, 4.995192, 4.998876, 5.002409, 
    5.00561, 5.008269, 5.010154, 5.011004, 5.010548, 5.008529, 5.004719,
  // totalHeight(26,24, 0-49)
    4.985459, 4.986189, 4.98672, 4.987087, 4.98732, 4.987445, 4.987481, 
    4.987444, 4.987351, 4.987216, 4.987059, 4.986901, 4.986779, 4.986742, 
    4.986866, 30, 4.954684, 4.956232, 4.958356, 4.960571, 4.962602, 4.959841, 
    4.957701, 4.955566, 4.954525, 4.954449, 4.955456, 4.957479, 4.960763, 
    4.964447, 4.969274, 4.970074, 4.971316, 4.973023, 4.975178, 4.977761, 
    4.980742, 4.984078, 4.98771, 4.991553, 4.995505, 4.999441, 5.003209, 
    5.006629, 5.009492, 5.011566, 5.012599, 5.012326, 5.010496, 5.006893,
  // totalHeight(26,25, 0-49)
    4.987332, 4.987795, 4.988081, 4.988227, 4.98826, 4.988207, 4.988082, 
    4.987899, 4.987672, 4.987413, 4.98714, 4.986873, 4.986648, 4.986516, 
    4.986553, 30, 4.952617, 4.954093, 4.956138, 4.958269, 4.960216, 4.957344, 
    4.955132, 4.95296, 4.95192, 4.951881, 4.952963, 4.955096, 4.958523, 
    4.962382, 4.96742, 4.968424, 4.96989, 4.971837, 4.974241, 4.977078, 
    4.980317, 4.983906, 4.987782, 4.991862, 4.996039, 5.000186, 5.004151, 
    5.007753, 5.010787, 5.013021, 5.014207, 5.014087, 5.012415, 5.008984,
  // totalHeight(26,26, 0-49)
    4.989085, 4.989303, 4.989362, 4.989299, 4.989142, 4.988912, 4.988623, 
    4.988289, 4.987917, 4.98752, 4.987116, 4.986723, 4.986379, 4.986131, 
    4.986053, 30, 4.951242, 4.952576, 4.954455, 4.95641, 4.958189, 4.955317, 
    4.953111, 4.950973, 4.949968, 4.949975, 4.951116, 4.953321, 4.956832, 
    4.960795, 4.965936, 4.967187, 4.96891, 4.971114, 4.973774, 4.976858, 
    4.980333, 4.984146, 4.988233, 4.992505, 4.996861, 5.001172, 5.005288, 
    5.009029, 5.012194, 5.014551, 5.015856, 5.015856, 5.014309, 5.011011,
  // totalHeight(26,27, 0-49)
    4.990705, 4.990705, 4.990558, 4.990302, 4.989961, 4.989553, 4.989096, 
    4.988595, 4.988062, 4.987507, 4.986948, 4.986408, 4.985921, 4.985535, 
    4.985317, 30, 4.950675, 4.9518, 4.953434, 4.955128, 4.956655, 4.953875, 
    4.951737, 4.949679, 4.948724, 4.948766, 4.949928, 4.952152, 4.955673, 
    4.959657, 4.964782, 4.966302, 4.968293, 4.970756, 4.97366, 4.976973, 
    4.980659, 4.984664, 4.988923, 4.993354, 4.997853, 5.002294, 5.00653, 
    5.010384, 5.013654, 5.016113, 5.017517, 5.017615, 5.016166, 5.012967,
  // totalHeight(26,28, 0-49)
    4.992178, 4.991997, 4.991673, 4.991239, 4.990721, 4.990136, 4.989495, 
    4.988809, 4.988087, 4.987344, 4.9866, 4.985881, 4.985225, 4.984678, 
    4.984301, 30, 4.951277, 4.95214, 4.953459, 4.954813, 4.956015, 4.953386, 
    4.95134, 4.949368, 4.948436, 4.948458, 4.949565, 4.951716, 4.955142, 
    4.959041, 4.964017, 4.965793, 4.968029, 4.970719, 4.973828, 4.977328, 
    4.981176, 4.985326, 4.989712, 4.994259, 4.998865, 5.003407, 5.007742, 
    5.011695, 5.015062, 5.017617, 5.019115, 5.019303, 5.017936, 5.014811,
  // totalHeight(26,29, 0-49)
    4.993492, 4.993173, 4.992706, 4.992117, 4.991431, 4.990662, 4.989821, 
    4.98892, 4.987972, 4.987, 4.986029, 4.985097, 4.984242, 4.98352, 
    4.982977, 30, 4.952824, 4.953395, 4.954348, 4.955293, 4.95609, 4.953598, 
    4.951597, 4.949647, 4.948653, 4.948557, 4.949506, 4.951476, 4.95469, 
    4.958384, 4.963066, 4.965036, 4.967458, 4.970321, 4.97359, 4.977238, 
    4.981226, 4.985511, 4.990031, 4.994714, 4.999458, 5.004147, 5.00863, 
    5.012733, 5.016247, 5.018942, 5.020564, 5.020856, 5.019571, 5.016503,
  // totalHeight(26,30, 0-49)
    4.99386, 4.992723, 4.991463, 4.990121, 4.988725, 4.987293, 4.985828, 
    4.984329, 4.982784, 4.98118, 4.979504, 4.977741, 4.975895, 4.973988, 
    4.972077, 4.969747, 4.956999, 4.956827, 4.957161, 4.957656, 4.958186, 
    4.95614, 4.954606, 4.953129, 4.952481, 4.952558, 4.953475, 4.955208, 
    4.957977, 4.961077, 4.964963, 4.966609, 4.968697, 4.971236, 4.974212, 
    4.977611, 4.981407, 4.985562, 4.990018, 4.994699, 4.999503, 5.004301, 
    5.008934, 5.013212, 5.016919, 5.019805, 5.021607, 5.022055, 5.020894, 
    5.017915,
  // totalHeight(26,31, 0-49)
    4.994776, 4.99362, 4.992315, 4.990895, 4.989389, 4.987814, 4.986178, 
    4.984484, 4.982728, 4.980905, 4.979011, 4.977039, 4.974996, 4.972894, 
    4.97077, 4.969105, 4.957089, 4.956472, 4.956341, 4.956375, 4.956476, 
    4.954564, 4.953073, 4.951636, 4.950986, 4.951061, 4.95199, 4.953743, 
    4.956496, 4.959546, 4.963222, 4.965158, 4.96754, 4.970372, 4.973639, 
    4.977323, 4.981398, 4.985823, 4.99054, 4.995468, 5.000506, 5.005515, 
    5.010334, 5.014765, 5.01858, 5.021528, 5.023334, 5.023723, 5.022443, 
    5.01929,
  // totalHeight(26,32, 0-49)
    4.995375, 4.994205, 4.99286, 4.991376, 4.989777, 4.988082, 4.986303, 
    4.984447, 4.982514, 4.980509, 4.978431, 4.976282, 4.974068, 4.971794, 
    4.969482, 4.968209, 4.95724, 4.956205, 4.955632, 4.955235, 4.954943, 
    4.953212, 4.951815, 4.950471, 4.949865, 4.949964, 4.950908, 4.952662, 
    4.955353, 4.958293, 4.961698, 4.963876, 4.966497, 4.969563, 4.973063, 
    4.976978, 4.981282, 4.985934, 4.990874, 4.996023, 5.001267, 5.006473, 
    5.011462, 5.016034, 5.019948, 5.022943, 5.024738, 5.025053, 5.023633, 
    5.020279,
  // totalHeight(26,33, 0-49)
    4.995639, 4.99447, 4.9931, 4.991568, 4.989897, 4.988105, 4.98621, 
    4.984221, 4.982143, 4.979988, 4.97776, 4.975465, 4.973111, 4.970702, 
    4.968242, 4.967098, 4.957392, 4.955994, 4.955024, 4.954244, 4.95361, 
    4.952107, 4.950858, 4.949664, 4.949143, 4.949293, 4.950252, 4.951982, 
    4.954559, 4.957333, 4.960416, 4.962787, 4.965594, 4.96884, 4.972515, 
    4.976605, 4.981087, 4.985918, 4.991039, 4.996368, 5.001789, 5.007158, 
    5.012293, 5.01698, 5.020972, 5.023992, 5.025752, 5.025967, 5.02438, 
    5.020803,
  // totalHeight(26,34, 0-49)
    4.995543, 4.994396, 4.993027, 4.99147, 4.98975, 4.98789, 4.985905, 
    4.983811, 4.98162, 4.979345, 4.976997, 4.97459, 4.97213, 4.969624, 
    4.967066, 4.965834, 4.957517, 4.955821, 4.954513, 4.953405, 4.952485, 
    4.951245, 4.95019, 4.9492, 4.948807, 4.949031, 4.950005, 4.951681, 
    4.954097, 4.956656, 4.959386, 4.961906, 4.964849, 4.968222, 4.972019, 
    4.97623, 4.980836, 4.985796, 4.991051, 4.996513, 5.002068, 5.007562, 
    5.012805, 5.017571, 5.021602, 5.024612, 5.026301, 5.026382, 5.024599, 
    5.020772,
  // totalHeight(26,35, 0-49)
    4.995066, 4.99397, 4.992628, 4.991074, 4.989336, 4.987434, 4.985391, 
    4.983224, 4.98095, 4.978586, 4.976151, 4.97366, 4.971129, 4.968563, 
    4.965956, 4.964484, 4.957617, 4.955689, 4.954103, 4.952727, 4.951577, 
    4.950626, 4.949806, 4.949069, 4.948839, 4.949157, 4.950138, 4.951736, 
    4.953943, 4.956252, 4.958614, 4.961243, 4.964278, 4.967728, 4.971596, 
    4.975876, 4.980554, 4.985588, 4.990923, 4.996468, 5.002102, 5.007667, 
    5.012964, 5.017759, 5.02178, 5.024729, 5.026304, 5.026208, 5.024194, 
    5.02009,
  // totalHeight(26,36, 0-49)
    4.99419, 4.993175, 4.991889, 4.99037, 4.988643, 4.986734, 4.984667, 
    4.98246, 4.980136, 4.977716, 4.975226, 4.972688, 4.970117, 4.967527, 
    4.964915, 4.96312, 4.957703, 4.95561, 4.953803, 4.952217, 4.950887, 
    4.950241, 4.949687, 4.949242, 4.949209, 4.949636, 4.95062, 4.952115, 
    4.954077, 4.95611, 4.958105, 4.960808, 4.963894, 4.967376, 4.971268, 
    4.975566, 4.98026, 4.985313, 4.990666, 4.996232, 5.001882, 5.007453, 
    5.012741, 5.017495, 5.021441, 5.024268, 5.025669, 5.02535, 5.023067, 
    5.018667,
  // totalHeight(26,37, 0-49)
    4.992908, 4.991998, 4.9908, 4.989348, 4.987668, 4.985786, 4.983728, 
    4.981519, 4.979182, 4.976744, 4.974233, 4.971678, 4.969099, 4.966518, 
    4.963937, 4.961798, 4.957793, 4.955594, 4.953619, 4.951871, 4.950411, 
    4.950073, 4.949806, 4.949687, 4.949876, 4.950426, 4.951407, 4.952781, 
    4.954471, 4.956215, 4.957856, 4.9606, 4.963703, 4.967181, 4.971049, 
    4.975317, 4.979972, 4.984982, 4.990291, 4.995806, 5.001399, 5.006898, 
    5.012094, 5.01673, 5.020518, 5.023149, 5.024311, 5.023713, 5.021127, 
    5.016415,
  // totalHeight(26,38, 0-49)
    4.991222, 4.990443, 4.98936, 4.988006, 4.986406, 4.984589, 4.98258, 
    4.980407, 4.978095, 4.975675, 4.97318, 4.970641, 4.968087, 4.965544, 
    4.963021, 4.960566, 4.957904, 4.955646, 4.953547, 4.951684, 4.950138, 
    4.950104, 4.950134, 4.950362, 4.950793, 4.951478, 4.952455, 4.953692, 
    4.955092, 4.956546, 4.957858, 4.960621, 4.96371, 4.967146, 4.970952, 
    4.975142, 4.979702, 4.98461, 4.989802, 4.995189, 5.000639, 5.005978, 
    5.010987, 5.015409, 5.01895, 5.021299, 5.022146, 5.021213, 5.018287, 
    5.013258,
  // totalHeight(26,39, 0-49)
    4.989146, 4.988517, 4.987576, 4.98635, 4.984865, 4.983149, 4.981227, 
    4.979128, 4.976882, 4.974522, 4.972079, 4.969591, 4.967091, 4.96461, 
    4.962165, 4.959454, 4.95805, 4.955768, 4.953585, 4.951646, 4.950048, 
    4.950306, 4.950636, 4.951224, 4.951909, 4.952735, 4.953708, 4.954801, 
    4.955904, 4.957078, 4.958095, 4.960857, 4.963908, 4.967274, 4.970981, 
    4.975045, 4.979459, 4.984196, 4.9892, 4.994374, 4.999588, 5.004664, 
    5.009383, 5.013483, 5.016672, 5.018644, 5.019099, 5.017773, 5.014479, 
    5.009132,
  // totalHeight(26,40, 0-49)
    4.986707, 4.986245, 4.985466, 4.984396, 4.983058, 4.981478, 4.979682, 
    4.977698, 4.975558, 4.973294, 4.970941, 4.968537, 4.966121, 4.963724, 
    4.961371, 4.958483, 4.95824, 4.95596, 4.953722, 4.951737, 4.950122, 
    4.950653, 4.951275, 4.952221, 4.953166, 4.954142, 4.955109, 4.956059, 
    4.956869, 4.957781, 4.958541, 4.961287, 4.964283, 4.967553, 4.97113, 
    4.975026, 4.979239, 4.983742, 4.988476, 4.993349, 4.998224, 5.002929, 
    5.007241, 5.010903, 5.013631, 5.015126, 5.015107, 5.013333, 5.009647, 
    5.004004,
  // totalHeight(26,41, 0-49)
    4.983946, 4.983662, 4.983064, 4.982172, 4.981009, 4.979598, 4.977962, 
    4.976132, 4.974137, 4.972007, 4.969779, 4.967493, 4.965187, 4.962894, 
    4.960647, 4.957664, 4.958471, 4.956212, 4.953946, 4.951943, 4.950333, 
    4.951114, 4.952014, 4.953312, 4.954513, 4.955637, 4.9566, 4.957409, 
    4.957942, 4.95862, 4.959163, 4.961884, 4.964809, 4.967964, 4.97138, 
    4.97507, 4.97903, 4.983232, 4.987618, 4.992094, 4.996525, 5.000741, 
    5.004525, 5.007628, 5.009777, 5.010693, 5.010121, 5.007853, 5.003766, 
    4.997855,
  // totalHeight(26,42, 0-49)
    4.980917, 4.980814, 4.98041, 4.979715, 4.978751, 4.977537, 4.976097, 
    4.974453, 4.972636, 4.970678, 4.968611, 4.966472, 4.964302, 4.962132, 
    4.959999, 4.957001, 4.958748, 4.95652, 4.954246, 4.952245, 4.950657, 
    4.95166, 4.952818, 4.954448, 4.955894, 4.957162, 4.958123, 4.958803, 
    4.95908, 4.959553, 4.959918, 4.962606, 4.965451, 4.968475, 4.971704, 
    4.97515, 4.978807, 4.982642, 4.986598, 4.990582, 4.994461, 4.998068, 
    5.0012, 5.003619, 5.005074, 5.005314, 5.004117, 5.001315, 4.996832, 
    4.990704,
  // totalHeight(26,43, 0-49)
    4.977679, 4.97776, 4.977554, 4.977072, 4.976327, 4.975336, 4.974116, 
    4.972692, 4.971086, 4.969328, 4.967451, 4.965489, 4.963478, 4.961449, 
    4.959437, 4.956493, 4.959065, 4.956875, 4.954607, 4.952624, 4.951071, 
    4.952264, 4.953651, 4.955585, 4.95726, 4.958661, 4.959623, 4.960185, 
    4.960233, 4.960534, 4.960759, 4.963408, 4.966163, 4.96904, 4.97206, 
    4.975228, 4.978531, 4.981936, 4.985381, 4.988777, 4.991995, 4.994875, 
    4.99723, 4.998845, 4.999496, 4.998971, 4.997089, 4.993732, 4.988872, 
    4.982594,
  // totalHeight(26,44, 0-49)
    4.974301, 4.974561, 4.974557, 4.974297, 4.973784, 4.973035, 4.972059, 
    4.970877, 4.96951, 4.967981, 4.966322, 4.964559, 4.962726, 4.960854, 
    4.958971, 4.956134, 4.959414, 4.957269, 4.955017, 4.953065, 4.951551, 
    4.952901, 4.954484, 4.956686, 4.958561, 4.960083, 4.961043, 4.961501, 
    4.961351, 4.961507, 4.961627, 4.964231, 4.966889, 4.969604, 4.972392, 
    4.975247, 4.97815, 4.981063, 4.983919, 4.986634, 4.989085, 4.991127, 
    4.992589, 4.993289, 4.99304, 4.991673, 4.989062, 4.985146, 4.979949, 
    4.973607,
  // totalHeight(26,45, 0-49)
    4.970855, 4.971286, 4.971483, 4.971446, 4.971176, 4.970679, 4.969965, 
    4.969045, 4.967938, 4.96666, 4.965239, 4.963696, 4.962062, 4.960358, 
    4.958611, 4.955917, 4.95979, 4.957693, 4.955468, 4.95355, 4.952076, 
    4.95355, 4.955291, 4.957713, 4.959756, 4.961379, 4.962333, 4.9627, 
    4.962382, 4.962423, 4.96246, 4.965011, 4.967559, 4.970098, 4.972632, 
    4.97514, 4.977598, 4.979958, 4.982154, 4.984101, 4.985687, 4.986785, 
    4.987253, 4.986942, 4.985713, 4.983451, 4.980091, 4.975633, 4.970161, 
    4.963855,
  // totalHeight(26,46, 0-49)
    4.967414, 4.968003, 4.968394, 4.968578, 4.968554, 4.968318, 4.967876, 
    4.967232, 4.9664, 4.96539, 4.964222, 4.962915, 4.961491, 4.959968, 
    4.958365, 4.955836, 4.960183, 4.95814, 4.955951, 4.954069, 4.952631, 
    4.954192, 4.956049, 4.95864, 4.960809, 4.962502, 4.963447, 4.963733, 
    4.963276, 4.963221, 4.963187, 4.965672, 4.968098, 4.970442, 4.972695, 
    4.974825, 4.976792, 4.978544, 4.980013, 4.981115, 4.981754, 4.981822, 
    4.98121, 4.979815, 4.977552, 4.974366, 4.970264, 4.965308, 4.959643, 
    4.953489,
  // totalHeight(26,47, 0-49)
    4.964046, 4.964777, 4.965352, 4.965752, 4.96597, 4.965997, 4.965829, 
    4.96547, 4.96492, 4.964187, 4.963284, 4.962223, 4.961019, 4.959685, 
    4.958235, 4.955878, 4.960584, 4.958601, 4.956454, 4.954607, 4.953197, 
    4.954808, 4.956738, 4.959435, 4.961684, 4.963416, 4.964339, 4.964552, 
    4.96398, 4.963842, 4.963738, 4.966136, 4.968418, 4.970546, 4.972489, 
    4.974205, 4.975642, 4.976735, 4.977419, 4.977613, 4.977237, 4.976211, 
    4.974462, 4.97194, 4.968619, 4.964515, 4.959707, 4.954324, 4.948567, 
    4.942689,
  // totalHeight(26,48, 0-49)
    4.96081, 4.961668, 4.962411, 4.963017, 4.963469, 4.963753, 4.96386, 
    4.963782, 4.963516, 4.963064, 4.962431, 4.961621, 4.960644, 4.959507, 
    4.958216, 4.956029, 4.960979, 4.959066, 4.956965, 4.955151, 4.953761, 
    4.955386, 4.957339, 4.960083, 4.962356, 4.964089, 4.964973, 4.965117, 
    4.964446, 4.964223, 4.964039, 4.966322, 4.968429, 4.970309, 4.971912, 
    4.973177, 4.974042, 4.974437, 4.974288, 4.973528, 4.972093, 4.969935, 
    4.967025, 4.963368, 4.959004, 4.954024, 4.948578, 4.942863, 4.937129, 
    4.93166,
  // totalHeight(26,49, 0-49)
    4.957191, 4.958059, 4.958873, 4.959602, 4.960219, 4.9607, 4.961027, 
    4.961179, 4.961144, 4.960912, 4.960473, 4.959821, 4.95895, 4.957851, 
    4.956515, 4.953525, 4.964903, 4.962058, 4.958658, 4.955644, 4.953284, 
    4.956749, 4.960586, 4.965696, 4.969499, 4.971891, 4.972278, 4.970906, 
    4.967642, 4.965106, 4.962541, 4.964893, 4.966942, 4.968615, 4.969858, 
    4.970594, 4.970757, 4.97027, 4.969067, 4.967099, 4.964337, 4.960783, 
    4.956475, 4.951499, 4.945994, 4.940145, 4.934196, 4.928425, 4.923135, 
    4.918625,
  // totalHeight(27,0, 0-49)
    4.952485, 4.956017, 4.95919, 4.962013, 4.964487, 4.966623, 4.968421, 
    4.969888, 4.971034, 4.971874, 4.972427, 4.972726, 4.972806, 4.972714, 
    4.972504, 4.972033, 4.971988, 4.9717, 4.971503, 4.971475, 4.971662, 
    4.97227, 4.973104, 4.974205, 4.975557, 4.977133, 4.978898, 4.980816, 
    4.982846, 4.984953, 4.987058, 4.989343, 4.991569, 4.993695, 4.995677, 
    4.997463, 4.998989, 5.00017, 5.000906, 5.001068, 5.000506, 4.999043, 
    4.996487, 4.992639, 4.987311, 4.98035, 4.971671, 4.961278, 4.9493, 
    4.936006,
  // totalHeight(27,1, 0-49)
    4.953785, 4.957267, 4.960383, 4.963142, 4.965549, 4.967614, 4.969344, 
    4.970743, 4.971827, 4.97261, 4.973116, 4.973373, 4.973421, 4.973308, 
    4.973083, 4.972408, 4.972571, 4.972211, 4.971914, 4.971784, 4.971873, 
    4.97256, 4.97343, 4.974563, 4.975933, 4.977504, 4.979235, 4.981091, 
    4.983034, 4.985042, 4.987011, 4.989357, 4.991658, 4.993884, 4.995999, 
    4.997962, 4.999713, 5.001177, 5.002253, 5.002817, 5.002716, 5.001765, 
    4.999763, 4.996496, 4.991755, 4.985361, 4.977194, 4.967225, 4.955546, 
    4.942395,
  // totalHeight(27,2, 0-49)
    4.9551, 4.958522, 4.961576, 4.964267, 4.96661, 4.96861, 4.970279, 
    4.971625, 4.97266, 4.973405, 4.97388, 4.974118, 4.974155, 4.974039, 
    4.97382, 4.972966, 4.973311, 4.972891, 4.972506, 4.972278, 4.972264, 
    4.973009, 4.97389, 4.975019, 4.976368, 4.9779, 4.979566, 4.981339, 
    4.983176, 4.985064, 4.98687, 4.989237, 4.991573, 4.993855, 4.996058, 
    4.998144, 5.000066, 5.00175, 5.003102, 5.003998, 5.004288, 5.003786, 
    5.002285, 4.999563, 4.995397, 4.989588, 4.981988, 4.972539, 4.961292, 
    4.948447,
  // totalHeight(27,3, 0-49)
    4.956424, 4.959782, 4.962767, 4.965392, 4.967669, 4.969612, 4.971227, 
    4.972527, 4.973528, 4.974247, 4.97471, 4.974946, 4.974991, 4.974892, 
    4.974695, 4.973688, 4.974173, 4.973708, 4.973245, 4.972928, 4.972816, 
    4.973597, 4.974463, 4.975552, 4.976844, 4.978302, 4.979884, 4.981561, 
    4.983288, 4.985043, 4.986671, 4.989024, 4.991359, 4.993658, 4.995905, 
    4.99807, 5.000108, 5.001954, 5.003517, 5.004678, 5.00529, 5.005171, 
    5.004114, 5.001892, 4.998278, 4.993056, 4.986063, 4.977203, 4.966496, 
    4.9541,
  // totalHeight(27,4, 0-49)
    4.957763, 4.961049, 4.963962, 4.966518, 4.968731, 4.970614, 4.97218, 
    4.973444, 4.974419, 4.975125, 4.975588, 4.975837, 4.975906, 4.975838, 
    4.975676, 4.974549, 4.975114, 4.974617, 4.974098, 4.973704, 4.973499, 
    4.974296, 4.97512, 4.976135, 4.977338, 4.978698, 4.980179, 4.981754, 
    4.983374, 4.984993, 4.986437, 4.988748, 4.991049, 4.993332, 4.995584, 
    4.997785, 4.999891, 5.001845, 5.003561, 5.004924, 5.005792, 5.005991, 
    5.00532, 5.003553, 5.000459, 4.995819, 4.98945, 4.981233, 4.971154, 
    4.959323,
  // totalHeight(27,5, 0-49)
    4.959124, 4.96233, 4.965165, 4.967649, 4.969796, 4.971621, 4.973139, 
    4.974367, 4.975321, 4.976024, 4.976496, 4.976768, 4.976871, 4.976844, 
    4.976726, 4.975518, 4.976087, 4.975574, 4.975018, 4.974565, 4.97428, 
    4.975071, 4.975831, 4.976738, 4.977826, 4.979064, 4.980437, 4.981911, 
    4.983433, 4.984925, 4.986189, 4.988428, 4.990667, 4.992902, 4.995128, 
    4.997325, 4.999457, 5.001471, 5.003284, 5.004794, 5.005862, 5.006324, 
    5.005984, 5.004626, 5.002022, 4.997947, 4.992211, 4.984674, 4.975287, 
    4.964118,
  // totalHeight(27,6, 0-49)
    4.960515, 4.963633, 4.966385, 4.96879, 4.970866, 4.972629, 4.974098, 
    4.975291, 4.976225, 4.976924, 4.97741, 4.977711, 4.977855, 4.977876, 
    4.977808, 4.976558, 4.977046, 4.976531, 4.97596, 4.975471, 4.975124, 
    4.975888, 4.976562, 4.977334, 4.978279, 4.979381, 4.980637, 4.982016, 
    4.983459, 4.984834, 4.985934, 4.988077, 4.990227, 4.992387, 4.994555, 
    4.996716, 4.998837, 5.000868, 5.002738, 5.004347, 5.005566, 5.006243, 
    5.006188, 5.005199, 5.003053, 4.999527, 4.994426, 4.987591, 4.978942, 
    4.968504,
  // totalHeight(27,7, 0-49)
    4.961944, 4.964969, 4.96763, 4.969948, 4.971945, 4.97364, 4.975054, 
    4.976207, 4.977119, 4.977812, 4.978312, 4.978641, 4.978827, 4.978899, 
    4.97888, 4.977633, 4.977947, 4.977446, 4.976884, 4.976382, 4.975995, 
    4.976711, 4.97728, 4.977891, 4.978675, 4.97963, 4.980768, 4.982057, 
    4.98344, 4.984717, 4.985673, 4.987694, 4.989734, 4.991795, 4.99388, 
    4.995977, 4.998057, 5.000075, 5.001965, 5.003634, 5.004968, 5.005818, 
    5.006014, 5.00536, 5.003646, 5.000652, 4.996178, 4.990054, 4.982172, 
    4.972516,
  // totalHeight(27,8, 0-49)
    4.96342, 4.966343, 4.968904, 4.971127, 4.973035, 4.974654, 4.976002, 
    4.977108, 4.977989, 4.978671, 4.979177, 4.979532, 4.979758, 4.979877, 
    4.979905, 4.978708, 4.978746, 4.978274, 4.97775, 4.977262, 4.976861, 
    4.977507, 4.977953, 4.978384, 4.978992, 4.979788, 4.980811, 4.982022, 
    4.983364, 4.984567, 4.985405, 4.987285, 4.989192, 4.991133, 4.993113, 
    4.995123, 4.997139, 4.999117, 5.001001, 5.002707, 5.004125, 5.005124, 
    5.005543, 5.005198, 5.003892, 5.001414, 4.997559, 4.992144, 4.985043, 
    4.976196,
  // totalHeight(27,9, 0-49)
    4.964952, 4.967762, 4.970212, 4.972329, 4.974138, 4.975667, 4.976941, 
    4.977984, 4.978825, 4.979486, 4.97999, 4.980362, 4.98062, 4.980781, 
    4.980847, 4.979746, 4.979405, 4.97898, 4.978518, 4.978075, 4.977688, 
    4.978245, 4.978553, 4.978786, 4.97921, 4.979844, 4.980752, 4.981893, 
    4.983215, 4.984366, 4.985122, 4.98684, 4.988597, 4.990402, 4.992261, 
    4.994167, 4.9961, 4.998025, 4.999886, 5.001608, 5.003094, 5.004222, 
    5.004846, 5.004794, 5.003879, 5.001898, 4.998647, 4.993936, 4.987614, 
    4.979589,
  // totalHeight(27,10, 0-49)
    4.966544, 4.969228, 4.971554, 4.973551, 4.975248, 4.976675, 4.977859, 
    4.97883, 4.979616, 4.980243, 4.980734, 4.981112, 4.98139, 4.981582, 
    4.981678, 4.980717, 4.979891, 4.979529, 4.979159, 4.978791, 4.978449, 
    4.978896, 4.979054, 4.97908, 4.979313, 4.979784, 4.980581, 4.981661, 
    4.982981, 4.984105, 4.984818, 4.986358, 4.987952, 4.989606, 4.991331, 
    4.993123, 4.994964, 4.996823, 4.998651, 5.000382, 5.001927, 5.003174, 
    5.003991, 5.00422, 5.003681, 5.002182, 4.999519, 4.995496, 4.989943, 
    4.982737,
  // totalHeight(27,11, 0-49)
    4.968184, 4.970732, 4.972922, 4.974787, 4.976358, 4.97767, 4.978752, 
    4.979636, 4.980354, 4.980931, 4.981393, 4.981763, 4.982052, 4.982261, 
    4.982378, 4.981594, 4.980174, 4.979899, 4.979648, 4.979387, 4.979123, 
    4.979436, 4.979437, 4.979248, 4.979291, 4.979603, 4.980292, 4.981318, 
    4.98265, 4.983774, 4.984485, 4.985836, 4.987253, 4.988749, 4.990333, 
    4.992004, 4.993749, 4.995539, 4.997333, 4.99907, 5.000671, 5.002034, 
    5.00304, 5.00354, 5.003365, 5.00233, 5.000237, 4.996881, 4.992076, 
    4.985673,
  // totalHeight(27,12, 0-49)
    4.969869, 4.972264, 4.974305, 4.976025, 4.977458, 4.978641, 4.979606, 
    4.98039, 4.981024, 4.981538, 4.981959, 4.982306, 4.982589, 4.982803, 
    4.982933, 4.982355, 4.980234, 4.98007, 4.979968, 4.979845, 4.979689, 
    4.97985, 4.979685, 4.979283, 4.979139, 4.979298, 4.979885, 4.980863, 
    4.982218, 4.983363, 4.984119, 4.985269, 4.986504, 4.987836, 4.989278, 
    4.990828, 4.992476, 4.9942, 4.995962, 4.997709, 4.999368, 5.000849, 
    5.002039, 5.002804, 5.002984, 5.002398, 5.00085, 4.998134, 4.99405, 
    4.988423,
  // totalHeight(27,13, 0-49)
    4.971578, 4.973805, 4.975684, 4.977247, 4.978529, 4.979571, 4.980408, 
    4.98108, 4.981618, 4.982056, 4.982419, 4.982728, 4.982991, 4.983199, 
    4.983337, 4.982982, 4.980053, 4.980028, 4.980104, 4.980148, 4.980134, 
    4.980123, 4.97979, 4.979178, 4.978858, 4.978872, 4.979362, 4.980295, 
    4.981681, 4.982868, 4.983716, 4.984661, 4.98571, 4.986878, 4.988178, 
    4.989611, 4.991169, 4.992833, 4.994571, 4.996334, 4.998056, 4.999658, 
    5.001034, 5.002057, 5.002578, 5.002422, 5.001395, 4.999288, 4.995888, 
    4.991003,
  // totalHeight(27,14, 0-49)
    4.973285, 4.975332, 4.977035, 4.978428, 4.979551, 4.980443, 4.981143, 
    4.981692, 4.982125, 4.982474, 4.982768, 4.983025, 4.983253, 4.983449, 
    4.983591, 4.983465, 4.979623, 4.979764, 4.980047, 4.980291, 4.980448, 
    4.980245, 4.979743, 4.978934, 4.978452, 4.978334, 4.978735, 4.979624, 
    4.981044, 4.98229, 4.983274, 4.984014, 4.98488, 4.985888, 4.987052, 
    4.988374, 4.98985, 4.991462, 4.993183, 4.994971, 4.996765, 4.998491, 
    5.000052, 5.001328, 5.002178, 5.002431, 5.001897, 5.000363, 4.99761, 
    4.993423,
  // totalHeight(27,15, 0-49)
    4.974969, 4.976818, 4.97833, 4.979544, 4.980499, 4.981234, 4.981791, 
    4.982209, 4.982529, 4.98278, 4.982994, 4.983189, 4.983375, 4.983549, 
    4.983696, 4.983794, 4.978942, 4.979278, 4.979795, 4.980265, 4.98062, 
    4.980211, 4.979545, 4.978554, 4.977929, 4.977694, 4.978014, 4.978863, 
    4.980318, 4.981638, 4.982798, 4.983336, 4.984023, 4.984879, 4.985915, 
    4.987135, 4.988539, 4.990111, 4.991827, 4.993648, 4.99552, 4.997373, 
    4.999117, 5.000638, 5.001802, 5.002442, 5.002368, 5.00137, 4.999219, 
    4.995688,
  // totalHeight(27,16, 0-49)
    4.9766, 4.978232, 4.979541, 4.980565, 4.981343, 4.981917, 4.982327, 
    4.982615, 4.982817, 4.982967, 4.983095, 4.98322, 4.983356, 4.983504, 
    4.983661, 4.983968, 4.978021, 4.978576, 4.979346, 4.980065, 4.980643, 
    4.980015, 4.979194, 4.97804, 4.977294, 4.976964, 4.977215, 4.978029, 
    4.979517, 4.980919, 4.982292, 4.982636, 4.983153, 4.983865, 4.984783, 
    4.985914, 4.987255, 4.988797, 4.990517, 4.992379, 4.994334, 4.996316, 
    4.99824, 4.999999, 5.001459, 5.002461, 5.002818, 5.002316, 5.000722, 
    4.997799,
  // totalHeight(27,17, 0-49)
    4.97815, 4.979545, 4.980634, 4.981458, 4.982053, 4.982463, 4.982728, 
    4.982884, 4.982973, 4.983024, 4.983063, 4.983118, 4.983199, 4.983321, 
    4.983489, 4.983988, 4.976887, 4.977677, 4.978717, 4.979698, 4.980515, 
    4.97966, 4.978692, 4.977397, 4.976559, 4.976156, 4.976355, 4.977139, 
    4.97866, 4.980151, 4.981763, 4.981924, 4.982281, 4.982859, 4.983669, 
    4.98472, 4.986009, 4.987531, 4.989263, 4.991172, 4.993215, 4.995326, 
    4.997425, 4.999409, 5.001151, 5.00249, 5.003245, 5.0032, 5.002119, 
    4.999754,
  // totalHeight(27,18, 0-49)
    4.979592, 4.980724, 4.981576, 4.982186, 4.982595, 4.982841, 4.982964, 
    4.983, 4.982983, 4.982941, 4.9829, 4.982886, 4.982915, 4.983007, 
    4.983186, 4.983865, 4.975588, 4.976619, 4.977927, 4.979177, 4.980241, 
    4.979152, 4.978045, 4.976635, 4.97573, 4.975284, 4.975449, 4.976212, 
    4.977769, 4.979352, 4.981221, 4.981211, 4.981418, 4.981871, 4.982583, 
    4.983562, 4.984807, 4.986314, 4.988064, 4.990025, 4.992156, 4.994394, 
    4.996664, 4.998864, 5.000867, 5.002522, 5.003644, 5.004018, 5.003407, 
    5.001557,
  // totalHeight(27,19, 0-49)
    4.980903, 4.98174, 4.98233, 4.982714, 4.982932, 4.983019, 4.98301, 
    4.982938, 4.982831, 4.982711, 4.982603, 4.982526, 4.982506, 4.982572, 
    4.982763, 4.983617, 4.9742, 4.975467, 4.977031, 4.978539, 4.979841, 
    4.978513, 4.97728, 4.975773, 4.974828, 4.974364, 4.974518, 4.975278, 
    4.976873, 4.978549, 4.980679, 4.98051, 4.980577, 4.980914, 4.981531, 
    4.982439, 4.983643, 4.985138, 4.986907, 4.988921, 4.991139, 4.993503, 
    4.995936, 4.998341, 5.000593, 5.002542, 5.004004, 5.004765, 5.004586, 
    5.00321,
  // totalHeight(27,20, 0-49)
    4.982862, 4.984146, 4.985185, 4.986007, 4.98664, 4.987111, 4.987448, 
    4.987677, 4.987826, 4.987921, 4.987986, 4.988048, 4.988135, 4.988278, 
    4.988526, 30, 4.972143, 4.973258, 4.97473, 4.976183, 4.977445, 4.975578, 
    4.973876, 4.971932, 4.970649, 4.969963, 4.970038, 4.970872, 4.97272, 
    4.974809, 4.977582, 4.977671, 4.978006, 4.978611, 4.979485, 4.980634, 
    4.982059, 4.983755, 4.985709, 4.987898, 4.990287, 4.992825, 4.995441, 
    4.998047, 5.000524, 5.002726, 5.004475, 5.005559, 5.005739, 5.004762,
  // totalHeight(27,21, 0-49)
    4.984021, 4.985055, 4.985878, 4.986519, 4.987, 4.98735, 4.987592, 
    4.987746, 4.987836, 4.987881, 4.987903, 4.987926, 4.987977, 4.98809, 
    4.988317, 30, 4.96787, 4.969113, 4.970778, 4.972454, 4.973938, 4.971829, 
    4.970017, 4.96804, 4.966849, 4.966359, 4.966709, 4.967876, 4.970111, 
    4.97262, 4.975931, 4.976147, 4.976643, 4.977433, 4.978511, 4.979876, 
    4.981517, 4.983426, 4.985584, 4.987966, 4.990533, 4.993235, 4.996002, 
    4.998747, 5.001359, 5.003693, 5.005579, 5.006813, 5.007162, 5.006378,
  // totalHeight(27,22, 0-49)
    4.9851, 4.985905, 4.986529, 4.987001, 4.987345, 4.987583, 4.987735, 
    4.987818, 4.987849, 4.987846, 4.987824, 4.987807, 4.987818, 4.987895, 
    4.988095, 30, 4.96427, 4.965615, 4.967438, 4.969296, 4.970961, 4.968601, 
    4.96665, 4.964593, 4.963428, 4.963049, 4.963583, 4.964988, 4.96751, 
    4.970334, 4.974064, 4.974349, 4.974948, 4.975873, 4.977114, 4.978661, 
    4.980502, 4.982621, 4.984995, 4.987593, 4.990371, 4.993275, 4.996236, 
    4.999167, 5.001956, 5.004463, 5.006518, 5.007926, 5.008459, 5.007876,
  // totalHeight(27,23, 0-49)
    4.986108, 4.986693, 4.987132, 4.98745, 4.987665, 4.987799, 4.987868, 
    4.987884, 4.987857, 4.987806, 4.987741, 4.98768, 4.987649, 4.987686, 
    4.987846, 30, 4.961174, 4.962575, 4.964491, 4.966458, 4.968225, 4.965626, 
    4.963521, 4.961361, 4.960176, 4.959849, 4.960501, 4.962069, 4.964801, 
    4.96786, 4.971903, 4.972238, 4.972919, 4.973962, 4.97535, 4.977074, 
    4.979115, 4.981455, 4.984063, 4.986903, 4.989927, 4.993075, 4.996275, 
    4.999434, 5.00244, 5.005151, 5.007399, 5.008994, 5.009711, 5.00932,
  // totalHeight(27,24, 0-49)
    4.987052, 4.987432, 4.987696, 4.987866, 4.987962, 4.987997, 4.987984, 
    4.987933, 4.987851, 4.98775, 4.987639, 4.987533, 4.987454, 4.987441, 
    4.987548, 30, 4.958886, 4.960289, 4.962229, 4.964231, 4.966028, 4.963264, 
    4.961052, 4.958817, 4.957613, 4.957313, 4.958032, 4.959703, 4.962571, 
    4.965787, 4.970043, 4.970445, 4.971216, 4.972371, 4.973891, 4.975769, 
    4.977979, 4.980506, 4.983313, 4.986362, 4.989601, 4.992966, 4.996381, 
    4.99975, 5.002959, 5.005866, 5.0083, 5.010072, 5.010966, 5.010753,
  // totalHeight(27,25, 0-49)
    4.987951, 4.988135, 4.988231, 4.988259, 4.988237, 4.988174, 4.98808, 
    4.987959, 4.987818, 4.987662, 4.987497, 4.987339, 4.987206, 4.987133, 
    4.987175, 30, 4.957164, 4.958512, 4.960404, 4.962363, 4.964118, 4.961286, 
    4.959035, 4.956786, 4.955588, 4.955317, 4.956082, 4.957819, 4.960765, 
    4.964076, 4.968446, 4.968953, 4.969841, 4.971123, 4.972783, 4.974807, 
    4.977177, 4.979869, 4.98285, 4.986078, 4.989499, 4.993052, 4.996652, 
    5.000207, 5.003596, 5.006678, 5.009283, 5.011218, 5.01227, 5.012215,
  // totalHeight(27,26, 0-49)
    4.988813, 4.988812, 4.98875, 4.988639, 4.9885, 4.988336, 4.988153, 
    4.987953, 4.987741, 4.987518, 4.98729, 4.987069, 4.986872, 4.986731, 
    4.986691, 30, 4.956017, 4.957257, 4.959034, 4.960871, 4.962512, 4.95972, 
    4.957509, 4.955312, 4.954154, 4.953917, 4.954714, 4.956479, 4.959447, 
    4.962788, 4.967175, 4.967828, 4.968863, 4.970294, 4.972103, 4.974275, 
    4.976792, 4.979629, 4.982756, 4.986129, 4.989699, 4.9934, 4.997152, 
    5.000857, 5.004397, 5.007628, 5.010381, 5.01246, 5.013651, 5.013734,
  // totalHeight(27,27, 0-49)
    4.98965, 4.989479, 4.989264, 4.98902, 4.988759, 4.988484, 4.9882, 
    4.987906, 4.987603, 4.987295, 4.986986, 4.986688, 4.986415, 4.986197, 
    4.986067, 30, 4.955529, 4.956617, 4.958216, 4.959864, 4.961324, 4.958663, 
    4.956551, 4.954452, 4.95335, 4.953136, 4.95393, 4.955672, 4.958594, 
    4.961887, 4.966184, 4.967004, 4.968203, 4.969788, 4.971744, 4.974054, 
    4.976701, 4.979663, 4.98291, 4.986403, 4.990092, 4.993917, 4.997795, 
    5.001633, 5.005309, 5.008677, 5.011567, 5.013782, 5.015105, 5.01531,
  // totalHeight(27,28, 0-49)
    4.990469, 4.990145, 4.989788, 4.989411, 4.989022, 4.988625, 4.988218, 
    4.987805, 4.987385, 4.986967, 4.986554, 4.98616, 4.985801, 4.9855, 
    4.985283, 30, 4.956028, 4.956934, 4.958307, 4.959707, 4.96093, 4.958463, 
    4.956476, 4.954484, 4.953412, 4.953169, 4.953884, 4.955516, 4.958292, 
    4.961439, 4.965523, 4.966502, 4.967848, 4.969568, 4.971642, 4.974057, 
    4.976798, 4.979848, 4.983181, 4.986762, 4.990545, 4.994473, 4.998466, 
    5.002428, 5.006239, 5.009749, 5.012783, 5.015139, 5.016596, 5.016923,
  // totalHeight(27,29, 0-49)
    4.991272, 4.99082, 4.990334, 4.989828, 4.989304, 4.988763, 4.988209, 
    4.987643, 4.987072, 4.986504, 4.985958, 4.985448, 4.984994, 4.984619, 
    4.984338, 30, 4.957261, 4.957983, 4.959101, 4.960205, 4.96113, 4.958851, 
    4.956955, 4.955013, 4.953891, 4.953528, 4.954064, 4.955482, 4.958002, 
    4.960886, 4.964627, 4.965713, 4.967158, 4.968967, 4.971126, 4.973623, 
    4.976449, 4.979589, 4.983022, 4.986718, 4.990633, 4.994709, 4.998869, 
    5.003012, 5.00701, 5.010713, 5.013935, 5.016467, 5.018081, 5.018536,
  // totalHeight(27,30, 0-49)
    4.991342, 4.990104, 4.98886, 4.987627, 4.986415, 4.985223, 4.984044, 
    4.982868, 4.981678, 4.980457, 4.979197, 4.977892, 4.976555, 4.975228, 
    4.973989, 4.972118, 4.961142, 4.961493, 4.962195, 4.962931, 4.963588, 
    4.961671, 4.96014, 4.958567, 4.957699, 4.957439, 4.957901, 4.95906, 
    4.961126, 4.963423, 4.966387, 4.96713, 4.968222, 4.969685, 4.971525, 
    4.973748, 4.976355, 4.979339, 4.982685, 4.986363, 4.990328, 4.994513, 
    4.998833, 5.003178, 5.007408, 5.011355, 5.014824, 5.017593, 5.019419, 
    5.020052,
  // totalHeight(27,31, 0-49)
    4.992085, 4.990796, 4.989485, 4.988165, 4.986845, 4.985525, 4.9842, 
    4.982865, 4.981511, 4.980129, 4.978714, 4.977267, 4.975796, 4.974329, 
    4.972923, 4.971511, 4.96095, 4.960932, 4.961246, 4.961601, 4.961905, 
    4.960153, 4.958697, 4.957186, 4.956329, 4.956063, 4.956516, 4.957662, 
    4.959669, 4.961869, 4.964588, 4.965552, 4.966871, 4.968566, 4.970642, 
    4.973103, 4.975951, 4.979178, 4.982767, 4.986686, 4.990888, 4.995302, 
    4.99984, 5.004383, 5.008787, 5.012877, 5.016449, 5.019275, 5.021107, 
    5.021693,
  // totalHeight(27,32, 0-49)
    4.992704, 4.991362, 4.989981, 4.988571, 4.987143, 4.985699, 4.984235, 
    4.982752, 4.981244, 4.979711, 4.978148, 4.976559, 4.974949, 4.97334, 
    4.971759, 4.970668, 4.96088, 4.960486, 4.96041, 4.960387, 4.96035, 
    4.958791, 4.957444, 4.956033, 4.955215, 4.954963, 4.95541, 4.956527, 
    4.958438, 4.960497, 4.962925, 4.964082, 4.965597, 4.967487, 4.969763, 
    4.972429, 4.975488, 4.97893, 4.982742, 4.986887, 4.991313, 4.995951, 
    5.000702, 5.005444, 5.010021, 5.014254, 5.017927, 5.020806, 5.022637, 
    5.023165,
  // totalHeight(27,33, 0-49)
    4.993176, 4.991786, 4.990337, 4.988843, 4.987313, 4.98575, 4.984156, 
    4.982533, 4.980882, 4.979203, 4.977501, 4.975778, 4.97404, 4.972296, 
    4.97056, 4.969613, 4.960853, 4.960111, 4.959667, 4.95929, 4.95894, 
    4.957603, 4.956401, 4.955134, 4.954391, 4.954172, 4.954613, 4.955681, 
    4.957458, 4.959333, 4.961436, 4.962754, 4.964429, 4.966482, 4.968922, 
    4.971757, 4.974994, 4.978625, 4.982632, 4.986979, 4.991614, 4.996459, 
    5.001411, 5.006339, 5.011081, 5.015445, 5.019209, 5.022128, 5.023943, 
    5.024394,
  // totalHeight(27,34, 0-49)
    4.993468, 4.992046, 4.990543, 4.988973, 4.98735, 4.985679, 4.983964, 
    4.982211, 4.980426, 4.978615, 4.976783, 4.974936, 4.973081, 4.971223, 
    4.96936, 4.968389, 4.960826, 4.959777, 4.958998, 4.958305, 4.957679, 
    4.956588, 4.955568, 4.954486, 4.953852, 4.953686, 4.95412, 4.955118, 
    4.956721, 4.958376, 4.960136, 4.961588, 4.963395, 4.965575, 4.968145, 
    4.971118, 4.974501, 4.978288, 4.98246, 4.986983, 4.9918, 4.996827, 
    5.001957, 5.00705, 5.011934, 5.016407, 5.020238, 5.023174, 5.024948, 
    5.025294,
  // totalHeight(27,35, 0-49)
    4.993543, 4.992109, 4.990572, 4.988945, 4.987246, 4.98548, 4.983659, 
    4.98179, 4.979885, 4.977952, 4.976004, 4.97405, 4.972095, 4.970143, 
    4.968186, 4.967057, 4.960784, 4.959477, 4.958406, 4.957438, 4.956577, 
    4.955748, 4.954938, 4.954085, 4.953589, 4.953495, 4.953919, 4.954828, 
    4.956221, 4.957632, 4.959045, 4.960607, 4.962515, 4.964794, 4.967463, 
    4.970541, 4.974034, 4.977944, 4.982249, 4.986913, 4.991876, 4.997052, 
    5.002326, 5.007547, 5.012538, 5.017087, 5.020951, 5.023866, 5.025561, 
    5.025771,
  // totalHeight(27,36, 0-49)
    4.993363, 4.991943, 4.990395, 4.988733, 4.986978, 4.985139, 4.983231, 
    4.981265, 4.979257, 4.977222, 4.975175, 4.973129, 4.971095, 4.969073, 
    4.967054, 4.965679, 4.960728, 4.959213, 4.957893, 4.956695, 4.95564, 
    4.955082, 4.954507, 4.953914, 4.953588, 4.953581, 4.953995, 4.954797, 
    4.955952, 4.957104, 4.958177, 4.959828, 4.961814, 4.964163, 4.966903, 
    4.970053, 4.973625, 4.977619, 4.982017, 4.986782, 4.991848, 4.997127, 
    5.002496, 5.007801, 5.012851, 5.017424, 5.021269, 5.024117, 5.025689, 
    5.025723,
  // totalHeight(27,37, 0-49)
    4.992894, 4.991515, 4.989983, 4.988314, 4.986529, 4.984643, 4.982672, 
    4.980633, 4.978547, 4.97643, 4.974305, 4.972188, 4.970094, 4.968026, 
    4.965975, 4.964311, 4.960664, 4.958989, 4.957465, 4.956078, 4.95487, 
    4.954582, 4.954257, 4.953956, 4.953823, 4.953918, 4.954322, 4.955003, 
    4.955902, 4.956789, 4.957542, 4.959267, 4.961312, 4.963708, 4.96649, 
    4.969682, 4.973296, 4.977336, 4.981783, 4.986598, 4.991717, 4.997042, 
    5.00245, 5.007774, 5.01282, 5.017355, 5.021121, 5.02384, 5.025236, 
    5.025045,
  // totalHeight(27,38, 0-49)
    4.992102, 4.990796, 4.989309, 4.987664, 4.985879, 4.983975, 4.981972, 
    4.979889, 4.977752, 4.97558, 4.973402, 4.971236, 4.969102, 4.967009, 
    4.964951, 4.962999, 4.960605, 4.958811, 4.957121, 4.955583, 4.954257, 
    4.954235, 4.954173, 4.954182, 4.954263, 4.954476, 4.954871, 4.955422, 
    4.956054, 4.956684, 4.957149, 4.958934, 4.961021, 4.963445, 4.966245, 
    4.969447, 4.97307, 4.977113, 4.981561, 4.986373, 4.991481, 4.996788, 
    5.002161, 5.007431, 5.012395, 5.016815, 5.020426, 5.022949, 5.024106, 
    5.023642,
  // totalHeight(27,39, 0-49)
    4.990971, 4.989764, 4.988355, 4.986764, 4.985014, 4.983126, 4.981123, 
    4.97903, 4.976871, 4.974676, 4.97247, 4.970282, 4.968132, 4.966033, 
    4.963985, 4.961775, 4.960558, 4.95868, 4.956858, 4.955204, 4.953793, 
    4.954025, 4.954226, 4.954561, 4.954874, 4.955217, 4.955606, 4.956029, 
    4.956393, 4.956779, 4.956996, 4.958832, 4.960948, 4.963384, 4.966179, 
    4.969365, 4.972958, 4.976961, 4.981358, 4.986107, 4.991138, 4.99635, 
    5.001607, 5.006737, 5.011529, 5.015744, 5.019113, 5.021358, 5.022209, 
    5.021421,
  // totalHeight(27,40, 0-49)
    4.989492, 4.988411, 4.987108, 4.985605, 4.983923, 4.982087, 4.980121, 
    4.978053, 4.975909, 4.973721, 4.971519, 4.969333, 4.96719, 4.965103, 
    4.963079, 4.960662, 4.960529, 4.958594, 4.956668, 4.954926, 4.953461, 
    4.953931, 4.954395, 4.955062, 4.955615, 4.956097, 4.956487, 4.956788, 
    4.956896, 4.957064, 4.957074, 4.958955, 4.961094, 4.963527, 4.966299, 
    4.96944, 4.972969, 4.976889, 4.98118, 4.9858, 4.990678, 4.995711, 
    5.000761, 5.005651, 5.010171, 5.01408, 5.017112, 5.018996, 5.019468, 
    5.018303,
  // totalHeight(27,41, 0-49)
    4.98767, 4.986738, 4.98557, 4.984185, 4.982606, 4.98086, 4.978968, 
    4.97696, 4.974867, 4.972721, 4.970555, 4.9684, 4.966283, 4.964226, 
    4.962235, 4.959669, 4.96052, 4.958544, 4.956538, 4.954738, 4.95324, 
    4.953933, 4.95465, 4.955646, 4.956444, 4.957076, 4.957476, 4.957663, 
    4.957536, 4.957518, 4.957366, 4.959292, 4.961448, 4.963868, 4.9666, 
    4.969671, 4.973102, 4.976892, 4.98102, 4.985444, 4.99009, 4.994852, 
    4.999594, 5.004138, 5.008276, 5.01177, 5.014363, 5.015793, 5.015814, 
    5.014226,
  // totalHeight(27,42, 0-49)
    4.985522, 4.98476, 4.983753, 4.982516, 4.981074, 4.97945, 4.977669, 
    4.975759, 4.973754, 4.971684, 4.969582, 4.967484, 4.965418, 4.963405, 
    4.961457, 4.958804, 4.960528, 4.958524, 4.956461, 4.954623, 4.953115, 
    4.954007, 4.954963, 4.956277, 4.957321, 4.958108, 4.958529, 4.958621, 
    4.958286, 4.958118, 4.957849, 4.959821, 4.961989, 4.96439, 4.967066, 
    4.970046, 4.973344, 4.976959, 4.980868, 4.985023, 4.989351, 4.993749, 
    4.998077, 5.002162, 5.005802, 5.008768, 5.010814, 5.011698, 5.011199, 
    5.009146,
  // totalHeight(27,43, 0-49)
    4.983078, 4.982504, 4.981679, 4.980618, 4.979343, 4.977874, 4.976239, 
    4.974464, 4.972579, 4.970617, 4.968614, 4.966598, 4.964602, 4.962647, 
    4.96075, 4.958064, 4.960546, 4.958526, 4.956423, 4.954565, 4.953062, 
    4.954131, 4.955307, 4.956923, 4.958204, 4.959147, 4.959601, 4.959621, 
    4.959113, 4.958833, 4.958492, 4.960511, 4.962692, 4.965067, 4.967675, 
    4.97054, 4.973672, 4.977067, 4.980697, 4.984512, 4.988438, 4.992373, 
    4.996177, 4.999687, 5.00271, 5.00503, 5.006423, 5.006673, 5.005592, 
    5.003043,
  // totalHeight(27,44, 0-49)
    4.980382, 4.980007, 4.979383, 4.978521, 4.97744, 4.976157, 4.974699, 
    4.973089, 4.971357, 4.969535, 4.967654, 4.965747, 4.963842, 4.961959, 
    4.960116, 4.957444, 4.96057, 4.958542, 4.956412, 4.954548, 4.953062, 
    4.954283, 4.955656, 4.957548, 4.959053, 4.960151, 4.960651, 4.960621, 
    4.959981, 4.95963, 4.959256, 4.961325, 4.963518, 4.965861, 4.968388, 
    4.971116, 4.974051, 4.97718, 4.980473, 4.983876, 4.987314, 4.990685, 
    4.993859, 4.996679, 4.998967, 5.000529, 5.001168, 5.000703, 4.998985, 
    4.995923,
  // totalHeight(27,45, 0-49)
    4.977487, 4.977318, 4.976908, 4.976263, 4.975397, 4.974328, 4.973073, 
    4.971658, 4.970108, 4.968452, 4.96672, 4.964941, 4.963143, 4.961346, 
    4.959565, 4.956938, 4.960594, 4.958564, 4.956421, 4.954561, 4.953098, 
    4.954445, 4.955987, 4.958123, 4.959834, 4.961078, 4.961632, 4.961581, 
    4.960852, 4.960466, 4.960093, 4.962214, 4.964419, 4.966725, 4.969159, 
    4.971728, 4.974432, 4.977252, 4.980149, 4.983069, 4.985935, 4.988648, 
    4.991086, 4.993104, 4.994545, 4.995243, 4.995037, 4.993789, 4.991396, 
    4.987819,
  // totalHeight(27,46, 0-49)
    4.974452, 4.974493, 4.974304, 4.97389, 4.973258, 4.972421, 4.971393, 
    4.970196, 4.968852, 4.967385, 4.965823, 4.964191, 4.962515, 4.960814, 
    4.959103, 4.956544, 4.960613, 4.958589, 4.956441, 4.954591, 4.953156, 
    4.954598, 4.956281, 4.95862, 4.960506, 4.961886, 4.962506, 4.96246, 
    4.961684, 4.961299, 4.960954, 4.963126, 4.965339, 4.9676, 4.969926, 
    4.972314, 4.974755, 4.97722, 4.979667, 4.982036, 4.98425, 4.986214, 
    4.987817, 4.988932, 4.989427, 4.989168, 4.988042, 4.98596, 4.982873, 
    4.9788,
  // totalHeight(27,47, 0-49)
    4.971342, 4.971589, 4.971627, 4.971451, 4.971065, 4.970476, 4.969693, 
    4.968733, 4.967612, 4.966353, 4.964977, 4.963507, 4.961967, 4.960371, 
    4.958735, 4.956259, 4.960622, 4.95861, 4.956469, 4.954632, 4.953219, 
    4.954731, 4.956517, 4.959014, 4.961045, 4.962544, 4.963233, 4.963216, 
    4.962434, 4.962078, 4.961781, 4.963998, 4.966213, 4.96842, 4.970622, 
    4.972805, 4.974948, 4.977016, 4.978959, 4.98071, 4.982198, 4.983331, 
    4.98401, 4.984134, 4.9836, 4.982316, 4.980217, 4.977271, 4.973495, 
    4.968967,
  // totalHeight(27,48, 0-49)
    4.968221, 4.96867, 4.968932, 4.968997, 4.968864, 4.968532, 4.968005, 
    4.967294, 4.966412, 4.965373, 4.964195, 4.962899, 4.961504, 4.960023, 
    4.958469, 4.956077, 4.960622, 4.958631, 4.9565, 4.954679, 4.953285, 
    4.954834, 4.956685, 4.959286, 4.961421, 4.963017, 4.963776, 4.963808, 
    4.963056, 4.96275, 4.962512, 4.964767, 4.96697, 4.969106, 4.971163, 
    4.973114, 4.974928, 4.976556, 4.977943, 4.97902, 4.979716, 4.979949, 
    4.979635, 4.978698, 4.977073, 4.974717, 4.971618, 4.96781, 4.963374, 
    4.958452,
  // totalHeight(27,49, 0-49)
    4.964688, 4.965261, 4.965686, 4.965944, 4.966022, 4.965912, 4.965609, 
    4.96511, 4.964419, 4.963542, 4.962485, 4.96126, 4.959875, 4.958338, 
    4.95665, 4.953324, 4.963948, 4.960972, 4.957505, 4.954463, 4.952101, 
    4.95546, 4.959188, 4.964164, 4.967905, 4.970287, 4.97073, 4.969472, 
    4.966397, 4.964046, 4.961688, 4.964251, 4.966651, 4.968855, 4.970845, 
    4.972581, 4.974022, 4.975112, 4.975787, 4.975982, 4.975631, 4.974669, 
    4.973047, 4.97073, 4.967712, 4.964019, 4.959729, 4.954966, 4.949904, 
    4.944765,
  // totalHeight(28,0, 0-49)
    4.963037, 4.965694, 4.96799, 4.96993, 4.971521, 4.972774, 4.973701, 
    4.974322, 4.97466, 4.974749, 4.974625, 4.974331, 4.973917, 4.973434, 
    4.972936, 4.972286, 4.972091, 4.971761, 4.971567, 4.971555, 4.971744, 
    4.972298, 4.973012, 4.97391, 4.974973, 4.97617, 4.977477, 4.978871, 
    4.980332, 4.981852, 4.983389, 4.985156, 4.986973, 4.988846, 4.990781, 
    4.992773, 4.99481, 4.99686, 4.998869, 5.000762, 5.002431, 5.003738, 
    5.00451, 5.00454, 5.003603, 5.00145, 4.997844, 4.992567, 4.985462, 
    4.976461,
  // totalHeight(28,1, 0-49)
    4.964329, 4.966931, 4.969166, 4.971049, 4.972588, 4.973791, 4.974676, 
    4.975263, 4.975576, 4.975647, 4.975512, 4.975218, 4.974807, 4.97433, 
    4.973841, 4.973016, 4.97299, 4.972588, 4.972288, 4.972158, 4.972225, 
    4.97281, 4.973512, 4.974387, 4.975416, 4.976565, 4.977803, 4.979111, 
    4.980468, 4.981872, 4.983257, 4.985047, 4.986896, 4.988817, 4.990819, 
    4.992906, 4.995065, 4.997271, 4.999474, 5.001599, 5.003541, 5.005161, 
    5.006287, 5.006708, 5.006192, 5.004486, 5.001334, 4.996506, 4.989824, 
    4.981192,
  // totalHeight(28,2, 0-49)
    4.965621, 4.968162, 4.970339, 4.972167, 4.973656, 4.974818, 4.975669, 
    4.976233, 4.976532, 4.976597, 4.976467, 4.976181, 4.975784, 4.975326, 
    4.974851, 4.973862, 4.973973, 4.973501, 4.973098, 4.972849, 4.972789, 
    4.973388, 4.974058, 4.974888, 4.97586, 4.976943, 4.978105, 4.979328, 
    4.98059, 4.981882, 4.983115, 4.984918, 4.986787, 4.988737, 4.990783, 
    4.992933, 4.995179, 4.997493, 4.999833, 5.002124, 5.004266, 5.00612, 
    5.007517, 5.00825, 5.008084, 5.006764, 5.004031, 4.999646, 4.993412, 
    4.985214,
  // totalHeight(28,3, 0-49)
    4.966917, 4.969394, 4.971512, 4.973285, 4.974725, 4.975849, 4.976673, 
    4.977219, 4.97751, 4.977582, 4.977464, 4.977196, 4.976823, 4.976389, 
    4.975935, 4.974799, 4.974998, 4.974462, 4.973961, 4.973601, 4.973414, 
    4.97401, 4.974627, 4.975387, 4.976283, 4.977287, 4.978371, 4.979517, 
    4.980698, 4.981891, 4.98298, 4.984787, 4.986662, 4.988626, 4.990697, 
    4.992883, 4.995177, 4.997558, 4.999983, 5.002381, 5.004653, 5.00667, 
    5.008263, 5.009232, 5.009345, 5.008354, 5.006002, 5.002043, 4.996274, 
    4.988564,
  // totalHeight(28,4, 0-49)
    4.968223, 4.970632, 4.972686, 4.974402, 4.975794, 4.97688, 4.977679, 
    4.97821, 4.978501, 4.97858, 4.978481, 4.97824, 4.977897, 4.977489, 
    4.97706, 4.975801, 4.976025, 4.975429, 4.974844, 4.97438, 4.974075, 
    4.974649, 4.975199, 4.975864, 4.976665, 4.977577, 4.978583, 4.979664, 
    4.980787, 4.981899, 4.982858, 4.984657, 4.986529, 4.988494, 4.99057, 
    4.992767, 4.99508, 4.997489, 4.999952, 5.002404, 5.004749, 5.006863, 
    5.008582, 5.00972, 5.010053, 5.009339, 5.007329, 5.00378, 4.998486, 
    4.991301,
  // totalHeight(28,5, 0-49)
    4.969545, 4.971881, 4.973867, 4.975522, 4.976862, 4.977907, 4.978678, 
    4.979195, 4.979484, 4.979575, 4.979497, 4.979285, 4.978973, 4.978598, 
    4.978193, 4.976839, 4.977013, 4.976367, 4.975714, 4.975161, 4.97475, 
    4.975285, 4.975749, 4.976297, 4.976986, 4.977798, 4.978731, 4.979761, 
    4.980849, 4.981899, 4.982753, 4.984535, 4.986391, 4.988342, 4.990406, 
    4.992593, 4.994897, 4.997301, 4.999764, 5.002223, 5.00459, 5.006744, 
    5.008537, 5.009789, 5.010285, 5.009804, 5.008102, 5.004949, 5.000133, 
    4.993503,
  // totalHeight(28,6, 0-49)
    4.970886, 4.97314, 4.975051, 4.976639, 4.977922, 4.978922, 4.979661, 
    4.98016, 4.980445, 4.980545, 4.980488, 4.980305, 4.980027, 4.979684, 
    4.979302, 4.977885, 4.977926, 4.977243, 4.97654, 4.975917, 4.975418, 
    4.975897, 4.97626, 4.976669, 4.977231, 4.977938, 4.978801, 4.979794, 
    4.980872, 4.981885, 4.982657, 4.984412, 4.986242, 4.988164, 4.990201, 
    4.992358, 4.994633, 4.997004, 4.999434, 5.001863, 5.00421, 5.006363, 
    5.008183, 5.0095, 5.010123, 5.009836, 5.008419, 5.005644, 5.001309, 
    4.995253,
  // totalHeight(28,7, 0-49)
    4.97225, 4.974414, 4.976242, 4.977755, 4.978972, 4.979918, 4.980618, 
    4.981094, 4.98137, 4.981475, 4.981435, 4.981279, 4.981033, 4.980721, 
    4.98036, 4.978918, 4.978734, 4.978028, 4.977297, 4.976627, 4.976062, 
    4.976467, 4.976714, 4.976967, 4.977389, 4.977985, 4.978783, 4.979753, 
    4.980847, 4.981849, 4.982569, 4.984282, 4.986072, 4.987955, 4.989949, 
    4.992061, 4.994284, 4.996599, 4.998971, 5.001343, 5.003639, 5.005757, 
    5.007569, 5.008923, 5.00964, 5.009525, 5.00837, 5.005964, 5.002109, 
    4.996638,
  // totalHeight(28,8, 0-49)
    4.973632, 4.975698, 4.977432, 4.978859, 4.980003, 4.980888, 4.981541, 
    4.981984, 4.982244, 4.982347, 4.98232, 4.982186, 4.981969, 4.981684, 
    4.98134, 4.979915, 4.979413, 4.978697, 4.977963, 4.977275, 4.97667, 
    4.976981, 4.977097, 4.97718, 4.977454, 4.977934, 4.978669, 4.97963, 
    4.980763, 4.981778, 4.982479, 4.984136, 4.985872, 4.987704, 4.989642, 
    4.991693, 4.99385, 4.996092, 4.998385, 5.00068, 5.002903, 5.004966, 
    5.006748, 5.008116, 5.00891, 5.00895, 5.008045, 5.005998, 5.00262, 
    4.997739,
  // totalHeight(28,9, 0-49)
    4.975026, 4.976983, 4.978614, 4.979947, 4.981006, 4.98182, 4.982415, 
    4.982818, 4.983053, 4.983148, 4.983126, 4.983008, 4.982814, 4.982553, 
    4.982228, 4.980858, 4.979939, 4.979236, 4.978528, 4.977848, 4.977229, 
    4.97743, 4.977406, 4.977305, 4.977422, 4.977784, 4.978463, 4.979421, 
    4.980612, 4.981666, 4.98238, 4.983967, 4.985638, 4.987401, 4.989273, 
    4.991251, 4.993327, 4.995483, 4.997686, 4.999889, 5.002028, 5.004021, 
    5.005765, 5.007137, 5.007996, 5.008182, 5.00752, 5.005828, 5.002922, 
    4.998632,
  // totalHeight(28,10, 0-49)
    4.976417, 4.978255, 4.979773, 4.981001, 4.981967, 4.9827, 4.98323, 
    4.983584, 4.983787, 4.983865, 4.98384, 4.983733, 4.983557, 4.983315, 
    4.983003, 4.981734, 4.980297, 4.979631, 4.978978, 4.97834, 4.977737, 
    4.977809, 4.977633, 4.977343, 4.9773, 4.977544, 4.978166, 4.979129, 
    4.980392, 4.981504, 4.982268, 4.983768, 4.985357, 4.987044, 4.988835, 
    4.990729, 4.992716, 4.994777, 4.996881, 4.998987, 5.001035, 5.002955, 
    5.004656, 5.00603, 5.006954, 5.007286, 5.006864, 5.005523, 5.003084, 
    4.999376,
  // totalHeight(28,11, 0-49)
    4.977788, 4.979498, 4.980894, 4.982008, 4.982872, 4.983517, 4.983973, 
    4.984268, 4.984429, 4.984483, 4.984451, 4.984347, 4.984181, 4.983957, 
    4.983658, 4.98253, 4.980477, 4.979874, 4.979309, 4.978745, 4.978193, 
    4.978118, 4.977784, 4.977296, 4.977094, 4.977222, 4.97779, 4.978761, 
    4.980103, 4.981291, 4.982141, 4.983537, 4.985031, 4.986626, 4.988327, 
    4.990128, 4.992017, 4.993978, 4.995981, 4.997988, 4.999948, 5.001796, 
    5.00346, 5.004842, 5.005836, 5.006314, 5.006134, 5.005139, 5.003159, 
    5.000023,
  // totalHeight(28,12, 0-49)
    4.979121, 4.98069, 4.981956, 4.982948, 4.983704, 4.984252, 4.984627, 
    4.984859, 4.984973, 4.984995, 4.984945, 4.984837, 4.984681, 4.984471, 
    4.984189, 4.983234, 4.980469, 4.979962, 4.979518, 4.979064, 4.978595, 
    4.978358, 4.977861, 4.977178, 4.976821, 4.976835, 4.97735, 4.978325, 
    4.979751, 4.981029, 4.981995, 4.983273, 4.984656, 4.986147, 4.987747, 
    4.989446, 4.991234, 4.993092, 4.994994, 4.996906, 4.998783, 5.000571, 
    5.002206, 5.003607, 5.004677, 5.00531, 5.005374, 5.004723, 5.003193, 
    5.000611,
  // totalHeight(28,13, 0-49)
    4.980392, 4.981812, 4.982938, 4.983803, 4.984443, 4.98489, 4.985179, 
    4.985341, 4.985403, 4.985387, 4.985314, 4.985199, 4.985044, 4.984848, 
    4.984589, 4.983837, 4.980271, 4.979891, 4.979608, 4.979298, 4.978949, 
    4.978534, 4.977874, 4.977001, 4.976495, 4.976401, 4.976861, 4.977839, 
    4.979345, 4.980719, 4.981833, 4.982975, 4.984235, 4.98561, 4.987098, 
    4.988689, 4.990372, 4.992128, 4.993932, 4.995756, 4.997561, 4.999301, 
    5.00092, 5.002353, 5.003514, 5.00431, 5.004621, 5.004309, 5.003215, 
    5.001168,
  // totalHeight(28,14, 0-49)
    4.981575, 4.982839, 4.983819, 4.984552, 4.985072, 4.985415, 4.985616, 
    4.985703, 4.985707, 4.98565, 4.98555, 4.985421, 4.985268, 4.985085, 
    4.984856, 4.98433, 4.97988, 4.979667, 4.979576, 4.979448, 4.979251, 
    4.97865, 4.977829, 4.976778, 4.976137, 4.975942, 4.976348, 4.97732, 
    4.978895, 4.98037, 4.981659, 4.982649, 4.98377, 4.985018, 4.986386, 
    4.987864, 4.989438, 4.991094, 4.992805, 4.99455, 4.996294, 4.998002, 
    4.999622, 5.001102, 5.002368, 5.003336, 5.003896, 5.003918, 5.003249, 
    5.001713,
  // totalHeight(28,15, 0-49)
    4.982654, 4.983751, 4.984578, 4.985173, 4.985571, 4.985808, 4.985918, 
    4.98593, 4.985873, 4.985772, 4.985643, 4.985499, 4.985344, 4.985178, 
    4.984991, 4.984704, 4.979304, 4.979292, 4.979429, 4.979517, 4.979506, 
    4.978709, 4.977736, 4.976521, 4.975759, 4.975474, 4.975827, 4.976785, 
    4.978418, 4.979989, 4.981472, 4.982297, 4.983266, 4.984376, 4.985615, 
    4.986974, 4.988441, 4.989997, 4.991624, 4.993299, 4.994998, 4.996687, 
    4.998328, 4.999872, 5.001257, 5.002406, 5.003217, 5.003567, 5.003305, 
    5.002254,
  // totalHeight(28,16, 0-49)
    4.983608, 4.984528, 4.985196, 4.98565, 4.985922, 4.986052, 4.98607, 
    4.986007, 4.98589, 4.985743, 4.985583, 4.985423, 4.985268, 4.985124, 
    4.984986, 4.984951, 4.978553, 4.978775, 4.979172, 4.979506, 4.979712, 
    4.978718, 4.977604, 4.976244, 4.975379, 4.975018, 4.975318, 4.976254, 
    4.977931, 4.979589, 4.981279, 4.981926, 4.98273, 4.983689, 4.984793, 
    4.986029, 4.987384, 4.988845, 4.990394, 4.992012, 4.993679, 4.995368, 
    4.997046, 4.998671, 5.000189, 5.001527, 5.002593, 5.003264, 5.003393, 
    5.002801,
  // totalHeight(28,17, 0-49)
    4.984422, 4.985153, 4.985654, 4.985961, 4.986106, 4.986128, 4.986056, 
    4.985919, 4.985743, 4.985553, 4.985363, 4.985186, 4.985034, 4.984914, 
    4.984838, 4.985061, 4.977653, 4.978134, 4.978813, 4.97942, 4.979869, 
    4.978677, 4.977434, 4.975953, 4.975008, 4.974584, 4.974835, 4.975744, 
    4.977448, 4.979182, 4.981081, 4.981539, 4.982168, 4.982968, 4.983927, 
    4.985033, 4.986276, 4.987643, 4.98912, 4.990694, 4.992342, 4.994048, 
    4.995781, 4.997505, 4.999168, 5.000705, 5.002026, 5.00301, 5.003512, 
    5.003355,
  // totalHeight(28,18, 0-49)
    4.985089, 4.985617, 4.985938, 4.98609, 4.986105, 4.986018, 4.985858, 
    4.985652, 4.985424, 4.985193, 4.984977, 4.984787, 4.98464, 4.984551, 
    4.984545, 4.985033, 4.976648, 4.977406, 4.978383, 4.979276, 4.979985, 
    4.978594, 4.977239, 4.975657, 4.97465, 4.974179, 4.974391, 4.975267, 
    4.976982, 4.978776, 4.980881, 4.981141, 4.981584, 4.982214, 4.98302, 
    4.983992, 4.985119, 4.986394, 4.987806, 4.989342, 4.990986, 4.992723, 
    4.994529, 4.996365, 4.998188, 4.999933, 5.00151, 5.002803, 5.003664, 
    5.003913,
  // totalHeight(28,19, 0-49)
    4.985601, 4.985903, 4.986029, 4.986017, 4.985898, 4.985704, 4.985462, 
    4.985194, 4.98492, 4.984657, 4.984419, 4.984222, 4.984084, 4.984033, 
    4.984104, 4.984866, 4.975602, 4.976647, 4.977926, 4.979109, 4.980078, 
    4.978496, 4.977036, 4.975368, 4.974319, 4.973816, 4.973994, 4.974836, 
    4.976551, 4.978387, 4.980682, 4.980737, 4.980986, 4.981435, 4.982077, 
    4.982903, 4.983911, 4.985092, 4.986441, 4.987948, 4.989601, 4.991385, 
    4.993277, 4.995243, 4.997238, 4.999198, 5.001037, 5.002635, 5.003841, 
    5.004478,
  // totalHeight(28,20, 0-49)
    4.986712, 4.987498, 4.98811, 4.988571, 4.988906, 4.989136, 4.989282, 
    4.98936, 4.98939, 4.989389, 4.989371, 4.989356, 4.989365, 4.989432, 
    4.989607, 30, 4.973971, 4.974906, 4.976127, 4.977295, 4.978267, 4.976232, 
    4.974376, 4.972327, 4.970971, 4.970251, 4.970322, 4.971179, 4.973058, 
    4.975195, 4.977999, 4.978202, 4.978607, 4.979215, 4.980005, 4.980972, 
    4.982105, 4.983404, 4.984862, 4.986478, 4.988243, 4.990149, 4.992177, 
    4.994302, 4.996484, 4.998657, 5.000737, 5.002606, 5.004115, 5.005083,
  // totalHeight(28,21, 0-49)
    4.987054, 4.987665, 4.988129, 4.988471, 4.988711, 4.988868, 4.988958, 
    4.989, 4.989004, 4.988986, 4.988958, 4.988937, 4.988944, 4.989013, 
    4.989195, 30, 4.970282, 4.971366, 4.97281, 4.974231, 4.975453, 4.973234, 
    4.971309, 4.969253, 4.967992, 4.967446, 4.967751, 4.968876, 4.971061, 
    4.973518, 4.976734, 4.976965, 4.977419, 4.978096, 4.978973, 4.980039, 
    4.981282, 4.982694, 4.984271, 4.986003, 4.987885, 4.989907, 4.992052, 
    4.994292, 4.996589, 4.998882, 5.001087, 5.003087, 5.004737, 5.00586,
  // totalHeight(28,22, 0-49)
    4.987328, 4.98778, 4.988113, 4.988348, 4.988502, 4.988594, 4.988635, 
    4.98864, 4.988618, 4.988581, 4.988539, 4.988505, 4.988502, 4.988559, 
    4.988728, 30, 4.967324, 4.968526, 4.970151, 4.971785, 4.973213, 4.970802, 
    4.968777, 4.96666, 4.965425, 4.964967, 4.965406, 4.966697, 4.969078, 
    4.97174, 4.975243, 4.975431, 4.975869, 4.976557, 4.977474, 4.978605, 
    4.979939, 4.981463, 4.98317, 4.985048, 4.987089, 4.989276, 4.991593, 
    4.994008, 4.996481, 4.99895, 5.001328, 5.003502, 5.005326, 5.006629,
  // totalHeight(28,23, 0-49)
    4.987549, 4.987857, 4.98807, 4.988206, 4.988283, 4.988314, 4.98831, 
    4.988281, 4.988234, 4.988175, 4.988117, 4.988068, 4.988048, 4.988085, 
    4.988226, 30, 4.964871, 4.966145, 4.967893, 4.969668, 4.971232, 4.968641, 
    4.966502, 4.964304, 4.963049, 4.962618, 4.963121, 4.964503, 4.966997, 
    4.96978, 4.973461, 4.973578, 4.97397, 4.974645, 4.975582, 4.976766, 
    4.978186, 4.979832, 4.981688, 4.983741, 4.985978, 4.988378, 4.990917, 
    4.993559, 4.996259, 4.998947, 5.001537, 5.003915, 5.005933, 5.007423,
  // totalHeight(28,24, 0-49)
    4.98774, 4.98791, 4.988009, 4.988055, 4.98806, 4.988034, 4.987987, 
    4.987925, 4.987851, 4.987772, 4.987696, 4.987629, 4.987588, 4.987599, 
    4.987702, 30, 4.963188, 4.964485, 4.966293, 4.968147, 4.969785, 4.967083, 
    4.964877, 4.962627, 4.961349, 4.960917, 4.961437, 4.962847, 4.965379, 
    4.968204, 4.971961, 4.972018, 4.972366, 4.973018, 4.973957, 4.975173, 
    4.976654, 4.97839, 4.980366, 4.982566, 4.984974, 4.987565, 4.990309, 
    4.993167, 4.996087, 4.998994, 5.001799, 5.004381, 5.006594, 5.00827,
  // totalHeight(28,25, 0-49)
    4.987918, 4.987956, 4.987947, 4.987906, 4.98784, 4.98776, 4.987669, 
    4.987572, 4.98747, 4.98737, 4.987273, 4.987188, 4.987124, 4.987105, 
    4.987164, 30, 4.961998, 4.963271, 4.96508, 4.966942, 4.96859, 4.965873, 
    4.963664, 4.961417, 4.960142, 4.95971, 4.960229, 4.96163, 4.964145, 
    4.966951, 4.9707, 4.97073, 4.971062, 4.971709, 4.972658, 4.973903, 
    4.975436, 4.977246, 4.979321, 4.981645, 4.984196, 4.986951, 4.989874, 
    4.992926, 4.996044, 4.999156, 5.002161, 5.00494, 5.007341, 5.009192,
  // totalHeight(28,26, 0-49)
    4.988102, 4.988014, 4.9879, 4.98777, 4.987633, 4.987494, 4.987355, 
    4.987218, 4.987085, 4.986959, 4.98684, 4.986735, 4.98665, 4.986601, 
    4.986614, 30, 4.96127, 4.962483, 4.964233, 4.96604, 4.967638, 4.965005, 
    4.962867, 4.960688, 4.95945, 4.959028, 4.95953, 4.960891, 4.963342, 
    4.966077, 4.969729, 4.969779, 4.970129, 4.970798, 4.971775, 4.973054, 
    4.974634, 4.976504, 4.978654, 4.98107, 4.983733, 4.986615, 4.989684, 
    4.992893, 4.996181, 4.99947, 5.002655, 5.005613, 5.008188, 5.010205,
  // totalHeight(28,27, 0-49)
    4.988311, 4.988101, 4.987882, 4.987662, 4.987448, 4.987243, 4.987047, 
    4.986861, 4.986687, 4.986527, 4.986381, 4.986256, 4.986153, 4.986082, 
    4.986058, 30, 4.961052, 4.962173, 4.963817, 4.96551, 4.967003, 4.964544, 
    4.962538, 4.960472, 4.959287, 4.958868, 4.959324, 4.960605, 4.962934, 
    4.965534, 4.969001, 4.969101, 4.969494, 4.970201, 4.971213, 4.972528, 
    4.974146, 4.97606, 4.978265, 4.980749, 4.983495, 4.986478, 4.989666, 
    4.993008, 4.996446, 4.999894, 5.003249, 5.006377, 5.009121, 5.011301,
  // totalHeight(28,28, 0-49)
    4.988558, 4.98823, 4.987906, 4.987594, 4.987296, 4.987011, 4.986745, 
    4.986495, 4.986266, 4.986061, 4.985881, 4.985734, 4.98562, 4.985543, 
    4.985505, 30, 4.961629, 4.962648, 4.964153, 4.965688, 4.967029, 4.964806, 
    4.962961, 4.961018, 4.959865, 4.959403, 4.959753, 4.960879, 4.963003, 
    4.965382, 4.968564, 4.968718, 4.969153, 4.969889, 4.97092, 4.97225, 
    4.973881, 4.975813, 4.978045, 4.980568, 4.983372, 4.986431, 4.989717, 
    4.993181, 4.996759, 5.000366, 5.003891, 5.007196, 5.010116, 5.012463,
  // totalHeight(28,29, 0-49)
    4.988853, 4.988415, 4.987991, 4.98758, 4.987185, 4.986807, 4.986447, 
    4.986111, 4.985805, 4.985536, 4.985315, 4.985149, 4.985041, 4.984988, 
    4.984979, 30, 4.96272, 4.963651, 4.965005, 4.966348, 4.967486, 4.965503, 
    4.96379, 4.961924, 4.960732, 4.960146, 4.960302, 4.961183, 4.963007, 
    4.965075, 4.967861, 4.968034, 4.96848, 4.969221, 4.970254, 4.97159, 
    4.973233, 4.975191, 4.977465, 4.980054, 4.982945, 4.986122, 4.989549, 
    4.993178, 4.996941, 5.000747, 5.004481, 5.007996, 5.01112, 5.013654,
  // totalHeight(28,30, 0-49)
    4.98853, 4.987349, 4.986206, 4.985108, 4.984058, 4.983053, 4.98209, 
    4.981159, 4.980254, 4.979371, 4.978508, 4.977676, 4.976903, 4.976246, 
    4.975795, 4.974938, 4.965952, 4.966966, 4.968203, 4.969349, 4.970299, 
    4.968656, 4.967254, 4.965686, 4.964678, 4.964137, 4.964175, 4.964772, 
    4.966136, 4.967617, 4.969641, 4.969453, 4.969526, 4.969896, 4.970581, 
    4.971605, 4.972989, 4.974744, 4.976882, 4.979402, 4.982292, 4.98553, 
    4.989075, 4.992872, 4.996842, 5.000887, 5.004877, 5.008653, 5.012033, 
    5.014809,
  // totalHeight(28,31, 0-49)
    4.988934, 4.987695, 4.986489, 4.98532, 4.98419, 4.983098, 4.982041, 
    4.981017, 4.980021, 4.979056, 4.978122, 4.977229, 4.976397, 4.975665, 
    4.975098, 4.974432, 4.965597, 4.966311, 4.967228, 4.96806, 4.968717, 
    4.96726, 4.965956, 4.96447, 4.963483, 4.962937, 4.96296, 4.963528, 
    4.964809, 4.96617, 4.967934, 4.96792, 4.968172, 4.968722, 4.969593, 
    4.970803, 4.972375, 4.97432, 4.976649, 4.979359, 4.982438, 4.985861, 
    4.989586, 4.993555, 4.997685, 5.001874, 5.005987, 5.009863, 5.013318, 
    5.016133,
  // totalHeight(28,32, 0-49)
    4.989329, 4.988023, 4.986743, 4.985494, 4.984277, 4.983092, 4.98194, 
    4.980819, 4.979729, 4.978675, 4.977658, 4.976685, 4.97577, 4.974939, 
    4.974227, 4.97373, 4.965408, 4.965789, 4.966353, 4.966842, 4.96719, 
    4.965924, 4.964731, 4.963346, 4.9624, 4.961866, 4.961875, 4.962408, 
    4.963588, 4.964805, 4.966289, 4.966444, 4.96687, 4.967595, 4.96864, 
    4.970027, 4.971777, 4.973903, 4.976413, 4.979305, 4.982565, 4.986166, 
    4.990065, 4.994201, 4.998487, 5.002816, 5.007049, 5.011023, 5.014543, 
    5.017394,
  // totalHeight(28,33, 0-49)
    4.989703, 4.988327, 4.986968, 4.985633, 4.984324, 4.983045, 4.981792, 
    4.980573, 4.979386, 4.978236, 4.977127, 4.976064, 4.975055, 4.974112, 
    4.973249, 4.97283, 4.965299, 4.96534, 4.965545, 4.96569, 4.965733, 
    4.964666, 4.963603, 4.962349, 4.961465, 4.960958, 4.96096, 4.961446, 
    4.962501, 4.963549, 4.96474, 4.96506, 4.965649, 4.966537, 4.967746, 
    4.969299, 4.971216, 4.973511, 4.976191, 4.979255, 4.982684, 4.986455, 
    4.990518, 4.994809, 4.99924, 5.003698, 5.008042, 5.0121, 5.015676, 
    5.018547,
  // totalHeight(28,34, 0-49)
    4.990031, 4.988589, 4.987155, 4.985735, 4.984336, 4.982958, 4.981607, 
    4.980285, 4.978996, 4.977746, 4.976541, 4.975382, 4.974274, 4.973217, 
    4.972211, 4.971758, 4.965207, 4.964923, 4.964778, 4.964593, 4.964345, 
    4.963485, 4.962573, 4.961481, 4.960687, 4.960222, 4.960217, 4.960645, 
    4.961547, 4.962411, 4.963303, 4.963782, 4.964528, 4.965569, 4.966932, 
    4.96864, 4.970713, 4.973166, 4.976003, 4.979225, 4.982812, 4.986735, 
    4.990946, 4.995378, 4.999937, 5.004506, 5.008938, 5.013061, 5.01667, 
    5.019539,
  // totalHeight(28,35, 0-49)
    4.990283, 4.988789, 4.987288, 4.985792, 4.984304, 4.982832, 4.981381, 
    4.979957, 4.978567, 4.977216, 4.97591, 4.974653, 4.973446, 4.97228, 
    4.971144, 4.970554, 4.965104, 4.964519, 4.964046, 4.963553, 4.96304, 
    4.962392, 4.96165, 4.960749, 4.960071, 4.959666, 4.959654, 4.960008, 
    4.960733, 4.961397, 4.961999, 4.96263, 4.963524, 4.964712, 4.966218, 
    4.96807, 4.970286, 4.972882, 4.975864, 4.979228, 4.982954, 4.987012, 
    4.991352, 4.995899, 5.000561, 5.005215, 5.009709, 5.013865, 5.017476, 
    5.020309,
  // totalHeight(28,36, 0-49)
    4.990426, 4.988896, 4.987345, 4.985782, 4.984218, 4.982658, 4.981112, 
    4.97959, 4.9781, 4.976649, 4.975245, 4.973891, 4.972588, 4.971323, 
    4.970076, 4.969267, 4.964972, 4.964121, 4.963349, 4.962579, 4.961828, 
    4.961393, 4.960837, 4.960156, 4.959619, 4.959288, 4.959268, 4.959536, 
    4.960064, 4.96052, 4.960848, 4.961624, 4.962659, 4.963984, 4.965623, 
    4.967606, 4.969953, 4.972678, 4.975785, 4.979272, 4.983116, 4.987284, 
    4.991723, 4.996358, 5.001091, 5.005792, 5.010311, 5.014461, 5.01803, 
    5.020787,
  // totalHeight(28,37, 0-49)
    4.99042, 4.988878, 4.987295, 4.985683, 4.984055, 4.98242, 4.980792, 
    4.97918, 4.977595, 4.97605, 4.974551, 4.973106, 4.971712, 4.970358, 
    4.969019, 4.967945, 4.964811, 4.963729, 4.962691, 4.961675, 4.960719, 
    4.960494, 4.960138, 4.959701, 4.959327, 4.959084, 4.959058, 4.959228, 
    4.959541, 4.959791, 4.959871, 4.960784, 4.961951, 4.963401, 4.965164, 
    4.967265, 4.969728, 4.972565, 4.975777, 4.979362, 4.983298, 4.987546, 
    4.992053, 4.996737, 5.001498, 5.006205, 5.0107, 5.014793, 5.018272, 5.0209,
  // totalHeight(28,38, 0-49)
    4.99023, 4.988701, 4.987109, 4.98547, 4.983797, 4.982105, 4.980407, 
    4.978717, 4.977051, 4.97542, 4.973835, 4.972305, 4.97083, 4.969398, 
    4.967984, 4.966624, 4.964621, 4.963344, 4.962071, 4.960845, 4.959713, 
    4.959695, 4.959548, 4.959376, 4.959183, 4.959043, 4.959011, 4.959078, 
    4.959167, 4.959216, 4.959079, 4.960124, 4.961415, 4.962979, 4.964853, 
    4.967059, 4.969621, 4.972549, 4.975846, 4.979504, 4.983499, 4.98779, 
    4.992322, 4.997014, 5.001755, 5.006413, 5.010828, 5.014806, 5.018132, 
    5.020571,
  // totalHeight(28,39, 0-49)
    4.98982, 4.988333, 4.986758, 4.985115, 4.983422, 4.981692, 4.979945, 
    4.978195, 4.976461, 4.974759, 4.973101, 4.971496, 4.969948, 4.968448, 
    4.966973, 4.965341, 4.964407, 4.962965, 4.961492, 4.960084, 4.958814, 
    4.958994, 4.959059, 4.959167, 4.959174, 4.959148, 4.959116, 4.959077, 
    4.958942, 4.958804, 4.958484, 4.959653, 4.96106, 4.962731, 4.964701, 
    4.966998, 4.96964, 4.972637, 4.975991, 4.979691, 4.983709, 4.988005, 
    4.992517, 4.997162, 5.001826, 5.006374, 5.010642, 5.014437, 5.017542, 
    5.019726,
  // totalHeight(28,40, 0-49)
    4.989163, 4.987743, 4.986215, 4.984596, 4.982908, 4.981167, 4.979392, 
    4.977604, 4.975822, 4.974064, 4.972347, 4.970681, 4.969072, 4.967516, 
    4.965992, 4.964116, 4.964172, 4.962595, 4.960951, 4.959398, 4.958017, 
    4.958385, 4.958663, 4.959061, 4.959281, 4.959382, 4.959355, 4.959212, 
    4.958863, 4.958557, 4.95809, 4.959379, 4.960891, 4.962658, 4.964714, 
    4.967083, 4.969785, 4.972829, 4.97621, 4.979917, 4.983921, 4.988175, 
    4.992615, 4.997153, 5.001677, 5.006044, 5.010092, 5.013627, 5.016435, 
    5.018291,
  // totalHeight(28,41, 0-49)
    4.988236, 4.986912, 4.985459, 4.983894, 4.982239, 4.980513, 4.978737, 
    4.976935, 4.975128, 4.973335, 4.971576, 4.969865, 4.968209, 4.966607, 
    4.965042, 4.962963, 4.963916, 4.962226, 4.960443, 4.958775, 4.957313, 
    4.957856, 4.958346, 4.959037, 4.959479, 4.959718, 4.959705, 4.959471, 
    4.958921, 4.958473, 4.957899, 4.959299, 4.96091, 4.962762, 4.96489, 
    4.967316, 4.970056, 4.973118, 4.976497, 4.980174, 4.984117, 4.988278, 
    4.992589, 4.996957, 5.001267, 5.005378, 5.009124, 5.012317, 5.014746, 
    5.016197,
  // totalHeight(28,42, 0-49)
    4.98703, 4.98583, 4.984478, 4.982997, 4.981404, 4.979722, 4.977974, 
    4.976183, 4.974374, 4.97257, 4.97079, 4.96905, 4.96736, 4.965723, 
    4.964126, 4.961891, 4.963639, 4.961859, 4.95996, 4.958206, 4.956691, 
    4.957398, 4.958096, 4.959077, 4.959745, 4.96013, 4.960144, 4.959831, 
    4.959105, 4.958547, 4.957901, 4.959409, 4.961112, 4.963038, 4.965222, 
    4.967688, 4.970444, 4.973498, 4.976838, 4.980443, 4.98428, 4.988293, 
    4.992411, 4.996538, 5.000558, 5.00433, 5.007689, 5.010449, 5.012415, 
    5.013385,
  // totalHeight(28,43, 0-49)
    4.98554, 4.984489, 4.983268, 4.981898, 4.980398, 4.978789, 4.977099, 
    4.975349, 4.973565, 4.971771, 4.96999, 4.96824, 4.96653, 4.964868, 
    4.963245, 4.9609, 4.963339, 4.961486, 4.959499, 4.957683, 4.956139, 
    4.956997, 4.957892, 4.959154, 4.960049, 4.960588, 4.96064, 4.960272, 
    4.959402, 4.958764, 4.958083, 4.959694, 4.961483, 4.963474, 4.965702, 
    4.968185, 4.970934, 4.973947, 4.977213, 4.980706, 4.984384, 4.988188, 
    4.992046, 4.99586, 4.999508, 5.002852, 5.005733, 5.007973, 5.009391, 
    5.009803,
  // totalHeight(28,44, 0-49)
    4.983782, 4.982901, 4.981836, 4.980603, 4.979224, 4.977719, 4.976113, 
    4.974431, 4.972697, 4.970939, 4.969179, 4.967435, 4.965723, 4.964047, 
    4.962406, 4.959991, 4.963014, 4.961103, 4.959048, 4.957194, 4.955643, 
    4.956639, 4.95772, 4.959247, 4.960364, 4.961061, 4.961168, 4.960768, 
    4.95979, 4.959107, 4.958425, 4.960135, 4.962002, 4.964049, 4.966306, 
    4.968788, 4.971504, 4.974445, 4.977598, 4.980931, 4.984395, 4.987931, 
    4.991458, 4.994877, 4.99807, 5.000897, 5.003209, 5.00484, 5.005627, 
    5.005414,
  // totalHeight(28,45, 0-49)
    4.981774, 4.981083, 4.980196, 4.979126, 4.977894, 4.97652, 4.975028, 
    4.973438, 4.971782, 4.970082, 4.968363, 4.966645, 4.964943, 4.963265, 
    4.961613, 4.959162, 4.962658, 4.960703, 4.958603, 4.956729, 4.955187, 
    4.956307, 4.957557, 4.959331, 4.960659, 4.961514, 4.961693, 4.961289, 
    4.960246, 4.959553, 4.958898, 4.960707, 4.962646, 4.964738, 4.967009, 
    4.969471, 4.972126, 4.974962, 4.977961, 4.981081, 4.984278, 4.987478, 
    4.990602, 4.993547, 4.996198, 4.998419, 5.000072, 5.001008, 5.001089, 
    5.000189,
  // totalHeight(28,46, 0-49)
    4.979548, 4.979063, 4.978371, 4.977488, 4.976427, 4.975208, 4.973854, 
    4.972385, 4.970828, 4.969208, 4.96755, 4.965873, 4.964198, 4.96253, 
    4.960874, 4.958412, 4.962271, 4.960286, 4.958158, 4.95628, 4.95476, 
    4.955986, 4.957387, 4.959378, 4.960902, 4.961915, 4.96218, 4.961805, 
    4.96074, 4.960072, 4.959472, 4.961374, 4.96338, 4.965507, 4.967777, 
    4.970197, 4.972763, 4.975461, 4.978261, 4.981122, 4.983987, 4.986786, 
    4.989431, 4.991823, 4.993845, 4.995374, 4.996282, 4.996446, 4.995755, 
    4.994122,
  // totalHeight(28,47, 0-49)
    4.977147, 4.976876, 4.976397, 4.975716, 4.974848, 4.973806, 4.972611, 
    4.971286, 4.96985, 4.968332, 4.966752, 4.965134, 4.963496, 4.961848, 
    4.960196, 4.957739, 4.96185, 4.959847, 4.957707, 4.955839, 4.95435, 
    4.955663, 4.957192, 4.959366, 4.961065, 4.962229, 4.962596, 4.962281, 
    4.96124, 4.96063, 4.960107, 4.962099, 4.964166, 4.966316, 4.96857, 
    4.970924, 4.973373, 4.975894, 4.978453, 4.981, 4.983474, 4.985802, 
    4.987894, 4.98965, 4.990963, 4.991716, 4.991806, 4.991132, 4.989618, 
    4.987222,
  // totalHeight(28,48, 0-49)
    4.974618, 4.974567, 4.974308, 4.973845, 4.973186, 4.972341, 4.971326, 
    4.970162, 4.968867, 4.967466, 4.965981, 4.964435, 4.962846, 4.961228, 
    4.959587, 4.957145, 4.961398, 4.959391, 4.957252, 4.9554, 4.953947, 
    4.955328, 4.956959, 4.959277, 4.961123, 4.962427, 4.962908, 4.962682, 
    4.96171, 4.961189, 4.960761, 4.962839, 4.964956, 4.967119, 4.969338, 
    4.971605, 4.973905, 4.976213, 4.978484, 4.980662, 4.982685, 4.984473, 
    4.98594, 4.986984, 4.987511, 4.987416, 4.986622, 4.985056, 4.982687, 
    4.979521,
  // totalHeight(28,49, 0-49)
    4.971751, 4.97187, 4.971794, 4.971513, 4.971032, 4.970352, 4.969482, 
    4.968434, 4.96722, 4.965861, 4.964369, 4.962768, 4.961073, 4.959293, 
    4.957433, 4.953966, 4.963982, 4.960976, 4.957507, 4.954463, 4.952083, 
    4.955269, 4.95878, 4.963472, 4.966963, 4.969119, 4.969381, 4.967987, 
    4.964842, 4.962405, 4.959975, 4.962437, 4.964849, 4.967206, 4.969516, 
    4.971771, 4.973949, 4.976017, 4.977924, 4.979613, 4.981015, 4.982051, 
    4.98264, 4.982693, 4.982131, 4.980882, 4.978908, 4.976194, 4.972773, 
    4.968725,
  // totalHeight(29,0, 0-49)
    4.971556, 4.973361, 4.974815, 4.975937, 4.976742, 4.97725, 4.977488, 
    4.977488, 4.977288, 4.976929, 4.976456, 4.97591, 4.975338, 4.97478, 
    4.974274, 4.973676, 4.973505, 4.973238, 4.973083, 4.97306, 4.973165, 
    4.973533, 4.973971, 4.974497, 4.975105, 4.975779, 4.976512, 4.977307, 
    4.978165, 4.979098, 4.980094, 4.981372, 4.982794, 4.984384, 4.986169, 
    4.988163, 4.99037, 4.992781, 4.995366, 4.998078, 5.000845, 5.003565, 
    5.00611, 5.008316, 5.009995, 5.010931, 5.010883, 5.009605, 5.006854, 
    5.002412,
  // totalHeight(29,1, 0-49)
    4.97285, 4.9746, 4.976003, 4.977079, 4.977844, 4.97832, 4.978535, 
    4.978521, 4.978314, 4.977955, 4.977486, 4.976948, 4.976385, 4.975832, 
    4.975327, 4.974553, 4.974493, 4.974136, 4.97386, 4.973703, 4.973669, 
    4.97404, 4.974442, 4.974925, 4.975485, 4.976109, 4.976785, 4.977513, 
    4.978296, 4.979141, 4.980009, 4.981315, 4.982766, 4.984389, 4.986212, 
    4.988253, 4.990514, 4.992992, 4.995659, 4.998469, 5.001352, 5.00421, 
    5.006918, 5.009318, 5.011222, 5.012416, 5.012663, 5.011715, 5.009322, 
    5.005255,
  // totalHeight(29,2, 0-49)
    4.974152, 4.975846, 4.977199, 4.978231, 4.97896, 4.979407, 4.979604, 
    4.979578, 4.979369, 4.979012, 4.978549, 4.978021, 4.977464, 4.976915, 
    4.976405, 4.97546, 4.975474, 4.975027, 4.974627, 4.974336, 4.974163, 
    4.974525, 4.97488, 4.975307, 4.975816, 4.976388, 4.977014, 4.977693, 
    4.978423, 4.979195, 4.979949, 4.981287, 4.982766, 4.984417, 4.986269, 
    4.988337, 4.990631, 4.993144, 4.995852, 4.998711, 5.001653, 5.004588, 
    5.007389, 5.009909, 5.011964, 5.013349, 5.013828, 5.013155, 5.011086, 
    5.007389,
  // totalHeight(29,3, 0-49)
    4.975455, 4.977093, 4.978398, 4.979385, 4.98008, 4.980501, 4.980679, 
    4.980646, 4.980434, 4.980083, 4.979627, 4.979106, 4.978555, 4.978006, 
    4.977489, 4.976379, 4.976416, 4.975876, 4.975358, 4.974937, 4.97463, 
    4.974973, 4.975272, 4.975631, 4.976077, 4.976596, 4.977183, 4.977833, 
    4.978536, 4.979261, 4.979921, 4.981289, 4.982796, 4.98447, 4.98634, 
    4.988424, 4.990729, 4.993248, 4.995963, 4.998829, 5.001781, 5.004733, 
    5.007569, 5.010144, 5.012286, 5.013795, 5.014449, 5.014008, 5.01223, 
    5.008885,
  // totalHeight(29,4, 0-49)
    4.976765, 4.978344, 4.979596, 4.980538, 4.981195, 4.981589, 4.981749, 
    4.981706, 4.981493, 4.981143, 4.980695, 4.980181, 4.979634, 4.979084, 
    4.978553, 4.977294, 4.977292, 4.976662, 4.976037, 4.975495, 4.975061, 
    4.975371, 4.975604, 4.975881, 4.976256, 4.976723, 4.97728, 4.97792, 
    4.978625, 4.979328, 4.979919, 4.98132, 4.982853, 4.984545, 4.986426, 
    4.988512, 4.990811, 4.993315, 4.996003, 4.99884, 5.00176, 5.004683, 
    5.0075, 5.010075, 5.012246, 5.013824, 5.0146, 5.014348, 5.012831, 5.009826,
  // totalHeight(29,5, 0-49)
    4.978075, 4.97959, 4.980784, 4.981678, 4.982295, 4.98266, 4.9828, 
    4.982745, 4.982529, 4.982182, 4.981737, 4.981228, 4.980682, 4.980126, 
    4.979578, 4.978192, 4.978077, 4.977365, 4.976644, 4.975996, 4.975449, 
    4.975712, 4.975867, 4.976048, 4.976345, 4.976757, 4.977293, 4.977944, 
    4.978681, 4.97939, 4.979939, 4.981371, 4.982926, 4.984634, 4.986518, 
    4.988595, 4.990872, 4.99334, 4.995981, 4.998755, 5.001609, 5.004463, 
    5.007217, 5.009746, 5.0119, 5.013502, 5.014358, 5.014255, 5.012973, 
    5.010293,
  // totalHeight(29,6, 0-49)
    4.979375, 4.980821, 4.981953, 4.982794, 4.983367, 4.983699, 4.983816, 
    4.983747, 4.983525, 4.983177, 4.982736, 4.982229, 4.981682, 4.981119, 
    4.980551, 4.979065, 4.978755, 4.977969, 4.97717, 4.976434, 4.975792, 
    4.975995, 4.976058, 4.976129, 4.976338, 4.976693, 4.977218, 4.977898, 
    4.978695, 4.979438, 4.979978, 4.981435, 4.98301, 4.984728, 4.986608, 
    4.988667, 4.990908, 4.993323, 4.995894, 4.998584, 5.00134, 5.004094, 
    5.006751, 5.009197, 5.011295, 5.012885, 5.013788, 5.013808, 5.012739, 
    5.010373,
  // totalHeight(29,7, 0-49)
    4.980656, 4.982026, 4.983089, 4.983871, 4.984396, 4.98469, 4.984782, 
    4.984697, 4.984466, 4.984116, 4.983675, 4.98317, 4.982621, 4.982047, 
    4.981458, 4.979904, 4.979315, 4.978468, 4.977612, 4.976809, 4.976092, 
    4.976218, 4.97618, 4.976123, 4.976236, 4.976532, 4.977053, 4.977777, 
    4.978659, 4.979466, 4.980029, 4.981503, 4.983092, 4.984814, 4.986686, 
    4.988718, 4.99091, 4.993259, 4.995742, 4.998327, 5.000965, 5.003592, 
    5.006126, 5.008463, 5.010478, 5.012031, 5.012955, 5.013077, 5.012204, 
    5.010143,
  // totalHeight(29,8, 0-49)
    4.981897, 4.983184, 4.984174, 4.984893, 4.985365, 4.98562, 4.985681, 
    4.985578, 4.985337, 4.984982, 4.984541, 4.984036, 4.983485, 4.982903, 
    4.982292, 4.980708, 4.979747, 4.978858, 4.977969, 4.977125, 4.976357, 
    4.976388, 4.976235, 4.976039, 4.976047, 4.976282, 4.976804, 4.977584, 
    4.978576, 4.979469, 4.980087, 4.981573, 4.983167, 4.984883, 4.986736, 
    4.988731, 4.990869, 4.993138, 4.99552, 4.997984, 5.000488, 5.002973, 
    5.005363, 5.007573, 5.009488, 5.010984, 5.011919, 5.012128, 5.011442, 
    5.009677,
  // totalHeight(29,9, 0-49)
    4.983086, 4.984283, 4.985192, 4.985842, 4.986258, 4.986469, 4.986499, 
    4.986375, 4.986122, 4.985764, 4.985322, 4.984818, 4.984266, 4.983675, 
    4.983043, 4.981473, 4.980051, 4.97914, 4.978247, 4.977389, 4.976596, 
    4.976516, 4.976236, 4.97589, 4.975786, 4.975957, 4.976483, 4.977327, 
    4.978443, 4.979445, 4.980153, 4.981635, 4.983224, 4.984926, 4.986752, 
    4.988701, 4.990771, 4.992952, 4.995222, 4.997556, 4.999913, 5.002243, 
    5.004482, 5.006552, 5.008358, 5.009792, 5.010726, 5.011018, 5.010513, 
    5.009043,
  // totalHeight(29,10, 0-49)
    4.984201, 4.9853, 4.986125, 4.986701, 4.987059, 4.987222, 4.987219, 
    4.987072, 4.986808, 4.986445, 4.986005, 4.985502, 4.984953, 4.984358, 
    4.983712, 4.982196, 4.980223, 4.979319, 4.978451, 4.977612, 4.976825, 
    4.976614, 4.976199, 4.975692, 4.975474, 4.975579, 4.976107, 4.977016, 
    4.978267, 4.979397, 4.980227, 4.981689, 4.983257, 4.984932, 4.986719, 
    4.988612, 4.990606, 4.992688, 4.99484, 4.997035, 4.99924, 5.001411, 
    5.003496, 5.005424, 5.007121, 5.008492, 5.009428, 5.009802, 5.009476, 
    5.008297,
  // totalHeight(29,11, 0-49)
    4.985221, 4.986217, 4.986951, 4.987451, 4.987747, 4.987863, 4.987825, 
    4.987659, 4.987381, 4.987016, 4.986578, 4.986081, 4.985535, 4.984943, 
    4.984293, 4.982874, 4.980265, 4.979398, 4.978592, 4.977806, 4.977054, 
    4.9767, 4.976141, 4.975471, 4.975133, 4.975172, 4.9757, 4.976673, 
    4.978061, 4.979329, 4.980305, 4.981731, 4.983263, 4.984897, 4.98663, 
    4.988455, 4.990363, 4.992339, 4.994365, 4.996418, 4.998469, 5.000483, 
    5.002415, 5.004209, 5.005803, 5.007117, 5.008061, 5.008524, 5.008382, 
    5.00749,
  // totalHeight(29,12, 0-49)
    4.986129, 4.987016, 4.987657, 4.988077, 4.98831, 4.988379, 4.988306, 
    4.988117, 4.987829, 4.987461, 4.98703, 4.986541, 4.986005, 4.985423, 
    4.984781, 4.983505, 4.980176, 4.979388, 4.978679, 4.977983, 4.977303, 
    4.976789, 4.976083, 4.975247, 4.974793, 4.974764, 4.975285, 4.976314, 
    4.977836, 4.979246, 4.980394, 4.981762, 4.983236, 4.98481, 4.986475, 
    4.98822, 4.99003, 4.991893, 4.99379, 4.9957, 4.997602, 4.999462, 5.00125, 
    5.002921, 5.004425, 5.005697, 5.00666, 5.007222, 5.007267, 5.006666,
  // totalHeight(29,13, 0-49)
    4.98691, 4.987683, 4.988225, 4.988565, 4.988734, 4.988751, 4.988646, 
    4.988435, 4.988138, 4.98777, 4.987345, 4.98687, 4.986352, 4.985789, 
    4.985172, 4.984077, 4.97996, 4.979289, 4.978722, 4.978153, 4.97758, 
    4.976897, 4.976046, 4.975048, 4.974481, 4.974383, 4.974892, 4.975965, 
    4.977607, 4.979157, 4.980497, 4.98178, 4.983175, 4.984669, 4.986247, 
    4.987896, 4.989599, 4.991342, 4.993107, 4.994876, 4.996633, 4.998353, 
    5.000012, 5.001576, 5.003008, 5.004256, 5.005257, 5.005929, 5.00617, 
    5.005861,
  // totalHeight(29,14, 0-49)
    4.987552, 4.988207, 4.988649, 4.988905, 4.989006, 4.988974, 4.988832, 
    4.988601, 4.988295, 4.987929, 4.987513, 4.987056, 4.986562, 4.986031, 
    4.985457, 4.984582, 4.97962, 4.979108, 4.978724, 4.978326, 4.977896, 
    4.977039, 4.976047, 4.974896, 4.974222, 4.974059, 4.974547, 4.975648, 
    4.977391, 4.979072, 4.980613, 4.981785, 4.983075, 4.984465, 4.985938, 
    4.987476, 4.989061, 4.990677, 4.992309, 4.993942, 4.995565, 4.997159, 
    4.998707, 5.000188, 5.001571, 5.002817, 5.003875, 5.004673, 5.00512, 
    5.005102,
  // totalHeight(29,15, 0-49)
    4.988047, 4.988579, 4.988916, 4.989087, 4.989118, 4.989033, 4.988854, 
    4.988601, 4.988286, 4.987922, 4.98752, 4.987084, 4.986623, 4.986136, 
    4.985628, 4.985004, 4.979161, 4.978853, 4.978694, 4.978505, 4.978258, 
    4.977225, 4.976098, 4.97481, 4.974041, 4.973814, 4.974275, 4.975384, 
    4.977204, 4.978997, 4.980742, 4.981776, 4.982933, 4.984197, 4.985542, 
    4.986952, 4.988406, 4.989891, 4.991391, 4.992896, 4.994396, 4.995882, 
    4.997343, 4.998764, 5.000125, 5.001397, 5.002533, 5.003475, 5.004138, 
    5.004411,
  // totalHeight(29,16, 0-49)
    4.988392, 4.988796, 4.989022, 4.989101, 4.98906, 4.98892, 4.988703, 
    4.988425, 4.988101, 4.987741, 4.987353, 4.986944, 4.986523, 4.986093, 
    4.985668, 4.985326, 4.978594, 4.978531, 4.978637, 4.978697, 4.978667, 
    4.977459, 4.976213, 4.974801, 4.973953, 4.973667, 4.974092, 4.975191, 
    4.977059, 4.978941, 4.980883, 4.98175, 4.982749, 4.983858, 4.985055, 
    4.986319, 4.987631, 4.988978, 4.990348, 4.991733, 4.993127, 4.994525, 
    4.995924, 4.997314, 4.998682, 5.000005, 5.001247, 5.002351, 5.00324, 
    5.003806,
  // totalHeight(29,17, 0-49)
    4.988588, 4.988854, 4.988962, 4.988945, 4.988825, 4.988625, 4.988366, 
    4.988063, 4.987727, 4.98737, 4.986999, 4.986622, 4.986247, 4.985889, 
    4.985566, 4.98553, 4.977942, 4.97816, 4.978563, 4.978907, 4.979125, 
    4.977752, 4.9764, 4.974884, 4.973968, 4.973629, 4.97401, 4.97508, 
    4.976967, 4.978909, 4.981034, 4.981708, 4.982517, 4.983448, 4.984474, 
    4.985574, 4.986732, 4.987938, 4.98918, 4.990454, 4.991757, 4.99309, 
    4.994452, 4.995841, 4.997247, 4.998652, 5.000022, 5.001309, 5.002435, 
    5.003295,
  // totalHeight(29,18, 0-49)
    4.988639, 4.988755, 4.988736, 4.98861, 4.988406, 4.988142, 4.987838, 
    4.987507, 4.987159, 4.986805, 4.986453, 4.986112, 4.985792, 4.985513, 
    4.98531, 4.985602, 4.977243, 4.977769, 4.978495, 4.979146, 4.979639, 
    4.978107, 4.976663, 4.97506, 4.974088, 4.973702, 4.974034, 4.975058, 
    4.976934, 4.978906, 4.981187, 4.981641, 4.982238, 4.982964, 4.983794, 
    4.984714, 4.985708, 4.986764, 4.987881, 4.989054, 4.990283, 4.991574, 
    4.992928, 4.994346, 4.995821, 4.997337, 4.998865, 5.000354, 5.001728, 
    5.002884,
  // totalHeight(29,19, 0-49)
    4.98855, 4.988499, 4.988338, 4.988094, 4.987796, 4.987462, 4.987109, 
    4.986747, 4.986388, 4.986039, 4.985707, 4.985406, 4.985149, 4.984963, 
    4.984892, 4.98553, 4.976555, 4.977411, 4.978475, 4.979445, 4.980222, 
    4.978542, 4.977019, 4.975341, 4.974323, 4.973892, 4.974168, 4.975128, 
    4.976965, 4.978934, 4.981341, 4.981552, 4.981909, 4.982407, 4.983021, 
    4.98374, 4.984555, 4.985459, 4.98645, 4.98753, 4.988702, 4.989972, 
    4.991343, 4.99282, 4.994395, 4.996053, 4.997765, 4.999477, 5.001114, 
    5.002572,
  // totalHeight(29,20, 0-49)
    4.989048, 4.989503, 4.989847, 4.990098, 4.99027, 4.990378, 4.990433, 
    4.990442, 4.990415, 4.99036, 4.990286, 4.990209, 4.990146, 4.990134, 
    4.990227, 30, 4.975359, 4.976153, 4.977207, 4.978203, 4.979018, 4.976952, 
    4.975087, 4.973069, 4.971763, 4.971109, 4.97125, 4.972173, 4.974099, 
    4.976275, 4.979077, 4.979346, 4.979769, 4.980332, 4.98101, 4.981788, 
    4.982655, 4.983606, 4.984644, 4.985774, 4.987006, 4.988348, 4.98981, 
    4.991399, 4.993111, 4.994935, 4.996837, 4.99877, 5.000656, 5.002386,
  // totalHeight(29,21, 0-49)
    4.988827, 4.98916, 4.989402, 4.98957, 4.989676, 4.989734, 4.989754, 
    4.989744, 4.989711, 4.98966, 4.9896, 4.989542, 4.989507, 4.989525, 
    4.989647, 30, 4.972302, 4.973264, 4.974558, 4.975825, 4.976907, 4.974704, 
    4.972797, 4.970784, 4.969567, 4.96906, 4.969389, 4.970522, 4.972679, 
    4.975086, 4.978195, 4.978409, 4.978792, 4.979332, 4.980003, 4.980789, 
    4.981676, 4.98266, 4.983741, 4.984922, 4.986211, 4.987618, 4.989153, 
    4.990819, 4.992617, 4.994532, 4.996534, 4.998575, 5.000577, 5.002439,
  // totalHeight(29,22, 0-49)
    4.988561, 4.988786, 4.988936, 4.989029, 4.989077, 4.989089, 4.989075, 
    4.989043, 4.988997, 4.988944, 4.988889, 4.988842, 4.988819, 4.988848, 
    4.988978, 30, 4.970036, 4.971129, 4.972622, 4.974118, 4.975419, 4.973063, 
    4.971076, 4.969011, 4.967807, 4.967357, 4.967772, 4.969004, 4.971275, 
    4.973795, 4.977079, 4.977161, 4.977431, 4.977885, 4.978497, 4.979252, 
    4.980139, 4.981151, 4.982288, 4.983549, 4.98494, 4.986465, 4.988132, 
    4.989944, 4.991897, 4.993972, 4.996139, 4.998345, 5.000515, 5.002546,
  // totalHeight(29,23, 0-49)
    4.988266, 4.988394, 4.988463, 4.988487, 4.988479, 4.988449, 4.988403, 
    4.988348, 4.988288, 4.988229, 4.988175, 4.988132, 4.988114, 4.988146, 
    4.988268, 30, 4.968285, 4.969466, 4.971102, 4.972762, 4.974215, 4.971715, 
    4.969638, 4.967495, 4.966257, 4.9658, 4.966229, 4.967482, 4.969783, 
    4.972326, 4.975673, 4.975587, 4.97571, 4.976046, 4.976573, 4.977282, 
    4.978163, 4.979208, 4.980416, 4.981785, 4.983315, 4.985008, 4.986862, 
    4.988875, 4.991038, 4.993327, 4.995707, 4.998123, 5.000495, 5.002719,
  // totalHeight(29,24, 0-49)
    4.987961, 4.987996, 4.987988, 4.98795, 4.987892, 4.987821, 4.987746, 
    4.98767, 4.987597, 4.987533, 4.987478, 4.987438, 4.987423, 4.987453, 
    4.987559, 30, 4.967278, 4.968503, 4.970228, 4.971992, 4.973543, 4.970967, 
    4.968838, 4.966646, 4.96537, 4.964878, 4.96527, 4.966482, 4.968736, 
    4.971223, 4.974539, 4.974289, 4.974264, 4.97447, 4.974896, 4.975535, 
    4.976382, 4.977432, 4.978685, 4.980134, 4.981779, 4.98362, 4.985648, 
    4.987854, 4.990224, 4.992731, 4.995331, 4.997964, 5.000548, 5.002974,
  // totalHeight(29,25, 0-49)
    4.98766, 4.987607, 4.987528, 4.98743, 4.987325, 4.987216, 4.987114, 
    4.987021, 4.986938, 4.986869, 4.986818, 4.986785, 4.986776, 4.986806, 
    4.986895, 30, 4.966704, 4.967937, 4.969695, 4.971504, 4.973098, 4.970532, 
    4.968414, 4.966226, 4.964935, 4.964411, 4.964749, 4.965886, 4.968045, 
    4.970422, 4.973626, 4.973247, 4.973096, 4.973194, 4.973528, 4.974099, 
    4.974905, 4.975947, 4.977223, 4.97873, 4.980465, 4.982426, 4.984601, 
    4.986979, 4.989538, 4.992245, 4.995053, 4.997897, 5.000687, 5.003313,
  // totalHeight(29,26, 0-49)
    4.987382, 4.987242, 4.987093, 4.986938, 4.986787, 4.986643, 4.986514, 
    4.986403, 4.986313, 4.986247, 4.986204, 4.986186, 4.986193, 4.986231, 
    4.986312, 30, 4.966497, 4.967708, 4.969454, 4.971251, 4.972836, 4.970378, 
    4.968344, 4.96622, 4.96495, 4.964405, 4.96468, 4.965718, 4.967741, 
    4.969964, 4.972982, 4.972522, 4.972288, 4.972305, 4.972567, 4.97308, 
    4.973845, 4.974867, 4.976147, 4.977685, 4.979478, 4.981522, 4.983808, 
    4.986319, 4.989032, 4.991911, 4.994902, 4.997937, 5.000921, 5.003737,
  // totalHeight(29,27, 0-49)
    4.987139, 4.986915, 4.986696, 4.986484, 4.986285, 4.986104, 4.98595, 
    4.985823, 4.985728, 4.985668, 4.985642, 4.98565, 4.985687, 4.985753, 
    4.985845, 30, 4.966663, 4.967835, 4.969529, 4.971269, 4.972798, 4.970535, 
    4.968647, 4.966635, 4.965405, 4.964836, 4.965031, 4.96594, 4.967781, 
    4.969799, 4.972559, 4.972056, 4.971772, 4.971733, 4.971939, 4.972399, 
    4.97312, 4.974112, 4.975377, 4.97692, 4.978742, 4.980838, 4.983202, 
    4.985818, 4.98866, 4.991688, 4.994846, 4.998058, 5.001228, 5.00423,
  // totalHeight(29,28, 0-49)
    4.986944, 4.986639, 4.986349, 4.986075, 4.985826, 4.985606, 4.985421, 
    4.985277, 4.985176, 4.985127, 4.985129, 4.985179, 4.985272, 4.985394, 
    4.985533, 30, 4.967456, 4.968589, 4.970207, 4.971852, 4.973289, 4.971285, 
    4.969576, 4.967695, 4.966493, 4.965866, 4.965929, 4.966646, 4.968236, 
    4.969983, 4.972405, 4.971874, 4.97155, 4.971457, 4.971603, 4.971999, 
    4.97266, 4.973596, 4.97482, 4.976341, 4.978161, 4.980283, 4.982701, 
    4.985398, 4.98835, 4.991515, 4.994833, 4.998222, 5.001579, 5.004774,
  // totalHeight(29,29, 0-49)
    4.986812, 4.986425, 4.986062, 4.985725, 4.98542, 4.985151, 4.984928, 
    4.984759, 4.984652, 4.984617, 4.984658, 4.984773, 4.984951, 4.985173, 
    4.985413, 30, 4.968573, 4.969682, 4.971219, 4.972744, 4.974048, 4.972317, 
    4.970768, 4.968982, 4.967752, 4.967, 4.966858, 4.967312, 4.968576, 
    4.969975, 4.971971, 4.971394, 4.971013, 4.970857, 4.970938, 4.971271, 
    4.971876, 4.97277, 4.97397, 4.975489, 4.977334, 4.979512, 4.982013, 
    4.984826, 4.987921, 4.991253, 4.994759, 4.998352, 5.001921, 5.005327,
  // totalHeight(29,30, 0-49)
    4.986113, 4.985028, 4.983992, 4.98301, 4.982088, 4.981229, 4.980436, 
    4.979713, 4.979061, 4.978491, 4.978013, 4.977649, 4.977439, 4.977439, 
    4.97774, 4.978108, 4.970986, 4.972597, 4.974332, 4.975877, 4.977121, 
    4.975759, 4.974507, 4.972983, 4.97189, 4.971142, 4.970854, 4.971008, 
    4.971807, 4.972627, 4.973881, 4.972935, 4.972168, 4.971625, 4.971332, 
    4.971322, 4.971624, 4.972265, 4.973269, 4.974652, 4.976425, 4.978588, 
    4.981136, 4.984048, 4.987289, 4.990808, 4.994532, 4.998365, 5.002188, 
    5.005852,
  // totalHeight(29,31, 0-49)
    4.986139, 4.985011, 4.983933, 4.982914, 4.981956, 4.981061, 4.980238, 
    4.979491, 4.978826, 4.978252, 4.977779, 4.977426, 4.97722, 4.9772, 
    4.977429, 4.977726, 4.970573, 4.971944, 4.973413, 4.974692, 4.97569, 
    4.974526, 4.973392, 4.971966, 4.970906, 4.970163, 4.969861, 4.969983, 
    4.970693, 4.971382, 4.972375, 4.971571, 4.970947, 4.970544, 4.970392, 
    4.970518, 4.970953, 4.971724, 4.972854, 4.974358, 4.976247, 4.978524, 
    4.98118, 4.984198, 4.987542, 4.991161, 4.99498, 4.998902, 5.002809, 
    5.006545,
  // totalHeight(29,32, 0-49)
    4.98621, 4.985024, 4.983895, 4.982825, 4.981821, 4.980885, 4.980024, 
    4.979245, 4.978554, 4.977959, 4.97747, 4.977098, 4.97686, 4.97678, 
    4.976899, 4.977179, 4.970335, 4.971414, 4.972563, 4.973532, 4.974247, 
    4.973269, 4.972249, 4.970926, 4.969913, 4.969187, 4.968878, 4.968968, 
    4.969584, 4.97014, 4.970872, 4.970227, 4.969762, 4.969515, 4.969513, 
    4.969784, 4.970358, 4.971261, 4.972516, 4.974138, 4.976139, 4.978522, 
    4.98128, 4.984394, 4.98783, 4.991536, 4.99544, 4.999442, 5.00342, 5.007222,
  // totalHeight(29,33, 0-49)
    4.986322, 4.985071, 4.98388, 4.982752, 4.981695, 4.980709, 4.979803, 
    4.978983, 4.978255, 4.977623, 4.977099, 4.976686, 4.976392, 4.976228, 
    4.976206, 4.976455, 4.97019, 4.970946, 4.971748, 4.972381, 4.972796, 
    4.971999, 4.971097, 4.969897, 4.968946, 4.968251, 4.967942, 4.968001, 
    4.96851, 4.968925, 4.969399, 4.968927, 4.968636, 4.968554, 4.968711, 
    4.969135, 4.969853, 4.970891, 4.972271, 4.97401, 4.976117, 4.978599, 
    4.981448, 4.984647, 4.988163, 4.991945, 4.995917, 4.999985, 5.00402, 
    5.007871,
  // totalHeight(29,34, 0-49)
    4.986467, 4.98515, 4.983893, 4.982704, 4.981585, 4.980543, 4.979585, 
    4.978714, 4.977937, 4.977258, 4.976682, 4.976209, 4.97584, 4.975573, 
    4.9754, 4.975558, 4.97007, 4.970491, 4.970932, 4.971223, 4.971337, 
    4.970714, 4.969939, 4.968884, 4.968016, 4.967366, 4.967063, 4.967083, 
    4.967473, 4.967741, 4.967969, 4.967685, 4.967576, 4.96767, 4.967996, 
    4.96858, 4.969448, 4.970625, 4.972131, 4.973985, 4.976196, 4.978769, 
    4.981701, 4.984973, 4.988553, 4.992392, 4.996415, 5.000526, 5.0046, 
    5.008479,
  // totalHeight(29,35, 0-49)
    4.986632, 4.985251, 4.98393, 4.982677, 4.981496, 4.980392, 4.979373, 
    4.978443, 4.977607, 4.976867, 4.976226, 4.97568, 4.975222, 4.97484, 
    4.974514, 4.974512, 4.969934, 4.970024, 4.970108, 4.97006, 4.969883, 
    4.969428, 4.968791, 4.967904, 4.967138, 4.966548, 4.966253, 4.966227, 
    4.96648, 4.966601, 4.966601, 4.96651, 4.966591, 4.96687, 4.967371, 
    4.968122, 4.969146, 4.970466, 4.972102, 4.974071, 4.976381, 4.979041, 
    4.982045, 4.985377, 4.989005, 4.99288, 4.996932, 5.001062, 5.005144, 
    5.009022,
  // totalHeight(29,36, 0-49)
    4.986797, 4.985363, 4.983984, 4.98267, 4.981424, 4.980255, 4.97917, 
    4.978174, 4.977268, 4.976458, 4.97574, 4.97511, 4.974553, 4.974052, 
    4.973577, 4.973351, 4.969756, 4.969531, 4.96927, 4.968902, 4.968448, 
    4.968158, 4.967667, 4.966969, 4.966328, 4.965811, 4.965522, 4.965443, 
    4.965545, 4.965516, 4.965311, 4.965418, 4.965693, 4.96616, 4.966842, 
    4.967765, 4.968948, 4.970416, 4.972183, 4.974266, 4.976675, 4.979414, 
    4.98248, 4.985857, 4.989515, 4.993406, 4.99746, 5.001577, 5.005634, 
    5.009474,
  // totalHeight(29,37, 0-49)
    4.986938, 4.985464, 4.984036, 4.982665, 4.981359, 4.980126, 4.978973, 
    4.977904, 4.976924, 4.976033, 4.97523, 4.974505, 4.973844, 4.973222, 
    4.972605, 4.972109, 4.969525, 4.969004, 4.968421, 4.967756, 4.967048, 
    4.966916, 4.966578, 4.966092, 4.965594, 4.965162, 4.964882, 4.964739, 
    4.964676, 4.9645, 4.964114, 4.96442, 4.964892, 4.965548, 4.966413, 
    4.96751, 4.968857, 4.970472, 4.972372, 4.974567, 4.97707, 4.979882, 
    4.983001, 4.986409, 4.990077, 4.993959, 4.997983, 5.002053, 5.006046, 
    5.009804,
  // totalHeight(29,38, 0-49)
    4.987028, 4.985529, 4.984065, 4.982647, 4.981288, 4.979993, 4.978771, 
    4.977629, 4.976569, 4.975593, 4.974696, 4.973871, 4.973101, 4.972361, 
    4.971611, 4.970821, 4.969233, 4.968444, 4.967564, 4.96663, 4.965697, 
    4.965714, 4.965539, 4.96528, 4.964942, 4.964607, 4.964337, 4.964119, 
    4.963884, 4.963566, 4.96303, 4.963531, 4.964195, 4.965038, 4.966087, 
    4.967357, 4.968866, 4.970628, 4.972659, 4.974966, 4.977559, 4.980438, 
    4.983595, 4.98702, 4.990678, 4.994521, 4.998483, 5.002466, 5.006349, 
    5.009973,
  // totalHeight(29,39, 0-49)
    4.98703, 4.985528, 4.984045, 4.982595, 4.981189, 4.97984, 4.978554, 
    4.977337, 4.976196, 4.975132, 4.974139, 4.97321, 4.972332, 4.971474, 
    4.970599, 4.969515, 4.96888, 4.967854, 4.966705, 4.965531, 4.964404, 
    4.964564, 4.964558, 4.964538, 4.964377, 4.964149, 4.963889, 4.963593, 
    4.96318, 4.96273, 4.962073, 4.962762, 4.963613, 4.964639, 4.965863, 
    4.967302, 4.96897, 4.970879, 4.973037, 4.975451, 4.978129, 4.981064, 
    4.984251, 4.987672, 4.991296, 4.995074, 4.998935, 5.002787, 5.006506, 
    5.009941,
  // totalHeight(29,40, 0-49)
    4.986917, 4.985433, 4.98395, 4.982483, 4.981046, 4.979649, 4.978304, 
    4.977018, 4.975799, 4.974646, 4.973557, 4.972527, 4.971539, 4.970568, 
    4.969579, 4.968217, 4.968469, 4.967233, 4.965849, 4.964469, 4.963177, 
    4.963475, 4.963636, 4.963868, 4.963894, 4.963784, 4.963535, 4.963162, 
    4.962571, 4.962003, 4.961255, 4.962122, 4.963151, 4.964351, 4.965744, 
    4.967346, 4.969165, 4.971212, 4.973492, 4.976008, 4.978761, 4.981743, 
    4.984945, 4.988344, 4.991908, 4.995585, 4.999307, 5.002978, 5.006479, 
    5.00966,
  // totalHeight(29,41, 0-49)
    4.986656, 4.985214, 4.983752, 4.982286, 4.980833, 4.979402, 4.978008, 
    4.976662, 4.975368, 4.97413, 4.97295, 4.971819, 4.970726, 4.969647, 
    4.968551, 4.96694, 4.968, 4.966581, 4.964995, 4.963443, 4.96202, 
    4.962448, 4.962779, 4.963267, 4.963491, 4.963505, 4.963273, 4.962823, 
    4.962065, 4.961395, 4.960584, 4.96162, 4.962814, 4.964176, 4.965727, 
    4.967481, 4.969442, 4.971618, 4.974011, 4.976619, 4.979436, 4.98245, 
    4.98565, 4.989006, 4.992481, 4.996022, 4.99956, 5.002998, 5.00622, 5.00908,
  // totalHeight(29,42, 0-49)
    4.986219, 4.984845, 4.983426, 4.981982, 4.980528, 4.979081, 4.977652, 
    4.976253, 4.974894, 4.973581, 4.972313, 4.971088, 4.969896, 4.968716, 
    4.96752, 4.965698, 4.967477, 4.965904, 4.964147, 4.962456, 4.960933, 
    4.961483, 4.961984, 4.962727, 4.963152, 4.963299, 4.96309, 4.962575, 
    4.961663, 4.96091, 4.960064, 4.961257, 4.962603, 4.964114, 4.96581, 
    4.967701, 4.969793, 4.972085, 4.974578, 4.977262, 4.980129, 4.98316, 
    4.986334, 4.989621, 4.992977, 4.996344, 4.99965, 5.0028, 5.00568, 5.00815,
  // totalHeight(29,43, 0-49)
    4.985586, 4.984303, 4.982952, 4.981551, 4.980116, 4.978669, 4.977219, 
    4.975782, 4.97437, 4.97299, 4.971644, 4.970334, 4.969049, 4.967778, 
    4.966492, 4.964496, 4.966899, 4.965197, 4.963301, 4.961505, 4.959913, 
    4.960582, 4.961247, 4.96224, 4.962868, 4.963152, 4.962977, 4.962408, 
    4.961366, 4.960551, 4.959695, 4.961031, 4.962516, 4.964162, 4.965988, 
    4.968001, 4.970206, 4.972599, 4.975173, 4.977917, 4.980814, 4.983839, 
    4.986966, 4.990153, 4.993352, 4.996504, 4.999529, 5.002333, 5.004804, 
    5.006812,
  // totalHeight(29,44, 0-49)
    4.984741, 4.983572, 4.98231, 4.980974, 4.979583, 4.978152, 4.9767, 
    4.975242, 4.973791, 4.972355, 4.970943, 4.969557, 4.968193, 4.966837, 
    4.96547, 4.96334, 4.966269, 4.964459, 4.962457, 4.960586, 4.958953, 
    4.959734, 4.960559, 4.961791, 4.962621, 4.963047, 4.962915, 4.962311, 
    4.961167, 4.960318, 4.959472, 4.96094, 4.96255, 4.964314, 4.966252, 
    4.968369, 4.970668, 4.973141, 4.975777, 4.978558, 4.981461, 4.984454, 
    4.987502, 4.990557, 4.993561, 4.996449, 4.999139, 5.001537, 5.003535, 
    5.00501,
  // totalHeight(29,45, 0-49)
    4.983676, 4.982643, 4.981495, 4.980247, 4.978919, 4.977528, 4.976092, 
    4.974628, 4.973153, 4.971678, 4.970212, 4.968764, 4.967327, 4.965899, 
    4.964459, 4.962228, 4.965582, 4.963693, 4.96161, 4.959693, 4.958048, 
    4.958934, 4.95991, 4.961367, 4.962389, 4.962958, 4.962886, 4.962271, 
    4.961058, 4.960199, 4.959386, 4.960973, 4.962695, 4.964563, 4.966595, 
    4.968796, 4.971167, 4.973697, 4.976369, 4.979159, 4.982038, 4.984967, 
    4.987901, 4.990783, 4.99355, 4.996124, 4.998423, 5.000354, 5.001812, 
    5.002688,
  // totalHeight(29,46, 0-49)
    4.982392, 4.981516, 4.980502, 4.979363, 4.978121, 4.976789, 4.97539, 
    4.973942, 4.972459, 4.970959, 4.969454, 4.967954, 4.96646, 4.964968, 
    4.963467, 4.961162, 4.96484, 4.962892, 4.96076, 4.958823, 4.957186, 
    4.958171, 4.959288, 4.960949, 4.962153, 4.962865, 4.962866, 4.962266, 
    4.961024, 4.960183, 4.959423, 4.961119, 4.962938, 4.964893, 4.967002, 
    4.969267, 4.971686, 4.974245, 4.976924, 4.979692, 4.982513, 4.985339, 
    4.988117, 4.990781, 4.993258, 4.995465, 4.997318, 4.998721, 4.999578, 
    4.999793,
  // totalHeight(29,47, 0-49)
    4.980901, 4.9802, 4.979339, 4.97833, 4.977193, 4.975943, 4.9746, 
    4.973184, 4.971713, 4.970206, 4.968677, 4.967138, 4.965598, 4.964054, 
    4.962501, 4.960147, 4.964045, 4.96206, 4.959902, 4.957967, 4.956358, 
    4.957434, 4.958677, 4.960518, 4.961888, 4.96274, 4.962831, 4.962277, 
    4.961047, 4.960255, 4.959564, 4.961359, 4.963265, 4.965293, 4.967459, 
    4.969764, 4.972204, 4.974763, 4.977415, 4.980123, 4.982846, 4.985526, 
    4.988099, 4.990493, 4.992628, 4.994412, 4.995758, 4.996574, 4.996771, 
    4.996272,
  // totalHeight(29,48, 0-49)
    4.979223, 4.978709, 4.978018, 4.977159, 4.976146, 4.974998, 4.973732, 
    4.972368, 4.970926, 4.969428, 4.967888, 4.966326, 4.96475, 4.963166, 
    4.961571, 4.959184, 4.963201, 4.961198, 4.959035, 4.957121, 4.955557, 
    4.956709, 4.958065, 4.960053, 4.961572, 4.96256, 4.962756, 4.96228, 
    4.961107, 4.960392, 4.959789, 4.961674, 4.963654, 4.965738, 4.967942, 
    4.970265, 4.972701, 4.975228, 4.977816, 4.980423, 4.983, 4.985481, 
    4.987796, 4.989864, 4.991597, 4.992898, 4.993679, 4.993851, 4.993337, 
    4.992082,
  // totalHeight(29,49, 0-49)
    4.977364, 4.976999, 4.976442, 4.975697, 4.974771, 4.973678, 4.972433, 
    4.97105, 4.96955, 4.967954, 4.966277, 4.964537, 4.96275, 4.960918, 
    4.959042, 4.955583, 4.965085, 4.962095, 4.958641, 4.955575, 4.95313, 
    4.956073, 4.959288, 4.963607, 4.966753, 4.968592, 4.96859, 4.966987, 
    4.963706, 4.96112, 4.958558, 4.960826, 4.963123, 4.965455, 4.967843, 
    4.970289, 4.972789, 4.975318, 4.977843, 4.980316, 4.982681, 4.984867, 
    4.986794, 4.988374, 4.989514, 4.990113, 4.990091, 4.989372, 4.987904, 
    4.98567 ;

 bathymetry =
  // bathymetry(0, 0-49)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  // bathymetry(1, 0-49)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  // bathymetry(2, 0-49)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  // bathymetry(3, 0-49)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  // bathymetry(4, 0-49)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  // bathymetry(5, 0-49)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  // bathymetry(6, 0-49)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  // bathymetry(7, 0-49)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  // bathymetry(8, 0-49)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  // bathymetry(9, 0-49)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  // bathymetry(10, 0-49)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  // bathymetry(11, 0-49)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  // bathymetry(12, 0-49)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  // bathymetry(13, 0-49)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  // bathymetry(14, 0-49)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  // bathymetry(15, 0-49)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  // bathymetry(16, 0-49)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  // bathymetry(17, 0-49)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  // bathymetry(18, 0-49)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  // bathymetry(19, 0-49)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  // bathymetry(20, 0-49)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  // bathymetry(21, 0-49)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  // bathymetry(22, 0-49)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  // bathymetry(23, 0-49)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  // bathymetry(24, 0-49)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  // bathymetry(25, 0-49)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  // bathymetry(26, 0-49)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  // bathymetry(27, 0-49)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  // bathymetry(28, 0-49)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  // bathymetry(29, 0-49)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  // bathymetry(30, 0-49)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  // bathymetry(31, 0-49)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  // bathymetry(32, 0-49)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  // bathymetry(33, 0-49)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  // bathymetry(34, 0-49)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  // bathymetry(35, 0-49)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  // bathymetry(36, 0-49)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  // bathymetry(37, 0-49)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  // bathymetry(38, 0-49)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  // bathymetry(39, 0-49)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  // bathymetry(40, 0-49)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  // bathymetry(41, 0-49)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  // bathymetry(42, 0-49)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  // bathymetry(43, 0-49)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  // bathymetry(44, 0-49)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  // bathymetry(45, 0-49)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  // bathymetry(46, 0-49)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  // bathymetry(47, 0-49)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  // bathymetry(48, 0-49)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  // bathymetry(49, 0-49)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0 ;

 momentumX =
  // momentumX(0,0, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumX(0,1, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumX(0,2, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumX(0,3, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumX(0,4, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumX(0,5, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumX(0,6, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumX(0,7, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumX(0,8, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumX(0,9, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumX(0,10, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumX(0,11, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumX(0,12, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumX(0,13, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumX(0,14, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumX(0,15, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumX(0,16, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumX(0,17, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumX(0,18, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumX(0,19, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumX(0,20, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 0, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumX(0,21, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 0, 5, 5, 5, 5, 5, 5, 5, 10, 
    10, 10, 10, 10, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5,
  // momentumX(0,22, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 0, 5, 5, 5, 5, 5, 5, 10, 10, 
    10, 10, 10, 10, 10, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5,
  // momentumX(0,23, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 0, 5, 5, 5, 5, 5, 10, 10, 
    10, 10, 10, 10, 10, 10, 10, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5,
  // momentumX(0,24, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 0, 5, 5, 5, 5, 5, 10, 10, 
    10, 10, 10, 10, 10, 10, 10, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5,
  // momentumX(0,25, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 0, 5, 5, 5, 5, 5, 10, 10, 
    10, 10, 10, 10, 10, 10, 10, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5,
  // momentumX(0,26, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 0, 5, 5, 5, 5, 5, 10, 10, 
    10, 10, 10, 10, 10, 10, 10, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5,
  // momentumX(0,27, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 0, 5, 5, 5, 5, 5, 10, 10, 
    10, 10, 10, 10, 10, 10, 10, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5,
  // momentumX(0,28, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 0, 5, 5, 5, 5, 5, 5, 10, 10, 
    10, 10, 10, 10, 10, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5,
  // momentumX(0,29, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 0, 5, 5, 5, 5, 5, 5, 5, 10, 
    10, 10, 10, 10, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5,
  // momentumX(0,30, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumX(0,31, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumX(0,32, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumX(0,33, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumX(0,34, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumX(0,35, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumX(0,36, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumX(0,37, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumX(0,38, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumX(0,39, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumX(0,40, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumX(0,41, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumX(0,42, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumX(0,43, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumX(0,44, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumX(0,45, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumX(0,46, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumX(0,47, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumX(0,48, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumX(0,49, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumX(1,0, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumX(1,1, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumX(1,2, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumX(1,3, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumX(1,4, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumX(1,5, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumX(1,6, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumX(1,7, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumX(1,8, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumX(1,9, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5.000001, 5.000003, 5.000003, 5.000003, 5.000003, 5.000003, 5.000001, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumX(1,10, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 
    5.00001, 5.000023, 5.000029, 5.00003, 5.000029, 5.000023, 5.00001, 
    5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumX(1,11, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000005, 
    5.000022, 5.000071, 5.000165, 5.000208, 5.000218, 5.000208, 5.000165, 
    5.000071, 5.000022, 5.000005, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5,
  // momentumX(1,12, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000009, 
    5.000041, 5.000161, 5.000472, 5.00103, 5.001293, 5.001361, 5.001293, 
    5.00103, 5.000472, 5.000161, 5.000041, 5.000009, 5.000001, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumX(1,13, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000013, 
    5.000065, 5.00028, 5.000989, 5.002667, 5.005479, 5.00688, 5.007271, 
    5.00688, 5.005479, 5.002667, 5.000989, 5.00028, 5.000065, 5.000013, 
    5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumX(1,14, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000016, 
    5.000087, 5.000412, 5.001609, 5.005196, 5.012874, 5.024823, 5.031068, 
    5.032917, 5.031068, 5.024823, 5.012874, 5.005196, 5.001609, 5.000412, 
    5.000087, 5.000016, 5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumX(1,15, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000018, 
    5.000104, 5.000527, 5.002232, 5.007843, 5.023126, 5.05233, 5.093832, 
    5.116333, 5.123362, 5.116333, 5.093832, 5.05233, 5.023126, 5.007843, 
    5.002232, 5.000527, 5.000104, 5.000018, 5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5,
  // momentumX(1,16, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000016, 5.000111, 
    5.000595, 5.002696, 5.010195, 5.032046, 5.08562, 5.174296, 5.284347, 
    5.345138, 5.365025, 5.345138, 5.284347, 5.174296, 5.08562, 5.032046, 
    5.010195, 5.002696, 5.000595, 5.00011, 5.000018, 5.000002, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5,
  // momentumX(1,17, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000013, 5.000091, 
    5.000609, 5.00287, 5.011568, 5.038834, 5.107607, 5.255316, 5.45458, 
    5.654781, 5.766831, 5.805127, 5.766831, 5.654781, 5.45458, 5.255316, 
    5.107607, 5.038834, 5.011568, 5.002866, 5.000595, 5.000104, 5.000016, 
    5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumX(1,18, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000008, 5.00006, 5.000425, 
    5.002811, 5.011596, 5.041329, 5.121252, 5.288161, 5.587032, 5.889495, 
    6.114048, 6.247925, 6.296353, 6.247925, 6.114048, 5.889495, 5.587032, 
    5.288161, 5.121252, 5.041325, 5.011568, 5.002696, 5.000527, 5.000087, 
    5.000013, 5.000001, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumX(1,19, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000003, 5.000028, 5.000218, 
    5.001533, 5.011003, 5.039038, 5.121291, 5.303221, 5.596775, 6.011393, 
    6.30257, 6.444544, 6.550306, 6.591668, 6.550305, 6.444544, 6.30257, 
    6.011393, 5.596775, 5.303215, 5.121252, 5.038834, 5.010195, 5.002232, 
    5.000412, 5.000065, 5.000009, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumX(1,20, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000014, 0, 5.039814, 
    5.109214, 5.288445, 5.596817, 5.95014, 6.326973, 6.498679, 6.541141, 
    6.600243, 6.624728, 6.600243, 6.541141, 6.498679, 6.326972, 5.950134, 
    5.596775, 5.288161, 5.107607, 5.032046, 5.007843, 5.001609, 5.00028, 
    5.000041, 5.000005, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumX(1,21, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 0, 5.108829, 
    5.260567, 5.588036, 6.011554, 6.326994, 6.546953, 6.566364, 6.535832, 
    6.558554, 6.576564, 6.558554, 6.535832, 6.566363, 6.546951, 6.326972, 
    6.011393, 5.587032, 5.255316, 5.08562, 5.023126, 5.005196, 5.000989, 
    5.000161, 5.000022, 5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumX(1,22, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 0, 5.226802, 5.467532, 
    5.892158, 6.303021, 6.498741, 6.56637, 6.621973, 6.765517, 6.920608, 
    6.987292, 6.920608, 6.765517, 6.621973, 6.566362, 6.498679, 6.30257, 
    5.889495, 5.45458, 5.174296, 5.05233, 5.012874, 5.002667, 5.000472, 
    5.000071, 5.00001, 5.000001, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumX(1,23, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 0, 5.378377, 5.679589, 
    6.119381, 6.445471, 6.541272, 6.535846, 6.765518, 7.138705, 7.442398, 
    7.559381, 7.442398, 7.138703, 6.765517, 6.535831, 6.541141, 6.444544, 
    6.114048, 5.654781, 5.284347, 5.093832, 5.024823, 5.005479, 5.00103, 
    5.000165, 5.000023, 5.000003, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumX(1,24, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 0, 5.461733, 5.797845, 
    6.254579, 6.551452, 6.600401, 6.558572, 6.920609, 7.442399, 7.841739, 
    7.990802, 7.841739, 7.442398, 6.920608, 6.558555, 6.600243, 6.550306, 
    6.247925, 5.766831, 5.345138, 5.116333, 5.031068, 5.00688, 5.001293, 
    5.000208, 5.000029, 5.000003, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumX(1,25, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 0, 5.488677, 5.83798, 
    6.303374, 6.592873, 6.624895, 6.576583, 6.987293, 7.559382, 7.990802, 
    8.150589, 7.990803, 7.559381, 6.987291, 6.576564, 6.624729, 6.591668, 
    6.296353, 5.805127, 5.365025, 5.123362, 5.032917, 5.007271, 5.001361, 
    5.000218, 5.00003, 5.000003, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumX(1,26, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 0, 5.461732, 5.797844, 
    6.254579, 6.551452, 6.600401, 6.558572, 6.920609, 7.442398, 7.841739, 
    7.990802, 7.841739, 7.442398, 6.920608, 6.558555, 6.600243, 6.550306, 
    6.247925, 5.766831, 5.345138, 5.116333, 5.031068, 5.00688, 5.001293, 
    5.000208, 5.000029, 5.000003, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumX(1,27, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 0, 5.378368, 
    5.679588, 6.119381, 6.445471, 6.541272, 6.535846, 6.765518, 7.138705, 
    7.442398, 7.55938, 7.442398, 7.138704, 6.765517, 6.535832, 6.541142, 
    6.444544, 6.114048, 5.654781, 5.284347, 5.093832, 5.024823, 5.005479, 
    5.00103, 5.000165, 5.000023, 5.000003, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumX(1,28, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000009, 0, 5.226734, 
    5.467518, 5.892155, 6.303021, 6.498741, 6.56637, 6.621974, 6.765516, 
    6.920608, 6.987291, 6.920608, 6.765516, 6.621973, 6.566363, 6.498679, 
    6.30257, 5.889495, 5.45458, 5.174296, 5.05233, 5.012874, 5.002667, 
    5.000472, 5.000071, 5.00001, 5.000001, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumX(1,29, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000013, 5.00007, 0, 
    5.108382, 5.260472, 5.588021, 6.011552, 6.326994, 6.546954, 6.566364, 
    6.535832, 6.558555, 6.576563, 6.558555, 6.535832, 6.566363, 6.546951, 
    6.326972, 6.011393, 5.587032, 5.255316, 5.08562, 5.023126, 5.005196, 
    5.000989, 5.000161, 5.000022, 5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumX(1,30, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000017, 5.000138, 5.000946, 
    5.005786, 5.03459, 5.108321, 5.288314, 5.5968, 5.950139, 6.326973, 
    6.49868, 6.541142, 6.600243, 6.624728, 6.600243, 6.541142, 6.498679, 
    6.326972, 5.950134, 5.596775, 5.288161, 5.107607, 5.032046, 5.007843, 
    5.001609, 5.00028, 5.000041, 5.000005, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumX(1,31, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000005, 5.000042, 5.000306, 
    5.001886, 5.010614, 5.038951, 5.121276, 5.303219, 5.596775, 6.011393, 
    6.30257, 6.444544, 6.550306, 6.591668, 6.550306, 6.444544, 6.30257, 
    6.011393, 5.596775, 5.303215, 5.121252, 5.038834, 5.010195, 5.002232, 
    5.000412, 5.000065, 5.000009, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumX(1,32, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000009, 5.000072, 5.000477, 
    5.002755, 5.011584, 5.041328, 5.121252, 5.288161, 5.587032, 5.889495, 
    6.114048, 6.247925, 6.296353, 6.247925, 6.114048, 5.889495, 5.587032, 
    5.288161, 5.121252, 5.041325, 5.011568, 5.002696, 5.000527, 5.000087, 
    5.000013, 5.000001, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumX(1,33, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000014, 5.000097, 
    5.000602, 5.002868, 5.011568, 5.038834, 5.107607, 5.255316, 5.45458, 
    5.654781, 5.766831, 5.805127, 5.766831, 5.654781, 5.45458, 5.255316, 
    5.107607, 5.038834, 5.011568, 5.002866, 5.000595, 5.000104, 5.000016, 
    5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumX(1,34, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000017, 5.00011, 
    5.000595, 5.002696, 5.010195, 5.032046, 5.08562, 5.174296, 5.284347, 
    5.345138, 5.365025, 5.345138, 5.284347, 5.174296, 5.08562, 5.032046, 
    5.010195, 5.002696, 5.000595, 5.00011, 5.000018, 5.000002, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5,
  // momentumX(1,35, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000018, 
    5.000104, 5.000527, 5.002232, 5.007843, 5.023126, 5.05233, 5.093832, 
    5.116333, 5.123362, 5.116333, 5.093832, 5.05233, 5.023126, 5.007843, 
    5.002232, 5.000527, 5.000104, 5.000018, 5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5,
  // momentumX(1,36, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000016, 
    5.000087, 5.000412, 5.001609, 5.005196, 5.012874, 5.024823, 5.031068, 
    5.032917, 5.031068, 5.024823, 5.012874, 5.005196, 5.001609, 5.000412, 
    5.000087, 5.000016, 5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumX(1,37, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000013, 
    5.000065, 5.00028, 5.000989, 5.002667, 5.005479, 5.00688, 5.007271, 
    5.00688, 5.005479, 5.002667, 5.000989, 5.00028, 5.000065, 5.000013, 
    5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumX(1,38, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000009, 
    5.000041, 5.000161, 5.000472, 5.00103, 5.001293, 5.001361, 5.001293, 
    5.00103, 5.000472, 5.000161, 5.000041, 5.000009, 5.000001, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumX(1,39, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000005, 
    5.000022, 5.000071, 5.000165, 5.000208, 5.000218, 5.000208, 5.000165, 
    5.000071, 5.000022, 5.000005, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5,
  // momentumX(1,40, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 
    5.00001, 5.000023, 5.000029, 5.00003, 5.000029, 5.000023, 5.00001, 
    5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumX(1,41, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5.000001, 5.000003, 5.000003, 5.000003, 5.000003, 5.000003, 5.000001, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumX(1,42, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumX(1,43, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumX(1,44, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumX(1,45, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumX(1,46, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumX(1,47, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumX(1,48, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumX(1,49, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumX(2,0, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumX(2,1, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumX(2,2, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumX(2,3, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5.000001, 5.000001, 5.000001, 5.000001, 5.000001, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumX(2,4, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 
    5.000003, 5.000006, 5.000008, 5.000009, 5.000008, 5.000006, 5.000003, 
    5.000001, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumX(2,5, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 
    5.000003, 5.000009, 5.000018, 5.00003, 5.000037, 5.000041, 5.000037, 
    5.00003, 5.000018, 5.000009, 5.000003, 5.000001, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumX(2,6, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000008, 
    5.00002, 5.000044, 5.000084, 5.000135, 5.000167, 5.000179, 5.000167, 
    5.000135, 5.000084, 5.000044, 5.00002, 5.000008, 5.000002, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumX(2,7, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000004, 5.000013, 
    5.000036, 5.000087, 5.000192, 5.000359, 5.000562, 5.000698, 5.000745, 
    5.000698, 5.000562, 5.000359, 5.000192, 5.000087, 5.000036, 5.000013, 
    5.000004, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumX(2,8, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000005, 
    5.000019, 5.000055, 5.000149, 5.000361, 5.000768, 5.001396, 5.002146, 
    5.002654, 5.002829, 5.002654, 5.002146, 5.001396, 5.000768, 5.000361, 
    5.000149, 5.000055, 5.000019, 5.000005, 5.000001, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5,
  // momentumX(2,9, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000007, 5.000025, 
    5.00008, 5.00023, 5.000596, 5.001375, 5.002819, 5.004971, 5.00749, 
    5.009201, 5.009799, 5.009201, 5.00749, 5.004971, 5.002819, 5.001375, 
    5.000596, 5.00023, 5.00008, 5.000025, 5.000007, 5.000001, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5,
  // momentumX(2,10, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000008, 5.000031, 
    5.000104, 5.000319, 5.000876, 5.002162, 5.004771, 5.009418, 5.016093, 
    5.023739, 5.028931, 5.030761, 5.028931, 5.023739, 5.016093, 5.009418, 
    5.004771, 5.002162, 5.000876, 5.000319, 5.000104, 5.000031, 5.000008, 
    5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumX(2,11, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.00001, 5.000034, 
    5.000126, 5.000408, 5.001172, 5.003046, 5.007127, 5.014987, 5.028435, 
    5.046975, 5.067611, 5.08152, 5.086449, 5.08152, 5.067611, 5.046975, 
    5.028435, 5.014987, 5.007127, 5.003045, 5.001171, 5.000405, 5.000127, 
    5.000036, 5.00001, 5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumX(2,12, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000009, 5.000036, 5.000136, 
    5.000466, 5.001442, 5.003905, 5.00958, 5.021203, 5.042273, 5.076715, 
    5.121716, 5.169673, 5.201324, 5.212531, 5.201324, 5.169673, 5.121716, 
    5.076715, 5.042273, 5.021201, 5.009576, 5.003897, 5.00143, 5.000474, 
    5.000143, 5.000039, 5.00001, 5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumX(2,13, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000008, 5.000033, 5.000133, 
    5.000481, 5.00157, 5.004634, 5.011772, 5.027131, 5.05641, 5.105655, 
    5.181499, 5.273223, 5.364344, 5.422204, 5.4425, 5.422204, 5.364344, 
    5.273223, 5.181498, 5.105653, 5.056403, 5.02711, 5.011728, 5.004572, 
    5.001609, 5.000513, 5.000149, 5.000039, 5.00001, 5.000002, 5, 5, 5, 5, 5, 
    5, 5, 5, 5,
  // momentumX(2,14, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000007, 5.000029, 5.000118, 5.000446, 
    5.001536, 5.004781, 5.013485, 5.031936, 5.068588, 5.132482, 5.229629, 
    5.367397, 5.516597, 5.650199, 5.73082, 5.75868, 5.73082, 5.650199, 
    5.516597, 5.367393, 5.229616, 5.132443, 5.068489, 5.031737, 5.013205, 
    5.004946, 5.001672, 5.000513, 5.000143, 5.000036, 5.000008, 5.000001, 5, 
    5, 5, 5, 5, 5, 5, 5,
  // momentumX(2,15, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000004, 5.000021, 5.000093, 5.000368, 
    5.001338, 5.004398, 5.013077, 5.035445, 5.07743, 5.152986, 5.270136, 
    5.425341, 5.623005, 5.808567, 5.954159, 6.038265, 6.066943, 6.038265, 
    5.954158, 5.808562, 5.622989, 5.425284, 5.269968, 5.152572, 5.076609, 
    5.034278, 5.01373, 5.004946, 5.001609, 5.000474, 5.000127, 5.000031, 
    5.000007, 5.000001, 5, 5, 5, 5, 5, 5, 5,
  // momentumX(2,16, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000014, 5.000063, 5.000268, 5.001024, 
    5.003561, 5.011195, 5.031907, 5.083897, 5.166404, 5.297246, 5.471339, 
    5.663941, 5.881144, 6.054009, 6.170801, 6.238191, 6.261086, 6.23819, 
    6.170798, 6.053992, 5.881079, 5.663725, 5.470706, 5.295689, 5.163324, 
    5.079466, 5.034278, 5.013205, 5.004572, 5.00143, 5.000405, 5.000104, 
    5.000025, 5.000005, 5, 5, 5, 5, 5, 5, 5,
  // momentumX(2,17, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000008, 5.000038, 5.000165, 5.00067, 
    5.002472, 5.008275, 5.024992, 5.068762, 5.178341, 5.314689, 5.498798, 
    5.701071, 5.878989, 6.057094, 6.174425, 6.241654, 6.28508, 6.300066, 
    6.285078, 6.24164, 6.174369, 6.056881, 5.878283, 5.699006, 5.493689, 
    5.304491, 5.163324, 5.076609, 5.031737, 5.011728, 5.003897, 5.001171, 
    5.000319, 5.00008, 5.000019, 5.000004, 5, 5, 5, 5, 5, 5,
  // momentumX(2,18, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5.000003, 5.000017, 5.000082, 5.000356, 5.001401, 
    5.005028, 5.016359, 5.047846, 5.129076, 5.339933, 5.523062, 5.725195, 
    5.900149, 6.010222, 6.107472, 6.153584, 6.174073, 6.196599, 6.204854, 
    6.196589, 6.174033, 6.153419, 6.106858, 6.008182, 5.894237, 5.710595, 
    5.493689, 5.295689, 5.152572, 5.068489, 5.02711, 5.009576, 5.003045, 
    5.000876, 5.00023, 5.000055, 5.000013, 5.000002, 5, 5, 5, 5, 5,
  // momentumX(2,19, 0-49)
    5, 5, 5, 5, 5, 5, 5.000001, 5.000007, 5.000029, 5.000135, 5.000575, 
    5.002245, 5.008015, 5.025926, 5.074886, 5.206708, 5.580922, 5.772137, 
    5.930871, 6.024444, 6.039964, 6.04226, 6.020387, 6.004436, 6.009708, 
    6.012484, 6.009684, 6.004327, 6.019951, 6.040654, 6.034697, 6.009424, 
    5.894236, 5.699005, 5.470706, 5.269968, 5.132443, 5.056403, 5.021201, 
    5.007127, 5.002162, 5.000596, 5.000149, 5.000036, 5.000008, 5.000001, 5, 
    5, 5, 5,
  // momentumX(2,20, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5.000001, 5.00001, 5.000042, 5.000171, 5.000613, 
    5.001966, 5.005518, 5.013143, 0, 6.070654, 6.10031, 6.109229, 6.073961, 
    5.989838, 5.897338, 5.812802, 5.764136, 5.750331, 5.746961, 5.750273, 
    5.763871, 5.811723, 5.893331, 5.976495, 6.034697, 6.008182, 5.878282, 
    5.663725, 5.425284, 5.229616, 5.105653, 5.042273, 5.014987, 5.004771, 
    5.001375, 5.000361, 5.000087, 5.00002, 5.000003, 5, 5, 5, 5,
  // momentumX(2,21, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5.000003, 5.000014, 5.000054, 5.000195, 5.00063, 
    5.001772, 5.004181, 0, 6.513035, 6.426273, 6.282675, 6.110457, 5.917133, 
    5.702082, 5.514227, 5.387189, 5.318944, 5.296926, 5.318848, 5.386738, 
    5.51234, 5.694969, 5.893331, 6.040654, 6.106857, 6.056882, 5.88108, 
    5.622988, 5.367393, 5.181498, 5.076715, 5.028435, 5.009418, 5.002819, 
    5.000768, 5.000192, 5.000044, 5.000009, 5.000001, 5, 5, 5,
  // momentumX(2,22, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000004, 5.000016, 5.000055, 5.000182, 
    5.000515, 5.001205, 0, 6.890601, 6.696692, 6.413081, 6.125101, 5.847679, 
    5.523096, 5.231614, 5.02129, 4.898302, 4.858558, 4.898164, 5.020628, 
    5.228783, 5.512339, 5.811723, 6.019951, 6.153419, 6.174369, 6.053992, 
    5.808561, 5.516597, 5.273223, 5.121716, 5.046975, 5.016093, 5.004971, 
    5.001396, 5.000359, 5.000084, 5.000018, 5.000003, 5, 5, 5,
  // momentumX(2,23, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000004, 5.000016, 5.000049, 5.000141, 
    5.000327, 0, 7.175317, 6.901651, 6.513165, 6.143483, 5.81144, 5.400992, 
    5.024344, 4.753988, 4.602839, 4.55656, 4.602668, 4.753143, 5.020628, 
    5.386737, 5.76387, 6.004326, 6.174033, 6.241639, 6.170797, 5.954158, 
    5.650199, 5.364344, 5.169673, 5.067611, 5.023739, 5.00749, 5.002146, 
    5.000562, 5.000135, 5.00003, 5.000006, 5.000001, 5, 5,
  // momentumX(2,24, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000006, 5.00002, 5.000057, 5.000128, 
    0, 7.33971, 7.028852, 6.586917, 6.171556, 5.805634, 5.335411, 4.902411, 
    4.603594, 4.448595, 4.40392, 4.448415, 4.602663, 4.89816, 5.318843, 
    5.750269, 6.009683, 6.196589, 6.285078, 6.23819, 6.038265, 5.73082, 
    5.422204, 5.201324, 5.08152, 5.028931, 5.009201, 5.002654, 5.000698, 
    5.000167, 5.000037, 5.000008, 5.000001, 5, 5,
  // momentumX(2,25, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000003, 5.000013, 5.000041, 5.000108, 
    5.000237, 0, 7.394997, 7.072412, 6.612961, 6.182293, 5.805012, 5.31426, 
    4.862948, 4.55748, 4.40407, 4.360934, 4.403889, 4.556526, 4.858529, 
    5.296904, 5.746947, 6.012478, 6.204852, 6.300065, 6.261086, 6.066943, 
    5.75868, 5.4425, 5.212531, 5.086449, 5.030761, 5.009799, 5.002829, 
    5.000745, 5.000179, 5.000041, 5.000009, 5.000001, 5, 5,
  // momentumX(2,26, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000003, 5.000014, 5.000048, 5.000146, 
    5.00039, 5.000851, 0, 7.33743, 7.027562, 6.586339, 6.171353, 5.805575, 
    5.335398, 4.902407, 4.603593, 4.448595, 4.403919, 4.448415, 4.602663, 
    4.898159, 5.318843, 5.750269, 6.009683, 6.196589, 6.285078, 6.23819, 
    6.038265, 5.73082, 5.422204, 5.201324, 5.08152, 5.028931, 5.009201, 
    5.002654, 5.000698, 5.000167, 5.000037, 5.000008, 5.000001, 5, 5,
  // momentumX(2,27, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5.000003, 5.000013, 5.000049, 5.000171, 5.000519, 
    5.001362, 5.002976, 0, 7.16783, 6.897426, 6.511255, 6.142797, 5.811236, 
    5.40094, 5.024333, 4.753986, 4.602839, 4.55656, 4.602669, 4.753144, 
    5.020627, 5.386737, 5.76387, 6.004327, 6.174033, 6.24164, 6.170797, 
    5.954158, 5.650199, 5.364344, 5.169673, 5.067611, 5.023739, 5.00749, 
    5.002146, 5.000562, 5.000135, 5.00003, 5.000006, 5.000001, 5, 5,
  // momentumX(2,28, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5.000002, 5.00001, 5.000044, 5.000165, 5.000557, 
    5.001666, 5.004333, 5.009483, 0, 6.869401, 6.684888, 6.407736, 6.123141, 
    5.847076, 5.522937, 5.231577, 5.021283, 4.898301, 4.858558, 4.898164, 
    5.020629, 5.228784, 5.51234, 5.811723, 6.019951, 6.153419, 6.174369, 
    6.053992, 5.808561, 5.516597, 5.273223, 5.121716, 5.046975, 5.016093, 
    5.004971, 5.001396, 5.000359, 5.000084, 5.000018, 5.000003, 5, 5, 5,
  // momentumX(2,29, 0-49)
    5, 5, 5, 5, 5, 5, 5.000001, 5.000007, 5.000031, 5.00013, 5.000485, 
    5.001624, 5.004813, 5.012438, 5.027185, 0, 6.458423, 6.39655, 6.269349, 
    6.105521, 5.915573, 5.701647, 5.514119, 5.387164, 5.318938, 5.296925, 
    5.318848, 5.386738, 5.51234, 5.694969, 5.893331, 6.040654, 6.106858, 
    6.056882, 5.88108, 5.622988, 5.367393, 5.181498, 5.076715, 5.028435, 
    5.009418, 5.002819, 5.000768, 5.000192, 5.000044, 5.000009, 5.000001, 5, 
    5, 5,
  // momentumX(2,30, 0-49)
    5, 5, 5, 5, 5, 5, 5.000004, 5.000019, 5.000091, 5.000392, 5.001544, 
    5.005568, 5.018255, 5.053765, 5.13902, 5.339774, 5.824156, 5.992731, 
    6.068674, 6.060568, 5.985876, 5.89627, 5.812539, 5.764076, 5.750317, 
    5.746958, 5.750272, 5.763871, 5.811723, 5.893331, 5.976495, 6.034697, 
    6.008182, 5.878283, 5.663725, 5.425284, 5.229616, 5.105653, 5.042273, 
    5.014987, 5.004771, 5.001375, 5.000361, 5.000087, 5.00002, 5.000003, 5, 
    5, 5, 5,
  // momentumX(2,31, 0-49)
    5, 5, 5, 5, 5, 5, 5.000002, 5.000012, 5.000059, 5.000257, 5.001028, 
    5.003737, 5.01235, 5.036781, 5.097425, 5.235366, 5.544514, 5.750298, 
    5.92068, 6.020491, 6.03864, 6.041875, 6.020286, 6.00441, 6.009703, 
    6.012483, 6.009684, 6.004327, 6.019951, 6.040655, 6.034697, 6.009424, 
    5.894237, 5.699006, 5.470706, 5.269968, 5.132443, 5.056403, 5.021201, 
    5.007127, 5.002162, 5.000596, 5.000149, 5.000036, 5.000008, 5.000001, 5, 
    5, 5, 5,
  // momentumX(2,32, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5.000005, 5.000028, 5.000126, 5.000518, 5.00194, 
    5.006609, 5.020349, 5.056161, 5.140028, 5.324083, 5.513662, 5.720868, 
    5.898491, 6.009674, 6.107315, 6.153543, 6.174064, 6.196596, 6.204853, 
    6.196589, 6.174033, 6.153419, 6.106858, 6.008182, 5.894237, 5.710595, 
    5.493689, 5.295689, 5.152572, 5.068489, 5.02711, 5.009576, 5.003045, 
    5.000876, 5.00023, 5.000055, 5.000013, 5.000002, 5, 5, 5, 5, 5,
  // momentumX(2,33, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000011, 5.000051, 5.000216, 5.000844, 
    5.002991, 5.009605, 5.02779, 5.072512, 5.172647, 5.311225, 5.497193, 
    5.700458, 5.878788, 6.057036, 6.17441, 6.241651, 6.28508, 6.300066, 
    6.285078, 6.241639, 6.174369, 6.056882, 5.878283, 5.699006, 5.493689, 
    5.304491, 5.163324, 5.076609, 5.031737, 5.011728, 5.003897, 5.001171, 
    5.000319, 5.00008, 5.000019, 5.000004, 5, 5, 5, 5, 5, 5,
  // momentumX(2,34, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5.000003, 5.000018, 5.000078, 5.000318, 5.001177, 
    5.003963, 5.012051, 5.033063, 5.082146, 5.165304, 5.29673, 5.471141, 
    5.663877, 5.881125, 6.054005, 6.170801, 6.238191, 6.261086, 6.238191, 
    6.170798, 6.053992, 5.88108, 5.663725, 5.470706, 5.295689, 5.163324, 
    5.079466, 5.034278, 5.013205, 5.004572, 5.00143, 5.000405, 5.000104, 
    5.000025, 5.000005, 5, 5, 5, 5, 5, 5, 5,
  // momentumX(2,35, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000006, 5.000025, 5.000106, 5.000411, 
    5.001449, 5.004638, 5.0134, 5.034968, 5.077124, 5.152843, 5.270081, 
    5.425323, 5.623, 5.808566, 5.954159, 6.038265, 6.066944, 6.038265, 
    5.954159, 5.808562, 5.622989, 5.425284, 5.269968, 5.152572, 5.076609, 
    5.034278, 5.01373, 5.004946, 5.001609, 5.000474, 5.000127, 5.000031, 
    5.000007, 5.000001, 5, 5, 5, 5, 5, 5, 5,
  // momentumX(2,36, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000007, 5.000031, 5.000127, 
    5.000473, 5.001596, 5.004863, 5.013367, 5.031859, 5.068552, 5.132469, 
    5.229624, 5.367395, 5.516597, 5.650199, 5.73082, 5.75868, 5.73082, 
    5.650199, 5.516597, 5.367393, 5.229616, 5.132443, 5.068489, 5.031737, 
    5.013205, 5.004946, 5.001672, 5.000513, 5.000143, 5.000036, 5.000008, 
    5.000001, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumX(2,37, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000009, 5.000036, 5.000139, 
    5.000494, 5.001589, 5.004607, 5.011755, 5.027123, 5.056408, 5.105654, 
    5.181498, 5.273223, 5.364344, 5.422204, 5.4425, 5.422204, 5.364344, 
    5.273223, 5.181498, 5.105653, 5.056403, 5.02711, 5.011728, 5.004572, 
    5.001609, 5.000513, 5.000149, 5.000039, 5.00001, 5.000002, 5, 5, 5, 5, 5, 
    5, 5, 5, 5,
  // momentumX(2,38, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.00001, 5.000037, 5.000138, 
    5.00047, 5.001437, 5.003901, 5.009578, 5.021202, 5.042273, 5.076715, 
    5.121716, 5.169673, 5.201324, 5.212531, 5.201324, 5.169673, 5.121716, 
    5.076715, 5.042273, 5.021201, 5.009576, 5.003897, 5.00143, 5.000474, 
    5.000143, 5.000039, 5.00001, 5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumX(2,39, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.00001, 5.000034, 
    5.000126, 5.000407, 5.001172, 5.003045, 5.007127, 5.014987, 5.028435, 
    5.046975, 5.067611, 5.08152, 5.086449, 5.08152, 5.067611, 5.046975, 
    5.028435, 5.014987, 5.007127, 5.003045, 5.001171, 5.000405, 5.000127, 
    5.000036, 5.00001, 5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumX(2,40, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000008, 5.000031, 
    5.000104, 5.000319, 5.000876, 5.002162, 5.004771, 5.009418, 5.016093, 
    5.023739, 5.028931, 5.030761, 5.028931, 5.023739, 5.016093, 5.009418, 
    5.004771, 5.002162, 5.000876, 5.000319, 5.000104, 5.000031, 5.000008, 
    5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumX(2,41, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000007, 5.000025, 
    5.00008, 5.00023, 5.000596, 5.001375, 5.002819, 5.004971, 5.00749, 
    5.009201, 5.009799, 5.009201, 5.00749, 5.004971, 5.002819, 5.001375, 
    5.000596, 5.00023, 5.00008, 5.000025, 5.000007, 5.000001, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5,
  // momentumX(2,42, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000005, 
    5.000019, 5.000055, 5.000149, 5.000361, 5.000768, 5.001396, 5.002146, 
    5.002654, 5.002829, 5.002654, 5.002146, 5.001396, 5.000768, 5.000361, 
    5.000149, 5.000055, 5.000019, 5.000005, 5.000001, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5,
  // momentumX(2,43, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000004, 5.000013, 
    5.000036, 5.000087, 5.000192, 5.000359, 5.000562, 5.000698, 5.000745, 
    5.000698, 5.000562, 5.000359, 5.000192, 5.000087, 5.000036, 5.000013, 
    5.000004, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumX(2,44, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000008, 
    5.00002, 5.000044, 5.000084, 5.000135, 5.000167, 5.000179, 5.000167, 
    5.000135, 5.000084, 5.000044, 5.00002, 5.000008, 5.000002, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumX(2,45, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 
    5.000003, 5.000009, 5.000018, 5.00003, 5.000037, 5.000041, 5.000037, 
    5.00003, 5.000018, 5.000009, 5.000003, 5.000001, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumX(2,46, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 
    5.000003, 5.000006, 5.000008, 5.000009, 5.000008, 5.000006, 5.000003, 
    5.000001, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumX(2,47, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5.000001, 5.000001, 5.000001, 5.000001, 5.000001, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumX(2,48, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumX(2,49, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumX(3,0, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 
    5.000003, 5.000006, 5.00001, 5.000014, 5.000018, 5.000019, 5.000018, 
    5.000014, 5.00001, 5.000006, 5.000003, 5.000001, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumX(3,1, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000007, 
    5.000014, 5.000024, 5.000038, 5.000054, 5.000065, 5.000069, 5.000065, 
    5.000054, 5.000038, 5.000024, 5.000014, 5.000007, 5.000002, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumX(3,2, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000005, 
    5.000013, 5.000025, 5.000051, 5.000089, 5.000139, 5.000192, 5.00023, 
    5.000245, 5.00023, 5.000192, 5.000139, 5.000089, 5.000051, 5.000025, 
    5.000013, 5.000005, 5.000001, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumX(3,3, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000003, 5.000008, 5.00002, 
    5.000045, 5.000092, 5.000175, 5.000303, 5.000471, 5.000645, 5.000771, 
    5.000815, 5.000771, 5.000645, 5.000471, 5.000303, 5.000175, 5.000092, 
    5.000045, 5.00002, 5.000008, 5.000003, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5,
  // momentumX(3,4, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000004, 5.000012, 5.00003, 
    5.00007, 5.000153, 5.000309, 5.000576, 5.000975, 5.001488, 5.002019, 
    5.0024, 5.002537, 5.0024, 5.002019, 5.001488, 5.000975, 5.000576, 
    5.000309, 5.000153, 5.00007, 5.00003, 5.000012, 5.000004, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5,
  // momentumX(3,5, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000005, 5.000016, 
    5.000041, 5.000101, 5.000232, 5.000495, 5.000975, 5.001767, 5.002935, 
    5.004404, 5.005916, 5.006993, 5.007383, 5.006993, 5.005916, 5.004404, 
    5.002935, 5.001767, 5.000974, 5.000495, 5.000232, 5.000101, 5.000041, 
    5.000016, 5.000005, 5.000001, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumX(3,6, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000007, 5.00002, 5.000052, 
    5.000135, 5.000328, 5.000727, 5.001502, 5.002871, 5.005065, 5.008235, 
    5.012152, 5.016148, 5.018981, 5.020005, 5.018981, 5.016148, 5.012152, 
    5.008235, 5.005065, 5.00287, 5.001501, 5.000726, 5.000327, 5.000136, 
    5.000052, 5.00002, 5.000007, 5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumX(3,7, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000008, 5.000022, 5.000062, 
    5.000168, 5.000426, 5.000994, 5.002136, 5.004256, 5.007876, 5.013505, 
    5.021459, 5.0311, 5.040833, 5.047673, 5.050141, 5.047673, 5.040833, 
    5.0311, 5.021459, 5.013503, 5.007874, 5.004254, 5.00213, 5.000989, 
    5.000427, 5.000171, 5.000064, 5.000023, 5.000008, 5.000002, 5, 5, 5, 5, 
    5, 5, 5, 5, 5,
  // momentumX(3,8, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000008, 5.000023, 5.000071, 
    5.000197, 5.000516, 5.001256, 5.002826, 5.005837, 5.011214, 5.020035, 
    5.033278, 5.051542, 5.073155, 5.094623, 5.109491, 5.114835, 5.109491, 
    5.094623, 5.073154, 5.05154, 5.033274, 5.020027, 5.011199, 5.005819, 
    5.002808, 5.001259, 5.000525, 5.000204, 5.000074, 5.000025, 5.000008, 
    5.000002, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumX(3,9, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000008, 5.000024, 5.000072, 5.000215, 
    5.000583, 5.001472, 5.003447, 5.007477, 5.01482, 5.027332, 5.046957, 
    5.07516, 5.112832, 5.155911, 5.197577, 5.225729, 5.235758, 5.225728, 
    5.197576, 5.155908, 5.112823, 5.075142, 5.046923, 5.027278, 5.014745, 
    5.00741, 5.003462, 5.001504, 5.000608, 5.000228, 5.00008, 5.000026, 
    5.000009, 5.000002, 5, 5, 5, 5, 5, 5, 5,
  // momentumX(3,10, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000007, 5.000022, 5.000071, 5.000216, 
    5.00061, 5.001602, 5.003899, 5.008797, 5.018371, 5.034782, 5.061243, 
    5.100461, 5.15364, 5.221577, 5.295402, 5.36382, 5.408352, 5.423996, 
    5.408351, 5.363815, 5.29539, 5.221547, 5.153577, 5.100338, 5.061041, 
    5.034512, 5.018124, 5.008841, 5.004006, 5.001688, 5.000662, 5.000242, 
    5.000082, 5.000026, 5.000008, 5.000002, 5, 5, 5, 5, 5, 5,
  // momentumX(3,11, 0-49)
    5, 5, 5, 5, 5, 5, 5.000001, 5.000006, 5.000021, 5.000064, 5.000203, 
    5.000594, 5.001617, 5.004089, 5.009582, 5.020787, 5.04175, 5.075024, 
    5.125049, 5.193873, 5.280046, 5.383638, 5.488432, 5.579867, 5.636599, 
    5.656176, 5.636593, 5.57985, 5.488389, 5.383534, 5.279824, 5.193449, 
    5.124352, 5.074101, 5.040899, 5.020916, 5.009921, 5.004369, 5.001788, 
    5.000681, 5.000242, 5.00008, 5.000025, 5.000008, 5.000002, 5, 5, 5, 5, 5,
  // momentumX(3,12, 0-49)
    5, 5, 5, 5, 5, 5, 5.000005, 5.000017, 5.000055, 5.000177, 5.000535, 
    5.001513, 5.003968, 5.009657, 5.021753, 5.045288, 5.087358, 5.14761, 
    5.230261, 5.333305, 5.449304, 5.57871, 5.698251, 5.795069, 5.852182, 
    5.871558, 5.852166, 5.795019, 5.698119, 5.578391, 5.448622, 5.331985, 
    5.228084, 5.144711, 5.084641, 5.045663, 5.022761, 5.010503, 5.004496, 
    5.001788, 5.000662, 5.000228, 5.000074, 5.000023, 5.000007, 5.000001, 5, 
    5, 5, 5,
  // momentumX(3,13, 0-49)
    5, 5, 5, 5, 5, 5.000002, 5.000013, 5.000043, 5.000142, 5.000446, 
    5.001304, 5.003549, 5.008974, 5.021013, 5.045398, 5.090425, 5.167326, 
    5.262846, 5.378967, 5.506453, 5.631666, 5.760675, 5.867614, 5.947062, 
    5.992007, 6.007091, 5.991964, 5.946927, 5.867256, 5.75981, 5.629799, 
    5.502812, 5.372893, 5.25464, 5.159427, 5.091476, 5.048205, 5.023404, 
    5.010503, 5.004369, 5.001688, 5.000608, 5.000204, 5.000064, 5.00002, 
    5.000005, 5, 5, 5, 5,
  // momentumX(3,14, 0-49)
    5, 5, 5, 5, 5.000001, 5.000009, 5.000031, 5.000105, 5.00034, 5.001029, 
    5.002908, 5.007648, 5.018635, 5.041913, 5.086556, 5.164249, 5.291772, 
    5.421392, 5.55587, 5.681244, 5.783919, 5.882294, 5.952684, 5.99908, 
    6.024866, 6.03354, 6.024758, 5.998743, 5.951796, 5.880162, 5.77933, 
    5.672307, 5.540854, 5.400769, 5.271254, 5.167127, 5.093842, 5.048205, 
    5.022761, 5.009921, 5.004006, 5.001504, 5.000525, 5.000171, 5.000052, 
    5.000016, 5.000004, 5, 5, 5,
  // momentumX(3,15, 0-49)
    5, 5, 5, 5, 5.000005, 5.00002, 5.000069, 5.000233, 5.000735, 5.002163, 
    5.005921, 5.015044, 5.035314, 5.076136, 5.14962, 5.26931, 5.461556, 
    5.608839, 5.731626, 5.821412, 5.873544, 5.920516, 5.942305, 5.950413, 
    5.955587, 5.957473, 5.955333, 5.949632, 5.940266, 5.915689, 5.863268, 
    5.801664, 5.698636, 5.56323, 5.414839, 5.276899, 5.167127, 5.091476, 
    5.045663, 5.020916, 5.00884, 5.003462, 5.001259, 5.000427, 5.000136, 
    5.000041, 5.000012, 5.000003, 5, 5,
  // momentumX(3,16, 0-49)
    5, 5, 5, 5.000002, 5.000011, 5.000041, 5.000143, 5.000468, 5.001436, 
    5.004103, 5.010897, 5.026792, 5.060598, 5.124972, 5.232549, 5.396155, 
    5.662586, 5.799902, 5.878317, 5.906157, 5.892824, 5.879972, 5.850737, 
    5.821409, 5.806584, 5.801819, 5.806024, 5.819709, 5.846377, 5.869823, 
    5.871604, 5.866385, 5.813318, 5.711125, 5.5706, 5.414839, 5.271254, 
    5.159427, 5.084641, 5.040899, 5.018124, 5.00741, 5.002808, 5.000989, 
    5.000327, 5.000101, 5.00003, 5.000008, 5.000001, 5,
  // momentumX(3,17, 0-49)
    5, 5, 5.000001, 5.000005, 5.000021, 5.000075, 5.000259, 5.000828, 
    5.002479, 5.006911, 5.017881, 5.042683, 5.093165, 5.18362, 5.322259, 
    5.521502, 5.866402, 5.969814, 5.983183, 5.936786, 5.854723, 5.780489, 
    5.701207, 5.636169, 5.601222, 5.58957, 5.600065, 5.632699, 5.692458, 
    5.76054, 5.814003, 5.863031, 5.867137, 5.816883, 5.711125, 5.56323, 
    5.400769, 5.25464, 5.144711, 5.0741, 5.034512, 5.014745, 5.005819, 
    5.00213, 5.000726, 5.000232, 5.00007, 5.00002, 5.000005, 5,
  // momentumX(3,18, 0-49)
    5, 5, 5.000002, 5.000009, 5.000031, 5.000117, 5.000395, 5.001246, 
    5.003667, 5.010052, 5.025521, 5.059556, 5.126149, 5.238306, 5.394081, 
    5.615667, 6.035935, 6.101533, 6.04922, 5.929343, 5.78085, 5.644381, 
    5.515065, 5.414158, 5.357251, 5.337825, 5.354997, 5.407474, 5.498516, 
    5.607554, 5.707836, 5.802571, 5.86004, 5.867137, 5.813318, 5.698636, 
    5.540854, 5.372893, 5.228083, 5.124352, 5.061041, 5.027278, 5.011199, 
    5.004254, 5.001501, 5.000495, 5.000153, 5.000045, 5.000013, 5.000002,
  // momentumX(3,19, 0-49)
    5, 5, 5.000002, 5.000011, 5.000038, 5.00014, 5.000471, 5.001475, 
    5.004326, 5.011827, 5.029943, 5.069492, 5.145236, 5.266404, 5.417098, 
    5.657688, 6.133231, 6.183744, 6.085767, 5.90326, 5.691944, 5.490312, 
    5.308599, 5.169163, 5.086947, 5.058302, 5.082806, 5.156998, 5.279012, 
    5.426208, 5.569045, 5.70021, 5.80257, 5.863031, 5.866385, 5.801664, 
    5.672307, 5.502812, 5.331985, 5.193449, 5.100338, 5.046923, 5.020027, 
    5.007874, 5.00287, 5.000974, 5.000309, 5.000092, 5.000025, 5.000007,
  // momentumX(3,20, 0-49)
    5, 5, 5.000001, 5.000006, 5.000022, 5.000076, 5.000246, 5.000745, 
    5.002099, 5.005454, 5.012992, 5.028082, 5.054316, 5.092286, 5.134862, 0, 
    6.537839, 6.444597, 6.224334, 5.931908, 5.627497, 5.341224, 5.09673, 
    4.91181, 4.799217, 4.759322, 4.791854, 4.890079, 5.043821, 5.226887, 
    5.408791, 5.569041, 5.707834, 5.814003, 5.871604, 5.863268, 5.779329, 
    5.629799, 5.448622, 5.279824, 5.153577, 5.075142, 5.033274, 5.013503, 
    5.005065, 5.001767, 5.000576, 5.000175, 5.000051, 5.000014,
  // momentumX(3,21, 0-49)
    5, 5, 5, 5.000002, 5.000011, 5.000037, 5.000119, 5.000364, 5.001029, 
    5.002694, 5.006472, 5.01416, 5.027897, 5.048741, 5.073972, 0, 6.715348, 
    6.582877, 6.306049, 5.934135, 5.539999, 5.157746, 4.834559, 4.587932, 
    4.433352, 4.378251, 4.422956, 4.55676, 4.757838, 4.992012, 5.226871, 
    5.426194, 5.607547, 5.760535, 5.869822, 5.915688, 5.880161, 5.75981, 
    5.578391, 5.383534, 5.221547, 5.112823, 5.05154, 5.021459, 5.008235, 
    5.002935, 5.000975, 5.000303, 5.000089, 5.000024,
  // momentumX(3,22, 0-49)
    5, 5, 5, 5, 5.000004, 5.000016, 5.000052, 5.00016, 5.000462, 5.001224, 
    5.002986, 5.006641, 5.013321, 5.023751, 5.036767, 0, 6.819324, 6.665093, 
    6.350619, 5.917248, 5.445622, 4.973551, 4.571023, 4.255342, 4.050066, 
    3.976002, 4.036703, 4.214768, 4.470624, 4.757758, 5.043741, 5.278961, 
    5.498487, 5.692443, 5.846371, 5.940264, 5.951795, 5.867255, 5.69812, 
    5.488389, 5.29539, 5.155908, 5.073154, 5.0311, 5.012152, 5.004404, 
    5.001488, 5.000471, 5.000139, 5.000038,
  // momentumX(3,23, 0-49)
    5, 5, 5, 5, 5.000001, 5.000007, 5.000022, 5.00007, 5.000204, 5.000552, 
    5.001373, 5.003109, 5.006342, 5.011469, 5.017878, 0, 6.881858, 6.715767, 
    6.377157, 5.89924, 5.365091, 4.814788, 4.335211, 3.944315, 3.680533, 
    3.584269, 3.664799, 3.895799, 4.214448, 4.556406, 4.88979, 5.156824, 
    5.407378, 5.63265, 5.819686, 5.949622, 5.99874, 5.946925, 5.795018, 
    5.57985, 5.363815, 5.197576, 5.094623, 5.040833, 5.016148, 5.005916, 
    5.002019, 5.000645, 5.000192, 5.000054,
  // momentumX(3,24, 0-49)
    5, 5, 5, 5, 5, 5.000004, 5.000014, 5.000044, 5.000131, 5.000354, 
    5.000885, 5.002009, 5.004103, 5.00741, 5.011444, 0, 6.913795, 6.743283, 
    6.393038, 5.88919, 5.313772, 4.708361, 4.169513, 3.717096, 3.405324, 
    3.291309, 3.388295, 3.663615, 4.035308, 4.421719, 4.790909, 5.082253, 
    5.354696, 5.599913, 5.805953, 5.955301, 6.024744, 5.991959, 5.852164, 
    5.636593, 5.40835, 5.225728, 5.109491, 5.047673, 5.018981, 5.006993, 
    5.0024, 5.000771, 5.00023, 5.000065,
  // momentumX(3,25, 0-49)
    5, 5, 5, 5, 5.000001, 5.000007, 5.000023, 5.000068, 5.000196, 5.000519, 
    5.001256, 5.00277, 5.005505, 5.009689, 5.014659, 0, 6.917509, 6.746934, 
    6.394336, 5.883124, 5.294426, 4.670211, 4.109842, 3.634244, 3.304592, 
    3.184185, 3.287201, 3.579186, 3.97121, 4.374317, 4.756428, 5.056643, 
    5.336924, 5.589113, 5.801601, 5.957374, 6.033497, 6.007074, 5.871552, 
    5.656174, 5.423996, 5.235758, 5.114835, 5.050141, 5.020005, 5.007383, 
    5.002537, 5.000815, 5.000245, 5.000069,
  // momentumX(3,26, 0-49)
    5, 5, 5, 5, 5.000005, 5.000018, 5.000054, 5.000162, 5.000451, 5.001157, 
    5.00272, 5.005827, 5.011258, 5.019319, 5.028754, 0, 6.889607, 6.723534, 
    6.378369, 5.879577, 5.308405, 4.705863, 4.168527, 3.716762, 3.405225, 
    3.291283, 3.388287, 3.663613, 4.035307, 4.421719, 4.790908, 5.082252, 
    5.354695, 5.599913, 5.805953, 5.955301, 6.024744, 5.991959, 5.852164, 
    5.636593, 5.40835, 5.225728, 5.109491, 5.047673, 5.018981, 5.006993, 
    5.0024, 5.000771, 5.00023, 5.000065,
  // momentumX(3,27, 0-49)
    5, 5, 5, 5.000003, 5.000013, 5.000042, 5.000131, 5.000385, 5.001048, 
    5.002628, 5.006048, 5.012661, 5.02387, 5.039977, 5.058367, 0, 6.826754, 
    6.670672, 6.343395, 5.876875, 5.352436, 4.808751, 4.332749, 3.943442, 
    3.680258, 3.58419, 3.664778, 3.895793, 4.214446, 4.556406, 4.889789, 
    5.156823, 5.407378, 5.63265, 5.819686, 5.949621, 5.99874, 5.946925, 
    5.795018, 5.57985, 5.363815, 5.197576, 5.094623, 5.040833, 5.016148, 
    5.005916, 5.002019, 5.000645, 5.000192, 5.000054,
  // momentumX(3,28, 0-49)
    5, 5, 5.000001, 5.000009, 5.000028, 5.000093, 5.000291, 5.000842, 
    5.002254, 5.005562, 5.012565, 5.025754, 5.047345, 5.076943, 5.108829, 0, 
    6.720564, 6.584433, 6.289873, 5.876649, 5.422355, 4.96215, 4.566208, 
    4.253551, 4.049467, 3.975818, 4.036649, 4.214753, 4.470621, 4.757757, 
    5.04374, 5.27896, 5.498487, 5.692443, 5.846371, 5.940264, 5.951794, 
    5.867256, 5.69812, 5.488389, 5.29539, 5.155908, 5.073154, 5.0311, 
    5.012152, 5.004404, 5.001488, 5.000471, 5.000139, 5.000038,
  // momentumX(3,29, 0-49)
    5, 5, 5.000004, 5.000016, 5.000057, 5.000186, 5.000579, 5.001659, 
    5.004405, 5.010764, 5.024003, 5.048273, 5.086257, 5.134563, 5.180684, 0, 
    6.556565, 6.454806, 6.209808, 5.869759, 5.502885, 5.139183, 4.826483, 
    4.584808, 4.432256, 4.377896, 4.422847, 4.556728, 4.757828, 4.99201, 
    5.226871, 5.426193, 5.607547, 5.760535, 5.869822, 5.915688, 5.880161, 
    5.75981, 5.578391, 5.383534, 5.221547, 5.112823, 5.05154, 5.021459, 
    5.008235, 5.002935, 5.000975, 5.000303, 5.000089, 5.000024,
  // momentumX(3,30, 0-49)
    5, 5.000002, 5.000008, 5.000027, 5.0001, 5.000338, 5.001072, 5.003178, 
    5.008781, 5.022519, 5.053143, 5.113769, 5.216212, 5.355342, 5.494076, 
    5.709598, 6.125762, 6.156536, 6.034242, 5.81732, 5.566053, 5.311934, 
    5.084235, 4.906974, 4.7975, 4.758753, 4.791675, 4.890025, 5.043805, 
    5.226883, 5.40879, 5.569041, 5.707834, 5.814003, 5.871604, 5.863268, 
    5.779329, 5.629799, 5.448622, 5.279824, 5.153577, 5.075142, 5.033274, 
    5.013503, 5.005065, 5.001767, 5.000576, 5.000175, 5.000051, 5.000014,
  // momentumX(3,31, 0-49)
    5, 5.000001, 5.000006, 5.000023, 5.000086, 5.000294, 5.000936, 5.002785, 
    5.007725, 5.019886, 5.047167, 5.101953, 5.197631, 5.337241, 5.499212, 
    5.707389, 6.101362, 6.130861, 6.032712, 5.862597, 5.666519, 5.477023, 
    5.3025, 5.166655, 5.086007, 5.057975, 5.082697, 5.156963, 5.279002, 
    5.426205, 5.569045, 5.70021, 5.80257, 5.863031, 5.866385, 5.801664, 
    5.672307, 5.502812, 5.331985, 5.193449, 5.100338, 5.046923, 5.020027, 
    5.007874, 5.00287, 5.000974, 5.000309, 5.000092, 5.000025, 5.000007,
  // momentumX(3,32, 0-49)
    5, 5, 5.000003, 5.000016, 5.000057, 5.000198, 5.000641, 5.001941, 
    5.005484, 5.014384, 5.034873, 5.077482, 5.155878, 5.27987, 5.442998, 
    5.649105, 5.993998, 6.054826, 6.009722, 5.902009, 5.764829, 5.636314, 
    5.511456, 5.412694, 5.356704, 5.337633, 5.354934, 5.407454, 5.49851, 
    5.607553, 5.707836, 5.802571, 5.86004, 5.867137, 5.813318, 5.698636, 
    5.540854, 5.372893, 5.228083, 5.124352, 5.061041, 5.027278, 5.011199, 
    5.004254, 5.001501, 5.000495, 5.000153, 5.000045, 5.000013, 5.000002,
  // momentumX(3,33, 0-49)
    5, 5, 5.000001, 5.000009, 5.000031, 5.000113, 5.000374, 5.00116, 
    5.003356, 5.009038, 5.022561, 5.051877, 5.108922, 5.206487, 5.349631, 
    5.540675, 5.829793, 5.934906, 5.95664, 5.919773, 5.845279, 5.775891, 
    5.699202, 5.635369, 5.600927, 5.589468, 5.600031, 5.632689, 5.692454, 
    5.760539, 5.814003, 5.863031, 5.867137, 5.816883, 5.711125, 5.563231, 
    5.400769, 5.25464, 5.144711, 5.0741, 5.034512, 5.014745, 5.005819, 
    5.00213, 5.000726, 5.000232, 5.00007, 5.00002, 5.000005, 5,
  // momentumX(3,34, 0-49)
    5, 5, 5, 5.000003, 5.000016, 5.000058, 5.000192, 5.000611, 5.001822, 
    5.00506, 5.013054, 5.031149, 5.068315, 5.13659, 5.246739, 5.405913, 
    5.637955, 5.777564, 5.862308, 5.896429, 5.887648, 5.877523, 5.849693, 
    5.821001, 5.806437, 5.801769, 5.806009, 5.819705, 5.846376, 5.869823, 
    5.871605, 5.866385, 5.813318, 5.711125, 5.5706, 5.414839, 5.271254, 
    5.159427, 5.084641, 5.040899, 5.018124, 5.00741, 5.002808, 5.000989, 
    5.000327, 5.000101, 5.00003, 5.000008, 5.000001, 5,
  // momentumX(3,35, 0-49)
    5, 5, 5, 5.000001, 5.000007, 5.000026, 5.000089, 5.00029, 5.000893, 
    5.002561, 5.006839, 5.016948, 5.038792, 5.081545, 5.156356, 5.273779, 
    5.448004, 5.596495, 5.722991, 5.816328, 5.870923, 5.919303, 5.941797, 
    5.950219, 5.955517, 5.957448, 5.955325, 5.949628, 5.940266, 5.915689, 
    5.863268, 5.801664, 5.698636, 5.56323, 5.414839, 5.276899, 5.167127, 
    5.091476, 5.045663, 5.020916, 5.00884, 5.003462, 5.001259, 5.000427, 
    5.000136, 5.000041, 5.000012, 5.000003, 5, 5,
  // momentumX(3,36, 0-49)
    5, 5, 5, 5, 5.000002, 5.000011, 5.000038, 5.000125, 5.000399, 5.001182, 
    5.00327, 5.008418, 5.020082, 5.044224, 5.089479, 5.166116, 5.285483, 
    5.41548, 5.55173, 5.678836, 5.782701, 5.881738, 5.952456, 5.998994, 
    6.024836, 6.033529, 6.024755, 5.998743, 5.951795, 5.880162, 5.77933, 
    5.672307, 5.540854, 5.400769, 5.271254, 5.167127, 5.093842, 5.048205, 
    5.022761, 5.009921, 5.004006, 5.001504, 5.000525, 5.000171, 5.000052, 
    5.000016, 5.000004, 5, 5, 5,
  // momentumX(3,37, 0-49)
    5, 5, 5, 5, 5, 5.000004, 5.000015, 5.000051, 5.000163, 5.000501, 
    5.001435, 5.003837, 5.00953, 5.021924, 5.046564, 5.091146, 5.164802, 
    5.260377, 5.377213, 5.50543, 5.631152, 5.760442, 5.867519, 5.947026, 
    5.991995, 6.007086, 5.991962, 5.946927, 5.867255, 5.75981, 5.629799, 
    5.502812, 5.372893, 5.25464, 5.159427, 5.091476, 5.048205, 5.023404, 
    5.010503, 5.004369, 5.001688, 5.000608, 5.000204, 5.000064, 5.00002, 
    5.000005, 5, 5, 5, 5,
  // momentumX(3,38, 0-49)
    5, 5, 5, 5, 5, 5, 5.000005, 5.00002, 5.000062, 5.000195, 5.00058, 
    5.001613, 5.004166, 5.009988, 5.022183, 5.045549, 5.086459, 5.146701, 
    5.229607, 5.33292, 5.449109, 5.578621, 5.698215, 5.795055, 5.852177, 
    5.871556, 5.852166, 5.79502, 5.69812, 5.578392, 5.448622, 5.331985, 
    5.228083, 5.144711, 5.084641, 5.045663, 5.022761, 5.010503, 5.004496, 
    5.001788, 5.000662, 5.000228, 5.000074, 5.000023, 5.000007, 5.000001, 5, 
    5, 5, 5,
  // momentumX(3,39, 0-49)
    5, 5, 5, 5, 5, 5, 5.000001, 5.000007, 5.000022, 5.000071, 5.000218, 
    5.000627, 5.001684, 5.004201, 5.00973, 5.020876, 5.04146, 5.074723, 
    5.124831, 5.193744, 5.27998, 5.383608, 5.48842, 5.579863, 5.636596, 
    5.656175, 5.636593, 5.57985, 5.488389, 5.383535, 5.279824, 5.193449, 
    5.124352, 5.0741, 5.040899, 5.020916, 5.009921, 5.004369, 5.001788, 
    5.000681, 5.000242, 5.00008, 5.000025, 5.000008, 5.000002, 5, 5, 5, 5, 5,
  // momentumX(3,40, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000008, 5.000024, 5.000075, 5.000226, 
    5.00063, 5.001637, 5.003948, 5.008826, 5.018284, 5.034691, 5.061178, 
    5.100423, 5.153621, 5.221567, 5.295398, 5.363819, 5.408352, 5.423996, 
    5.408351, 5.363815, 5.29539, 5.221547, 5.153577, 5.100338, 5.061041, 
    5.034512, 5.018124, 5.00884, 5.004006, 5.001688, 5.000662, 5.000242, 
    5.000082, 5.000026, 5.000008, 5.000002, 5, 5, 5, 5, 5, 5,
  // momentumX(3,41, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000008, 5.000024, 5.000076, 5.00022, 
    5.000594, 5.001486, 5.003456, 5.007452, 5.014793, 5.027314, 5.046945, 
    5.075154, 5.112829, 5.15591, 5.197577, 5.225729, 5.235758, 5.225728, 
    5.197576, 5.155908, 5.112823, 5.075142, 5.046923, 5.027278, 5.014745, 
    5.00741, 5.003462, 5.001504, 5.000608, 5.000228, 5.00008, 5.000026, 
    5.000009, 5.000002, 5, 5, 5, 5, 5, 5, 5,
  // momentumX(3,42, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000008, 5.000024, 5.000072, 
    5.0002, 5.000521, 5.001258, 5.002819, 5.00583, 5.011209, 5.020034, 
    5.033277, 5.051541, 5.073155, 5.094623, 5.109491, 5.114835, 5.109491, 
    5.094623, 5.073154, 5.05154, 5.033274, 5.020027, 5.011199, 5.005819, 
    5.002808, 5.001259, 5.000525, 5.000204, 5.000074, 5.000025, 5.000008, 
    5.000002, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumX(3,43, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000008, 5.000023, 5.000063, 
    5.00017, 5.000428, 5.000993, 5.002134, 5.004256, 5.007876, 5.013503, 
    5.021459, 5.0311, 5.040833, 5.047673, 5.050141, 5.047673, 5.040833, 
    5.0311, 5.021459, 5.013503, 5.007874, 5.004254, 5.00213, 5.000989, 
    5.000427, 5.000171, 5.000064, 5.000023, 5.000008, 5.000002, 5, 5, 5, 5, 
    5, 5, 5, 5, 5,
  // momentumX(3,44, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000007, 5.00002, 5.000052, 
    5.000136, 5.000328, 5.000727, 5.001502, 5.002871, 5.005065, 5.008235, 
    5.012152, 5.016148, 5.018981, 5.020005, 5.018981, 5.016148, 5.012152, 
    5.008235, 5.005065, 5.00287, 5.001501, 5.000726, 5.000327, 5.000136, 
    5.000052, 5.00002, 5.000007, 5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumX(3,45, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000005, 5.000016, 
    5.000041, 5.000101, 5.000232, 5.000495, 5.000975, 5.001767, 5.002935, 
    5.004404, 5.005916, 5.006993, 5.007383, 5.006993, 5.005916, 5.004404, 
    5.002935, 5.001767, 5.000974, 5.000495, 5.000232, 5.000101, 5.000041, 
    5.000016, 5.000005, 5.000001, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumX(3,46, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000004, 5.000012, 5.00003, 
    5.00007, 5.000153, 5.000309, 5.000576, 5.000975, 5.001488, 5.002019, 
    5.0024, 5.002537, 5.0024, 5.002019, 5.001488, 5.000975, 5.000576, 
    5.000309, 5.000153, 5.00007, 5.00003, 5.000012, 5.000004, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5,
  // momentumX(3,47, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000003, 5.000008, 5.00002, 
    5.000045, 5.000092, 5.000175, 5.000303, 5.000471, 5.000645, 5.000771, 
    5.000815, 5.000771, 5.000645, 5.000471, 5.000303, 5.000175, 5.000092, 
    5.000045, 5.00002, 5.000008, 5.000003, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5,
  // momentumX(3,48, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000005, 
    5.000013, 5.000025, 5.000051, 5.000089, 5.000139, 5.000192, 5.000231, 
    5.000245, 5.000231, 5.000192, 5.000139, 5.000089, 5.000051, 5.000025, 
    5.000013, 5.000005, 5.000001, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumX(3,49, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000006, 
    5.000012, 5.000023, 5.000038, 5.000055, 5.000067, 5.000071, 5.000067, 
    5.000055, 5.000038, 5.000023, 5.000012, 5.000006, 5.000002, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumX(4,0, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000006, 5.000013, 
    5.000028, 5.000057, 5.000112, 5.000206, 5.000354, 5.000569, 5.00085, 
    5.001171, 5.001479, 5.001697, 5.001776, 5.001697, 5.001479, 5.001171, 
    5.00085, 5.000569, 5.000354, 5.000206, 5.000112, 5.000057, 5.000028, 
    5.000013, 5.000006, 5.000001, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumX(4,1, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000003, 5.000008, 5.000018, 5.000039, 
    5.000082, 5.000166, 5.000319, 5.000575, 5.000974, 5.001544, 5.002285, 
    5.003127, 5.003933, 5.004504, 5.00471, 5.004504, 5.003933, 5.003127, 
    5.002285, 5.001544, 5.000974, 5.000575, 5.000319, 5.000166, 5.000082, 
    5.000038, 5.000018, 5.000008, 5.000003, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumX(4,2, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000004, 5.00001, 5.000022, 5.00005, 
    5.000111, 5.000235, 5.000467, 5.000876, 5.001545, 5.002564, 5.003994, 
    5.005826, 5.00789, 5.009855, 5.011244, 5.011746, 5.011244, 5.009855, 
    5.00789, 5.005825, 5.003993, 5.002563, 5.001543, 5.000874, 5.000466, 
    5.000235, 5.000111, 5.00005, 5.000022, 5.00001, 5.000004, 5, 5, 5, 5, 5, 
    5, 5, 5, 5,
  // momentumX(4,3, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000005, 5.000011, 5.000026, 5.000062, 
    5.000142, 5.000312, 5.000645, 5.001252, 5.002286, 5.003933, 5.006382, 
    5.00975, 5.014007, 5.018755, 5.023253, 5.026416, 5.027557, 5.026416, 
    5.023252, 5.018755, 5.014006, 5.009748, 5.006378, 5.003928, 5.002279, 
    5.001247, 5.000645, 5.000314, 5.000144, 5.000063, 5.000027, 5.000011, 
    5.000005, 5.000001, 5, 5, 5, 5, 5, 5, 5,
  // momentumX(4,4, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000005, 5.000012, 5.00003, 5.000073, 
    5.000174, 5.000391, 5.000835, 5.001678, 5.003172, 5.005635, 5.009448, 
    5.014966, 5.022386, 5.031617, 5.041789, 5.051358, 5.058033, 5.060435, 
    5.058033, 5.051356, 5.041786, 5.031611, 5.022377, 5.014951, 5.009429, 
    5.005613, 5.003155, 5.001675, 5.00084, 5.000397, 5.000178, 5.000076, 
    5.000031, 5.000013, 5.000005, 5.000001, 5, 5, 5, 5, 5, 5,
  // momentumX(4,5, 0-49)
    5, 5, 5, 5, 5, 5, 5.000002, 5.000006, 5.000013, 5.000031, 5.000082, 
    5.0002, 5.000464, 5.00102, 5.002115, 5.004128, 5.00759, 5.013093, 
    5.021336, 5.032907, 5.048047, 5.066521, 5.086531, 5.105149, 5.117974, 
    5.122565, 5.117973, 5.105145, 5.086521, 5.066501, 5.048014, 5.032856, 
    5.021269, 5.01302, 5.007533, 5.004119, 5.002128, 5.001039, 5.00048, 
    5.00021, 5.000087, 5.000034, 5.000014, 5.000006, 5.000002, 5, 5, 5, 5, 5,
  // momentumX(4,6, 0-49)
    5, 5, 5, 5, 5, 5.000001, 5.000006, 5.000013, 5.000033, 5.000086, 
    5.000218, 5.00052, 5.001176, 5.002513, 5.005054, 5.009583, 5.017104, 
    5.028571, 5.04509, 5.06742, 5.095617, 5.129127, 5.164507, 5.196824, 
    5.218638, 5.226384, 5.218632, 5.196807, 5.164472, 5.12906, 5.095507, 
    5.067253, 5.04487, 5.028332, 5.016919, 5.009551, 5.005095, 5.002568, 
    5.001224, 5.00055, 5.000236, 5.000094, 5.000036, 5.000015, 5.000007, 
    5.000002, 5, 5, 5, 5,
  // momentumX(4,7, 0-49)
    5, 5, 5, 5, 5, 5.000005, 5.000013, 5.000032, 5.000086, 5.000224, 
    5.000552, 5.001284, 5.002817, 5.005834, 5.011383, 5.020915, 5.036179, 
    5.058282, 5.0886, 5.12762, 5.174555, 5.228317, 5.28298, 5.331494, 
    5.363276, 5.374424, 5.363256, 5.331442, 5.282871, 5.228115, 5.174216, 
    5.12711, 5.08793, 5.057558, 5.035612, 5.020813, 5.011489, 5.00599, 
    5.002948, 5.001372, 5.000603, 5.00025, 5.000099, 5.000037, 5.000015, 
    5.000006, 5.000001, 5, 5, 5,
  // momentumX(4,8, 0-49)
    5, 5, 5, 5, 5.000004, 5.000011, 5.00003, 5.000083, 5.000219, 5.000553, 
    5.001321, 5.002983, 5.00635, 5.012745, 5.024074, 5.042771, 5.071508, 
    5.110453, 5.160557, 5.220954, 5.288945, 5.363122, 5.434719, 5.495795, 
    5.534249, 5.547521, 5.534192, 5.49565, 5.434417, 5.36256, 5.288007, 
    5.219527, 5.158675, 5.108407, 5.069887, 5.04248, 5.024346, 5.013159, 
    5.006711, 5.003231, 5.001469, 5.000631, 5.000257, 5.000099, 5.000036, 
    5.000014, 5.000005, 5.000001, 5, 5,
  // momentumX(4,9, 0-49)
    5, 5, 5, 5.000003, 5.00001, 5.000027, 5.000073, 5.000201, 5.000522, 
    5.001283, 5.002978, 5.006522, 5.013456, 5.026117, 5.047627, 5.081541, 
    5.131313, 5.193063, 5.26604, 5.346703, 5.429886, 5.515448, 5.592755, 
    5.65555, 5.693194, 5.705945, 5.693052, 5.655185, 5.592003, 5.51405, 
    5.427536, 5.343099, 5.261235, 5.187773, 5.12704, 5.0808, 5.048308, 
    5.027168, 5.014386, 5.00718, 5.00338, 5.001504, 5.000631, 5.00025, 
    5.000094, 5.000034, 5.000013, 5.000005, 5, 5,
  // momentumX(4,10, 0-49)
    5, 5, 5.000001, 5.000008, 5.000023, 5.000062, 5.000174, 5.000464, 
    5.001174, 5.002803, 5.006311, 5.01339, 5.026711, 5.050013, 5.087704, 
    5.143996, 5.222599, 5.309128, 5.400571, 5.490787, 5.573659, 5.653591, 
    5.720015, 5.770827, 5.799431, 5.808886, 5.799106, 5.770001, 5.718316, 
    5.65044, 5.568353, 5.482604, 5.389545, 5.296785, 5.212377, 5.142366, 
    5.089346, 5.052536, 5.028989, 5.015037, 5.007341, 5.00338, 5.001469, 
    5.000603, 5.000236, 5.000087, 5.000031, 5.000011, 5.000004, 5,
  // momentumX(4,11, 0-49)
    5, 5.000001, 5.000006, 5.000018, 5.000051, 5.000142, 5.000389, 5.00101, 
    5.002481, 5.005745, 5.012537, 5.025723, 5.049498, 5.089058, 5.149407, 
    5.233919, 5.346392, 5.451672, 5.547588, 5.628493, 5.690985, 5.747229, 
    5.788034, 5.816257, 5.830287, 5.834641, 5.829595, 5.814518, 5.784492, 
    5.740716, 5.680092, 5.611754, 5.524933, 5.425946, 5.324495, 5.230956, 
    5.153233, 5.094786, 5.05476, 5.029618, 5.015037, 5.00718, 5.003231, 
    5.001372, 5.00055, 5.00021, 5.000076, 5.000027, 5.00001, 5.000003,
  // momentumX(4,12, 0-49)
    5, 5.000003, 5.000013, 5.000038, 5.000109, 5.000305, 5.000814, 5.002055, 
    5.004901, 5.011015, 5.023273, 5.046094, 5.08526, 5.146695, 5.233996, 
    5.347453, 5.493467, 5.603019, 5.683767, 5.735504, 5.761001, 5.781113, 
    5.78789, 5.788424, 5.785759, 5.784305, 5.784378, 5.784986, 5.780982, 
    5.768596, 5.740397, 5.704315, 5.641876, 5.555245, 5.451858, 5.343374, 
    5.242486, 5.158862, 5.096653, 5.05476, 5.028989, 5.014386, 5.006711, 
    5.002948, 5.001224, 5.00048, 5.000178, 5.000063, 5.000022, 5.000008,
  // momentumX(4,13, 0-49)
    5.000001, 5.000009, 5.000026, 5.000077, 5.000224, 5.000611, 5.001587, 
    5.003901, 5.009038, 5.019696, 5.040237, 5.07673, 5.135884, 5.222372, 
    5.33526, 5.470407, 5.644621, 5.740721, 5.789155, 5.798397, 5.778439, 
    5.757261, 5.727443, 5.699325, 5.679906, 5.672492, 5.677281, 5.692876, 
    5.71471, 5.734662, 5.742108, 5.744841, 5.718772, 5.661288, 5.574646, 
    5.467301, 5.352917, 5.246391, 5.158862, 5.094786, 5.052536, 5.027167, 
    5.013159, 5.00599, 5.002568, 5.001039, 5.000397, 5.000144, 5.00005, 
    5.000018,
  // momentumX(4,14, 0-49)
    5.000004, 5.000016, 5.000051, 5.00015, 5.000423, 5.001134, 5.002876, 
    5.006879, 5.015491, 5.032723, 5.064547, 5.118182, 5.199555, 5.309104, 
    5.438466, 5.581018, 5.776528, 5.845946, 5.853991, 5.817026, 5.75099, 
    5.688416, 5.622475, 5.56643, 5.530651, 5.517122, 5.525881, 5.554883, 
    5.600159, 5.649828, 5.690797, 5.731436, 5.745387, 5.726641, 5.672071, 
    5.58408, 5.472425, 5.352917, 5.242486, 5.153233, 5.089346, 5.048308, 
    5.024346, 5.011489, 5.005095, 5.002128, 5.00084, 5.000314, 5.000111, 
    5.000039,
  // momentumX(4,15, 0-49)
    5.000009, 5.00003, 5.000093, 5.000268, 5.000741, 5.001943, 5.004808, 
    5.011213, 5.02456, 5.050291, 5.095673, 5.167803, 5.269303, 5.393564, 
    5.523967, 5.657652, 5.868953, 5.907986, 5.878179, 5.799743, 5.692262, 
    5.590435, 5.489555, 5.406311, 5.354075, 5.333925, 5.345757, 5.386508, 
    5.452232, 5.527853, 5.598085, 5.67159, 5.722934, 5.744675, 5.730055, 
    5.67552, 5.58408, 5.467301, 5.343374, 5.230956, 5.142365, 5.080799, 
    5.04248, 5.020813, 5.009551, 5.004119, 5.001675, 5.000645, 5.000236, 
    5.000084,
  // momentumX(4,16, 0-49)
    5.000016, 5.000051, 5.000154, 5.000436, 5.001185, 5.003041, 5.007361, 
    5.016769, 5.035784, 5.071095, 5.130445, 5.218989, 5.333667, 5.459665, 
    5.573878, 5.686548, 5.908281, 5.92311, 5.866307, 5.756901, 5.615705, 
    5.477578, 5.342819, 5.232497, 5.162915, 5.135132, 5.148944, 5.199866, 
    5.28306, 5.380913, 5.476108, 5.57633, 5.659531, 5.718256, 5.744269, 
    5.730054, 5.672071, 5.574646, 5.451857, 5.324495, 5.212377, 5.12704, 
    5.069887, 5.035612, 5.016918, 5.007533, 5.003155, 5.001247, 5.000467, 
    5.000169,
  // momentumX(4,17, 0-49)
    5.000024, 5.000076, 5.000226, 5.000637, 5.0017, 5.004287, 5.01019, 
    5.022752, 5.047452, 5.091729, 5.162721, 5.26203, 5.379788, 5.493896, 
    5.577772, 5.66574, 5.886785, 5.890759, 5.822771, 5.696401, 5.531397, 
    5.360797, 5.193435, 5.055688, 4.967145, 4.93014, 4.944488, 5.003893, 
    5.101617, 5.218238, 5.334838, 5.456188, 5.56532, 5.655404, 5.718253, 
    5.744672, 5.726639, 5.661288, 5.555245, 5.425946, 5.296785, 5.187774, 
    5.108407, 5.057558, 5.028332, 5.01302, 5.005613, 5.00228, 5.000876, 
    5.000325,
  // momentumX(4,18, 0-49)
    5.000031, 5.000098, 5.00029, 5.000809, 5.002132, 5.005311, 5.012467, 
    5.027443, 5.05629, 5.106589, 5.184099, 5.286392, 5.397364, 5.489583, 
    5.535452, 5.605662, 5.800894, 5.810308, 5.749249, 5.622153, 5.445377, 
    5.247847, 5.050285, 4.884759, 4.775092, 4.726635, 4.739514, 4.805339, 
    4.914531, 5.046517, 5.181646, 5.319603, 5.449533, 5.565309, 5.659521, 
    5.722928, 5.745382, 5.718771, 5.641876, 5.524933, 5.389545, 5.261234, 
    5.158674, 5.08793, 5.04487, 5.021269, 5.009429, 5.003929, 5.001545, 
    5.000584,
  // momentumX(4,19, 0-49)
    5.000033, 5.000104, 5.000303, 5.000842, 5.002212, 5.00549, 5.012845, 
    5.02818, 5.057574, 5.108389, 5.185361, 5.283393, 5.381967, 5.449668, 
    5.45941, 5.528225, 5.651516, 5.679839, 5.644249, 5.534561, 5.360603, 
    5.14432, 4.920958, 4.727758, 4.594412, 4.531527, 4.540184, 4.609795, 
    4.727152, 4.870959, 5.022038, 5.172999, 5.319552, 5.45614, 5.576295, 
    5.67157, 5.731426, 5.744835, 5.704313, 5.611754, 5.482604, 5.343098, 
    5.219526, 5.12711, 5.067253, 5.032856, 5.014951, 5.00638, 5.002567, 
    5.000986,
  // momentumX(4,20, 0-49)
    5.000022, 5.000071, 5.000206, 5.000566, 5.001461, 5.003547, 5.008075, 
    5.017149, 5.033758, 5.061057, 5.100434, 5.148736, 5.196876, 5.232886, 
    5.249486, 0, 5.72522, 5.722096, 5.663104, 5.536474, 5.342846, 5.092929, 
    4.832631, 4.601823, 4.436234, 4.352537, 4.352442, 4.422397, 4.544476, 
    4.696456, 4.860911, 5.021814, 5.181428, 5.334681, 5.476007, 5.598027, 
    5.690766, 5.742093, 5.74039, 5.680089, 5.568351, 5.427535, 5.288007, 
    5.174216, 5.095507, 5.048014, 5.022378, 5.00975, 5.003997, 5.001556,
  // momentumX(4,21, 0-49)
    5.000014, 5.000044, 5.000126, 5.000348, 5.000903, 5.002204, 5.005051, 
    5.010816, 5.021541, 5.039646, 5.06693, 5.102845, 5.142964, 5.179457, 
    5.204838, 0, 5.693264, 5.683771, 5.624491, 5.49779, 5.296422, 5.020554, 
    4.725423, 4.45422, 4.252345, 4.146114, 4.139155, 4.214416, 4.347202, 
    4.512626, 4.695527, 4.870046, 5.045835, 5.217789, 5.380641, 5.527698, 
    5.649745, 5.734621, 5.768576, 5.740706, 5.650436, 5.514049, 5.36256, 
    5.228116, 5.12906, 5.066501, 5.031611, 5.014006, 5.005826, 5.002292,
  // momentumX(4,22, 0-49)
    5.000008, 5.000024, 5.000072, 5.000199, 5.000521, 5.00129, 5.002997, 
    5.006517, 5.013214, 5.024857, 5.043125, 5.068581, 5.099402, 5.130821, 
    5.156437, 0, 5.645344, 5.631002, 5.571152, 5.445369, 5.241158, 4.948497, 
    4.63036, 4.328893, 4.096667, 3.969621, 3.954431, 4.03174, 4.170502, 
    4.343932, 4.540859, 4.72441, 4.91267, 5.100444, 5.282361, 5.451836, 
    5.599946, 5.7146, 5.780928, 5.784469, 5.718306, 5.591999, 5.434416, 
    5.28287, 5.164471, 5.086521, 5.041785, 5.018754, 5.007888, 5.003124,
  // momentumX(4,23, 0-49)
    5.000003, 5.000014, 5.000041, 5.000118, 5.000312, 5.000783, 5.001848, 
    5.004087, 5.008446, 5.016229, 5.028857, 5.047226, 5.070715, 5.096325, 
    5.118713, 0, 5.596464, 5.578844, 5.518146, 5.392861, 5.187092, 4.88203, 
    4.546795, 4.220427, 3.96124, 3.815448, 3.794108, 3.875613, 4.021391, 
    4.202407, 4.412063, 4.602664, 4.800696, 5.001018, 5.198163, 5.385542, 
    5.554357, 5.692601, 5.784849, 5.814455, 5.769972, 5.655174, 5.495645, 
    5.33144, 5.196806, 5.105144, 5.051356, 5.023251, 5.009851, 5.003916,
  // momentumX(4,24, 0-49)
    5.000002, 5.000011, 5.000033, 5.000093, 5.000248, 5.000626, 5.001483, 
    5.003294, 5.006839, 5.01322, 5.023686, 5.039129, 5.059257, 5.081702, 
    5.101663, 0, 5.556334, 5.537187, 5.476232, 5.351586, 5.145324, 4.83245, 
    4.485684, 4.140932, 3.860631, 3.700632, 3.676901, 3.765053, 3.9187, 
    4.106887, 4.327, 4.52336, 4.728728, 4.937836, 5.14499, 5.343493, 
    5.524635, 5.676622, 5.784046, 5.829436, 5.799034, 5.693022, 5.534179, 
    5.363252, 5.21863, 5.117971, 5.058032, 5.026413, 5.011236, 5.004478,
  // momentumX(4,25, 0-49)
    5.000005, 5.000016, 5.000045, 5.000125, 5.000327, 5.000806, 5.00187, 
    5.004066, 5.00826, 5.015623, 5.027387, 5.044277, 5.06568, 5.088906, 
    5.109101, 0, 5.530094, 5.511153, 5.450953, 5.327627, 5.122614, 4.808633, 
    4.459426, 4.109352, 3.822037, 3.657288, 3.633398, 3.724782, 3.881723, 
    4.07268, 4.296721, 4.495244, 4.70334, 4.915673, 5.126443, 5.328887, 
    5.514308, 5.670983, 5.783531, 5.834264, 5.808712, 5.705871, 5.54749, 
    5.374413, 5.226382, 5.122564, 5.060434, 5.027554, 5.011736, 5.004682,
  // momentumX(4,26, 0-49)
    5.00001, 5.00003, 5.000083, 5.000225, 5.000573, 5.001377, 5.003111, 
    5.006579, 5.012978, 5.023774, 5.040254, 5.062696, 5.089457, 5.116624, 
    5.138906, 0, 5.520136, 5.503262, 5.445169, 5.324215, 5.122498, 4.814704, 
    4.473166, 4.133136, 3.856438, 3.698707, 3.676142, 3.764788, 3.918613, 
    4.10686, 4.326991, 4.523357, 4.728727, 4.937836, 5.144989, 5.343493, 
    5.524634, 5.676622, 5.784046, 5.829436, 5.799034, 5.693022, 5.534179, 
    5.363252, 5.21863, 5.117971, 5.058032, 5.026413, 5.011236, 5.004478,
  // momentumX(4,27, 0-49)
    5.000019, 5.000056, 5.000157, 5.000415, 5.001042, 5.002456, 5.005435, 
    5.011232, 5.021597, 5.038417, 5.062864, 5.094123, 5.128512, 5.160077, 
    5.183197, 0, 5.526995, 5.513671, 5.458173, 5.339542, 5.142099, 4.846486, 
    4.52138, 4.204391, 3.952483, 3.811342, 3.79244, 3.875007, 4.021184, 
    4.202338, 4.412041, 4.602656, 4.800694, 5.001017, 5.198163, 5.385541, 
    5.554357, 5.692601, 5.784849, 5.814455, 5.769972, 5.655174, 5.495645, 
    5.33144, 5.196806, 5.105144, 5.051356, 5.023251, 5.009851, 5.003916,
  // momentumX(4,28, 0-49)
    5.000035, 5.0001, 5.000277, 5.000724, 5.001793, 5.004173, 5.009095, 
    5.018476, 5.034788, 5.060286, 5.095444, 5.137174, 5.178433, 5.210751, 
    5.229156, 0, 5.549765, 5.540964, 5.487337, 5.369511, 5.17579, 4.895623, 
    4.591888, 4.304254, 4.082989, 3.963053, 3.951664, 4.030686, 4.170128, 
    4.343802, 4.540814, 4.724395, 4.912664, 5.100442, 5.28236, 5.451836, 
    5.599946, 5.7146, 5.780928, 5.784469, 5.718305, 5.591999, 5.434416, 
    5.28287, 5.164471, 5.086521, 5.041785, 5.018754, 5.007888, 5.003124,
  // momentumX(4,29, 0-49)
    5.000054, 5.000159, 5.000442, 5.001153, 5.00284, 5.006568, 5.014205, 
    5.028555, 5.05294, 5.08968, 5.137436, 5.189026, 5.232651, 5.257787, 
    5.262488, 0, 5.584862, 5.579939, 5.525392, 5.405305, 5.214372, 4.952533, 
    4.675216, 4.421723, 4.234072, 4.137152, 4.135252, 4.212865, 4.346626, 
    4.51242, 4.695455, 4.870021, 5.045825, 5.217786, 5.380639, 5.527698, 
    5.649745, 5.734621, 5.768576, 5.740706, 5.650436, 5.514049, 5.36256, 
    5.228116, 5.12906, 5.066501, 5.031611, 5.014006, 5.005826, 5.002292,
  // momentumX(4,30, 0-49)
    5.000076, 5.000227, 5.000637, 5.001688, 5.004233, 5.010009, 5.022226, 
    5.046075, 5.08837, 5.154881, 5.244466, 5.342824, 5.423133, 5.457164, 
    5.429102, 5.460217, 5.513269, 5.527208, 5.492916, 5.390181, 5.221525, 
    4.998848, 4.766492, 4.560466, 4.413423, 4.341393, 4.347546, 4.42042, 
    4.543725, 4.696185, 4.860814, 5.02178, 5.181416, 5.334677, 5.476006, 
    5.598026, 5.690766, 5.742093, 5.74039, 5.680089, 5.568351, 5.427535, 
    5.288007, 5.174216, 5.095507, 5.048014, 5.022378, 5.00975, 5.003997, 
    5.001556,
  // momentumX(4,31, 0-49)
    5.000073, 5.000221, 5.000621, 5.001653, 5.00416, 5.009876, 5.02202, 
    5.045835, 5.088351, 5.155962, 5.249051, 5.356033, 5.453192, 5.513427, 
    5.51753, 5.549628, 5.688647, 5.683352, 5.618227, 5.4899, 5.309708, 
    5.098572, 4.885837, 4.704521, 4.580997, 4.524658, 4.537004, 4.608436, 
    4.726605, 4.870749, 5.021959, 5.17297, 5.319542, 5.456137, 5.576294, 
    5.671569, 5.731426, 5.744835, 5.704313, 5.611754, 5.482604, 5.343098, 
    5.219526, 5.12711, 5.067253, 5.032856, 5.014951, 5.00638, 5.002567, 
    5.000986,
  // momentumX(4,32, 0-49)
    5.000058, 5.000175, 5.000499, 5.001343, 5.003422, 5.008226, 5.018595, 
    5.039321, 5.077241, 5.13961, 5.229686, 5.340741, 5.453701, 5.542929, 
    5.586711, 5.634364, 5.810377, 5.794869, 5.715106, 5.578702, 5.402011, 
    5.211908, 5.024439, 4.868459, 4.765963, 4.722025, 4.737376, 4.804413, 
    4.91415, 5.046367, 5.181589, 5.319583, 5.449525, 5.565306, 5.65952, 
    5.722928, 5.745382, 5.718771, 5.641876, 5.524932, 5.389545, 5.261234, 
    5.158674, 5.08793, 5.04487, 5.021269, 5.009429, 5.003929, 5.001545, 
    5.000584,
  // momentumX(4,33, 0-49)
    5.00004, 5.000121, 5.000348, 5.000955, 5.002475, 5.006059, 5.013967, 
    5.030193, 5.060858, 5.113483, 5.193935, 5.30105, 5.422253, 5.535433, 
    5.617548, 5.69124, 5.875936, 5.864213, 5.786301, 5.657351, 5.496267, 
    5.333714, 5.17509, 5.044634, 4.961142, 4.927159, 4.943112, 5.003295, 
    5.101369, 5.218139, 5.334802, 5.456174, 5.565315, 5.655402, 5.718253, 
    5.744672, 5.726639, 5.661288, 5.555245, 5.425946, 5.296785, 5.187774, 
    5.108407, 5.057558, 5.028332, 5.01302, 5.005613, 5.00228, 5.000876, 
    5.000325,
  // momentumX(4,34, 0-49)
    5.000024, 5.000075, 5.000218, 5.000609, 5.001614, 5.004035, 5.009521, 
    5.021117, 5.043819, 5.084566, 5.150602, 5.245469, 5.363938, 5.490148, 
    5.602442, 5.704795, 5.886364, 5.892461, 5.832005, 5.724312, 5.588806, 
    5.458125, 5.330325, 5.225271, 5.159105, 5.133275, 5.148096, 5.1995, 
    5.282907, 5.380851, 5.476084, 5.576321, 5.659528, 5.718254, 5.744268, 
    5.730054, 5.672071, 5.574646, 5.451857, 5.324495, 5.212377, 5.12704, 
    5.069887, 5.035612, 5.016918, 5.007533, 5.003155, 5.001247, 5.000467, 
    5.000169,
  // momentumX(4,35, 0-49)
    5.000014, 5.000041, 5.000124, 5.000355, 5.000961, 5.002462, 5.00596, 
    5.013583, 5.029061, 5.058093, 5.107836, 5.184575, 5.289448, 5.414499, 
    5.54309, 5.668658, 5.844255, 5.878744, 5.849082, 5.774486, 5.672875, 
    5.577171, 5.48142, 5.401774, 5.351748, 5.332812, 5.345255, 5.386293, 
    5.452143, 5.527818, 5.598071, 5.671585, 5.722932, 5.744674, 5.730054, 
    5.67552, 5.58408, 5.467301, 5.343374, 5.230956, 5.142365, 5.080799, 
    5.04248, 5.020813, 5.009551, 5.004119, 5.001675, 5.000645, 5.000236, 
    5.000084,
  // momentumX(4,36, 0-49)
    5.000007, 5.000022, 5.000065, 5.00019, 5.000528, 5.001387, 5.003449, 
    5.008088, 5.01785, 5.036942, 5.071377, 5.128031, 5.211954, 5.322424, 
    5.450345, 5.586574, 5.754741, 5.821698, 5.831575, 5.79887, 5.73787, 
    5.679853, 5.617424, 5.563701, 5.529284, 5.51648, 5.525597, 5.554762, 
    5.600111, 5.649807, 5.69079, 5.731433, 5.745385, 5.72664, 5.672071, 
    5.58408, 5.472425, 5.352917, 5.242486, 5.153233, 5.089346, 5.048308, 
    5.024346, 5.011489, 5.005095, 5.002128, 5.00084, 5.000314, 5.000111, 
    5.000039,
  // momentumX(4,37, 0-49)
    5.000002, 5.000011, 5.000032, 5.000094, 5.00027, 5.000727, 5.001855, 
    5.004479, 5.010196, 5.021828, 5.043808, 5.082083, 5.142909, 5.230166, 
    5.342067, 5.472644, 5.628459, 5.722989, 5.773468, 5.786318, 5.77012, 
    5.752038, 5.724462, 5.697757, 5.679138, 5.672138, 5.677126, 5.692811, 
    5.714684, 5.734652, 5.742105, 5.744839, 5.718772, 5.661288, 5.574646, 
    5.467301, 5.352917, 5.246391, 5.158862, 5.094786, 5.052536, 5.027167, 
    5.013159, 5.00599, 5.002568, 5.001039, 5.000397, 5.000144, 5.00005, 
    5.000018,
  // momentumX(4,38, 0-49)
    5, 5.000005, 5.000015, 5.000044, 5.000129, 5.000355, 5.000931, 5.002315, 
    5.005435, 5.012023, 5.025013, 5.048794, 5.088931, 5.150884, 5.237588, 
    5.348084, 5.483159, 5.591568, 5.673834, 5.728097, 5.756079, 5.778114, 
    5.786222, 5.787565, 5.785347, 5.784119, 5.784297, 5.784952, 5.780969, 
    5.768591, 5.740396, 5.704315, 5.641877, 5.555245, 5.451857, 5.343374, 
    5.242486, 5.158862, 5.096653, 5.05476, 5.028989, 5.014386, 5.006711, 
    5.002948, 5.001224, 5.00048, 5.000178, 5.000063, 5.000022, 5.000008,
  // momentumX(4,39, 0-49)
    5, 5.000001, 5.000007, 5.00002, 5.000057, 5.000163, 5.000438, 5.00112, 
    5.002711, 5.006193, 5.013331, 5.026992, 5.051274, 5.091135, 5.151162, 
    5.233976, 5.340683, 5.445152, 5.541938, 5.624341, 5.688284, 5.745618, 
    5.787155, 5.815814, 5.830077, 5.834549, 5.829556, 5.814503, 5.784487, 
    5.740712, 5.680091, 5.611754, 5.524933, 5.425946, 5.324495, 5.230956, 
    5.153233, 5.094786, 5.05476, 5.029618, 5.015037, 5.00718, 5.003231, 
    5.001372, 5.00055, 5.00021, 5.000076, 5.000027, 5.00001, 5.000003,
  // momentumX(4,40, 0-49)
    5, 5, 5.000002, 5.000009, 5.000025, 5.00007, 5.000193, 5.000509, 
    5.001269, 5.002991, 5.006652, 5.013947, 5.027512, 5.050968, 5.088504, 
    5.143935, 5.219826, 5.305856, 5.397701, 5.488678, 5.572298, 5.652788, 
    5.719582, 5.770612, 5.799332, 5.808841, 5.799087, 5.769994, 5.718313, 
    5.650439, 5.568352, 5.482605, 5.389545, 5.296785, 5.212377, 5.142365, 
    5.089346, 5.052536, 5.028989, 5.015037, 5.007341, 5.00338, 5.001469, 
    5.000603, 5.000236, 5.000087, 5.000031, 5.000011, 5.000004, 5,
  // momentumX(4,41, 0-49)
    5, 5, 5, 5.000003, 5.000011, 5.000029, 5.000081, 5.000217, 5.000558, 
    5.001357, 5.003117, 5.006752, 5.013795, 5.026531, 5.047973, 5.081492, 
    5.130116, 5.191607, 5.264742, 5.345742, 5.429265, 5.515083, 5.592558, 
    5.655453, 5.693151, 5.705927, 5.693044, 5.655183, 5.592001, 5.51405, 
    5.427535, 5.343099, 5.261235, 5.187774, 5.12704, 5.080799, 5.048308, 
    5.027167, 5.014386, 5.00718, 5.00338, 5.001504, 5.000631, 5.00025, 
    5.000094, 5.000034, 5.000013, 5.000005, 5, 5,
  // momentumX(4,42, 0-49)
    5, 5, 5, 5, 5.000005, 5.000012, 5.000032, 5.000088, 5.000232, 5.00058, 
    5.001373, 5.003073, 5.006487, 5.012912, 5.024214, 5.042749, 5.071041, 
    5.10987, 5.16003, 5.220561, 5.28869, 5.362971, 5.434639, 5.495757, 
    5.534231, 5.547513, 5.534188, 5.495649, 5.434417, 5.36256, 5.288007, 
    5.219526, 5.158674, 5.108407, 5.069887, 5.04248, 5.024346, 5.013159, 
    5.006711, 5.003231, 5.001469, 5.000631, 5.000257, 5.000099, 5.000036, 
    5.000014, 5.000005, 5.000001, 5, 5,
  // momentumX(4,43, 0-49)
    5, 5, 5, 5, 5.000001, 5.000005, 5.000013, 5.000034, 5.000092, 5.000234, 
    5.000571, 5.001317, 5.002868, 5.005898, 5.011437, 5.020907, 5.036011, 
    5.058069, 5.088407, 5.127475, 5.17446, 5.228262, 5.28295, 5.331479, 
    5.36327, 5.374421, 5.363255, 5.331441, 5.28287, 5.228115, 5.174216, 
    5.12711, 5.08793, 5.057558, 5.035612, 5.020813, 5.011489, 5.00599, 
    5.002948, 5.001372, 5.000603, 5.00025, 5.000099, 5.000037, 5.000015, 
    5.000006, 5.000001, 5, 5, 5,
  // momentumX(4,44, 0-49)
    5, 5, 5, 5, 5, 5.000001, 5.000006, 5.000014, 5.000034, 5.00009, 5.000225, 
    5.000533, 5.001195, 5.002535, 5.005076, 5.009581, 5.017048, 5.028498, 
    5.045024, 5.067372, 5.095585, 5.129107, 5.164498, 5.196819, 5.218636, 
    5.226383, 5.218631, 5.196807, 5.164472, 5.12906, 5.095506, 5.067253, 
    5.044869, 5.028332, 5.016918, 5.009551, 5.005095, 5.002568, 5.001224, 
    5.00055, 5.000236, 5.000094, 5.000036, 5.000015, 5.000007, 5.000002, 5, 
    5, 5, 5,
  // momentumX(4,45, 0-49)
    5, 5, 5, 5, 5, 5, 5.000002, 5.000006, 5.000013, 5.000032, 5.000083, 
    5.000204, 5.000471, 5.001028, 5.002122, 5.004128, 5.007573, 5.013069, 
    5.021315, 5.032892, 5.048037, 5.066514, 5.086528, 5.105148, 5.117975, 
    5.122566, 5.117973, 5.105145, 5.086521, 5.0665, 5.048013, 5.032856, 
    5.021268, 5.013019, 5.007533, 5.004119, 5.002128, 5.001039, 5.00048, 
    5.00021, 5.000087, 5.000034, 5.000014, 5.000006, 5.000002, 5, 5, 5, 5, 5,
  // momentumX(4,46, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000005, 5.000012, 5.00003, 5.000074, 
    5.000175, 5.000395, 5.000838, 5.001678, 5.003167, 5.005628, 5.009441, 
    5.01496, 5.022381, 5.031613, 5.041788, 5.051359, 5.058036, 5.060439, 
    5.058036, 5.051358, 5.041786, 5.03161, 5.022376, 5.014949, 5.009427, 
    5.005613, 5.003155, 5.001675, 5.00084, 5.000397, 5.000178, 5.000076, 
    5.000031, 5.000013, 5.000005, 5.000001, 5, 5, 5, 5, 5, 5,
  // momentumX(4,47, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000005, 5.000011, 5.000026, 5.000062, 
    5.000143, 5.000313, 5.000644, 5.001248, 5.002281, 5.003928, 5.006376, 
    5.009744, 5.014003, 5.018755, 5.023259, 5.026426, 5.027568, 5.026426, 
    5.023259, 5.018755, 5.014002, 5.009743, 5.006373, 5.003924, 5.002277, 
    5.001245, 5.000643, 5.000314, 5.000143, 5.000063, 5.000027, 5.000011, 
    5.000005, 5.000001, 5, 5, 5, 5, 5, 5, 5,
  // momentumX(4,48, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000004, 5.00001, 5.000022, 5.000049, 
    5.000109, 5.000232, 5.000462, 5.000867, 5.001534, 5.002549, 5.003979, 
    5.005815, 5.007891, 5.009873, 5.011274, 5.01178, 5.011274, 5.009873, 
    5.007891, 5.005815, 5.003978, 5.002548, 5.001532, 5.000866, 5.000462, 
    5.000232, 5.000109, 5.000049, 5.000022, 5.00001, 5.000004, 5, 5, 5, 5, 5, 
    5, 5, 5, 5,
  // momentumX(4,49, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000005, 5.000012, 5.00003, 
    5.000065, 5.000139, 5.000275, 5.000512, 5.000896, 5.001465, 5.002233, 
    5.00314, 5.004033, 5.004668, 5.004897, 5.004668, 5.004033, 5.00314, 
    5.002233, 5.001465, 5.000896, 5.000512, 5.000275, 5.000139, 5.000065, 
    5.00003, 5.000012, 5.000005, 5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumX(5,0, 0-49)
    5, 5, 5, 5, 5, 5, 5.000002, 5.000006, 5.000013, 5.000028, 5.000061, 
    5.00013, 5.000265, 5.000516, 5.00096, 5.001699, 5.002862, 5.004584, 
    5.006996, 5.010178, 5.014109, 5.018611, 5.023259, 5.027408, 5.030265, 
    5.031285, 5.030264, 5.027405, 5.023253, 5.018603, 5.014096, 5.010162, 
    5.006977, 5.004565, 5.002849, 5.001694, 5.000961, 5.00052, 5.000268, 
    5.000132, 5.000062, 5.000028, 5.000013, 5.000006, 5.000002, 5, 5, 5, 5, 5,
  // momentumX(5,1, 0-49)
    5, 5, 5, 5, 5, 5.000004, 5.000008, 5.000015, 5.000031, 5.000068, 
    5.000149, 5.000312, 5.000626, 5.0012, 5.002189, 5.003802, 5.006291, 
    5.0099, 5.01486, 5.021302, 5.029162, 5.038113, 5.047316, 5.055529, 
    5.06116, 5.063167, 5.061155, 5.05552, 5.047298, 5.038086, 5.029122, 
    5.021251, 5.0148, 5.00984, 5.006246, 5.003785, 5.002189, 5.001209, 
    5.000637, 5.00032, 5.000154, 5.000071, 5.000032, 5.000015, 5.000008, 
    5.000004, 5, 5, 5, 5,
  // momentumX(5,2, 0-49)
    5, 5, 5, 5, 5.000005, 5.000009, 5.000016, 5.000033, 5.000074, 5.000168, 
    5.000363, 5.000746, 5.001466, 5.00274, 5.004883, 5.00829, 5.013408, 
    5.020618, 5.030261, 5.042474, 5.057049, 5.073393, 5.08998, 5.104668, 
    5.114639, 5.118178, 5.114626, 5.10464, 5.089929, 5.07331, 5.056931, 
    5.042319, 5.030082, 5.020443, 5.013276, 5.008237, 5.00488, 5.002761, 
    5.001492, 5.000769, 5.000379, 5.000178, 5.000082, 5.000035, 5.000017, 
    5.000009, 5.000005, 5.000001, 5, 5,
  // momentumX(5,3, 0-49)
    5, 5, 5, 5.000004, 5.000009, 5.000016, 5.000034, 5.000081, 5.000184, 
    5.000405, 5.000853, 5.001713, 5.00328, 5.005985, 5.010404, 5.017234, 
    5.027194, 5.040734, 5.058229, 5.079662, 5.104465, 5.131642, 5.158663, 
    5.182254, 5.198014, 5.203566, 5.197978, 5.182171, 5.158515, 5.131409, 
    5.104133, 5.079228, 5.057729, 5.040246, 5.026826, 5.017087, 5.010396, 
    5.006039, 5.00335, 5.001772, 5.000896, 5.000432, 5.000201, 5.000089, 
    5.000038, 5.000018, 5.00001, 5.000006, 5.000001, 5,
  // momentumX(5,4, 0-49)
    5, 5, 5.000002, 5.000008, 5.000016, 5.000034, 5.000082, 5.000193, 
    5.000432, 5.000931, 5.001913, 5.003746, 5.006992, 5.012434, 5.021055, 
    5.033954, 5.052146, 5.075799, 5.105033, 5.139303, 5.177319, 5.217662, 
    5.25659, 5.289864, 5.311574, 5.319134, 5.311477, 5.289647, 5.256206, 
    5.217056, 5.176451, 5.13817, 5.103726, 5.074522, 5.051179, 5.033571, 
    5.021023, 5.012565, 5.007167, 5.003901, 5.002026, 5.001004, 5.000476, 
    5.000216, 5.000093, 5.00004, 5.000018, 5.00001, 5.000005, 5,
  // momentumX(5,5, 0-49)
    5, 5.000001, 5.000006, 5.000015, 5.000033, 5.000081, 5.000193, 5.000442, 
    5.000971, 5.002039, 5.004083, 5.00779, 5.014157, 5.024488, 5.040304, 
    5.063102, 5.094024, 5.131987, 5.176251, 5.225178, 5.276432, 5.328592, 
    5.376917, 5.417064, 5.442416, 5.451099, 5.442188, 5.416547, 5.376002, 
    5.32715, 5.274362, 5.222458, 5.173093, 5.128881, 5.09165, 5.062176, 
    5.040218, 5.024799, 5.014578, 5.008171, 5.004367, 5.002228, 5.001084, 
    5.000504, 5.000224, 5.000095, 5.00004, 5.000018, 5.000009, 5.000004,
  // momentumX(5,6, 0-49)
    5.000001, 5.000005, 5.000013, 5.000031, 5.000074, 5.000183, 5.00043, 
    5.000967, 5.002075, 5.004246, 5.008282, 5.015374, 5.02715, 5.045572, 
    5.072659, 5.110019, 5.15846, 5.213607, 5.273174, 5.334088, 5.393208, 
    5.450352, 5.500582, 5.540859, 5.565177, 5.573293, 5.564681, 5.539737, 
    5.498604, 5.447233, 5.388718, 5.328151, 5.266213, 5.206674, 5.153087, 
    5.107989, 5.072482, 5.046282, 5.028121, 5.016266, 5.008961, 5.004705, 
    5.002356, 5.001125, 5.000514, 5.000224, 5.000093, 5.000038, 5.000018, 
    5.000008,
  // momentumX(5,7, 0-49)
    5.000004, 5.00001, 5.000028, 5.000067, 5.000166, 5.0004, 5.000918, 
    5.002015, 5.004214, 5.008401, 5.015932, 5.02872, 5.04916, 5.079797, 
    5.122718, 5.178854, 5.248075, 5.319426, 5.389174, 5.453479, 5.509659, 
    5.560696, 5.602446, 5.634424, 5.65239, 5.658066, 5.651396, 5.632189, 
    5.598525, 5.554535, 5.500804, 5.441733, 5.375283, 5.305392, 5.237004, 
    5.174875, 5.122472, 5.081369, 5.051301, 5.030718, 5.017484, 5.009469, 
    5.004883, 5.002399, 5.001125, 5.000504, 5.000216, 5.000089, 5.000036, 
    5.000016,
  // momentumX(5,8, 0-49)
    5.000009, 5.000022, 5.000058, 5.000145, 5.000354, 5.000831, 5.001863, 
    5.003988, 5.008126, 5.015749, 5.028997, 5.050632, 5.083705, 5.130813, 
    5.193053, 5.269456, 5.35902, 5.440007, 5.509358, 5.56441, 5.604834, 
    5.638444, 5.662354, 5.67907, 5.686673, 5.688493, 5.684813, 5.674917, 
    5.655134, 5.627209, 5.588828, 5.543271, 5.484299, 5.414421, 5.338465, 
    5.262632, 5.193025, 5.134175, 5.088205, 5.054886, 5.03237, 5.018123, 
    5.009644, 5.004883, 5.002356, 5.001084, 5.000476, 5.000201, 5.000082, 
    5.000034,
  // momentumX(5,9, 0-49)
    5.000019, 5.000048, 5.00012, 5.000298, 5.000716, 5.001643, 5.003593, 
    5.007489, 5.014842, 5.027926, 5.049793, 5.083932, 5.133445, 5.199761, 
    5.281408, 5.374544, 5.47942, 5.558947, 5.615193, 5.648915, 5.663444, 
    5.671911, 5.672351, 5.669973, 5.665254, 5.662431, 5.661954, 5.662679, 
    5.659845, 5.652761, 5.636622, 5.613993, 5.574114, 5.516903, 5.445178, 
    5.364569, 5.282547, 5.20661, 5.142382, 5.092508, 5.056751, 5.032938, 
    5.018123, 5.009469, 5.004705, 5.002228, 5.001004, 5.000433, 5.00018, 
    5.000075,
  // momentumX(5,10, 0-49)
    5.000036, 5.000093, 5.000239, 5.000585, 5.001373, 5.003076, 5.006561, 
    5.013308, 5.02562, 5.046711, 5.08042, 5.130344, 5.198357, 5.283011, 
    5.378876, 5.479668, 5.591911, 5.658225, 5.691349, 5.696425, 5.68037, 
    5.66087, 5.636159, 5.613672, 5.596256, 5.58842, 5.590661, 5.601462, 
    5.615591, 5.630049, 5.638243, 5.642887, 5.629557, 5.59555, 5.540604, 
    5.467718, 5.383308, 5.296116, 5.215004, 5.146606, 5.093976, 5.056751, 
    5.03237, 5.017484, 5.008961, 5.004367, 5.002027, 5.000896, 5.000381, 
    5.000162,
  // momentumX(5,11, 0-49)
    5.000071, 5.000181, 5.000453, 5.001088, 5.002494, 5.005449, 5.011323, 
    5.022336, 5.041712, 5.073508, 5.121789, 5.189017, 5.274099, 5.371275, 
    5.471056, 5.567159, 5.679311, 5.724144, 5.729917, 5.705225, 5.659316, 
    5.612999, 5.564149, 5.522204, 5.492456, 5.479336, 5.483345, 5.502607, 
    5.531834, 5.56584, 5.596796, 5.628322, 5.64375, 5.638568, 5.609673, 
    5.556548, 5.482425, 5.39456, 5.302978, 5.217842, 5.146606, 5.092508, 
    5.054886, 5.030718, 5.016266, 5.008171, 5.003901, 5.001774, 5.000774, 
    5.000335,
  // momentumX(5,12, 0-49)
    5.000131, 5.00033, 5.000812, 5.001908, 5.004274, 5.00911, 5.018438, 
    5.035336, 5.0639, 5.108568, 5.172517, 5.255433, 5.351807, 5.45142, 
    5.54234, 5.622025, 5.729712, 5.750149, 5.730207, 5.67971, 5.608513, 
    5.538956, 5.468381, 5.40834, 5.366759, 5.347938, 5.352461, 5.37809, 
    5.419709, 5.470071, 5.520361, 5.575464, 5.617815, 5.642097, 5.643387, 
    5.618141, 5.565696, 5.48967, 5.398307, 5.302978, 5.215004, 5.142382, 
    5.088205, 5.051301, 5.028121, 5.014579, 5.007169, 5.003353, 5.001502, 
    5.000663,
  // momentumX(5,13, 0-49)
    5.000229, 5.000569, 5.001369, 5.00315, 5.006894, 5.014339, 5.02826, 
    5.052577, 5.091915, 5.1502, 5.228284, 5.321659, 5.420121, 5.510469, 
    5.580884, 5.636158, 5.738116, 5.735927, 5.695858, 5.626519, 5.536742, 
    5.448798, 5.359662, 5.283228, 5.230228, 5.205044, 5.208557, 5.238231, 
    5.289241, 5.352497, 5.418259, 5.492509, 5.55786, 5.608896, 5.639956, 
    5.645646, 5.622089, 5.568675, 5.48967, 5.39456, 5.296116, 5.20661, 
    5.134175, 5.081369, 5.046282, 5.0248, 5.012568, 5.006046, 5.00278, 
    5.001256,
  // momentumX(5,14, 0-49)
    5.000374, 5.000917, 5.002163, 5.004873, 5.010436, 5.021191, 5.040668, 
    5.073408, 5.123923, 5.194474, 5.282308, 5.378265, 5.468612, 5.539557, 
    5.581494, 5.609149, 5.704862, 5.684734, 5.631863, 5.551764, 5.45104, 
    5.350298, 5.246478, 5.15581, 5.091814, 5.059381, 5.060057, 5.091223, 
    5.148467, 5.22124, 5.298869, 5.387869, 5.471773, 5.545377, 5.60301, 
    5.638582, 5.646293, 5.622088, 5.565695, 5.482424, 5.383307, 5.282547, 
    5.193025, 5.122472, 5.072483, 5.040219, 5.021027, 5.010407, 5.004912, 
    5.002266,
  // momentumX(5,15, 0-49)
    5.000567, 5.001374, 5.003187, 5.00704, 5.014763, 5.029299, 5.054786, 
    5.09597, 5.156433, 5.235746, 5.326997, 5.417121, 5.49086, 5.535902, 
    5.545708, 5.546775, 5.632914, 5.60088, 5.542744, 5.459904, 5.356049, 
    5.248635, 5.134977, 5.033073, 4.95883, 4.918158, 4.913803, 4.943549, 
    5.003622, 5.082602, 5.168946, 5.268797, 5.367137, 5.458964, 5.538911, 
    5.600954, 5.638575, 5.645641, 5.618137, 5.556546, 5.467716, 5.364568, 
    5.262632, 5.174875, 5.10799, 5.062179, 5.033578, 5.017106, 5.008286, 
    5.003901,
  // momentumX(5,16, 0-49)
    5.000793, 5.001904, 5.004345, 5.009432, 5.01941, 5.037717, 5.06884, 
    5.117216, 5.184804, 5.268004, 5.356136, 5.433732, 5.48586, 5.502688, 
    5.480472, 5.459173, 5.525829, 5.488203, 5.431913, 5.353796, 5.254422, 
    5.146871, 5.029435, 4.92056, 4.837578, 4.787774, 4.775797, 4.80067, 
    4.859735, 4.941498, 5.033751, 5.14112, 5.250391, 5.356567, 5.454606, 
    5.538887, 5.602984, 5.639937, 5.643376, 5.609665, 5.5406, 5.445177, 
    5.338465, 5.237003, 5.153089, 5.091654, 5.05119, 5.026856, 5.013346, 
    5.006411,
  // momentumX(5,17, 0-49)
    5.001009, 5.002405, 5.005424, 5.01161, 5.023516, 5.044888, 5.080247, 
    5.133332, 5.204224, 5.28643, 5.36658, 5.428285, 5.457914, 5.448078, 
    5.397178, 5.359798, 5.38727, 5.349489, 5.301646, 5.235264, 5.147697, 
    5.046798, 4.932895, 4.822896, 4.733915, 4.674499, 4.651908, 4.667727, 
    4.721311, 4.802092, 4.897588, 5.009571, 5.126815, 5.244068, 5.35647, 
    5.458864, 5.5453, 5.608845, 5.642067, 5.638551, 5.595541, 5.5169, 
    5.414419, 5.305392, 5.206675, 5.128885, 5.074537, 5.040285, 5.020535, 
    5.010053,
  // momentumX(5,18, 0-49)
    5.001149, 5.002726, 5.006095, 5.012916, 5.025878, 5.048788, 5.085967, 
    5.140407, 5.210714, 5.288495, 5.358942, 5.405567, 5.415976, 5.384698, 
    5.312162, 5.264491, 5.221843, 5.186554, 5.153127, 5.1055, 5.037116, 
    4.949855, 4.847899, 4.744311, 4.653742, 4.585035, 4.548517, 4.550172, 
    4.592954, 4.668444, 4.76445, 4.87837, 5.000965, 5.126472, 5.250022, 
    5.366846, 5.471569, 5.55773, 5.617738, 5.643708, 5.629535, 5.574101, 
    5.484294, 5.375281, 5.266214, 5.1731, 5.103745, 5.057774, 5.03019, 
    5.015046,
  // momentumX(5,19, 0-49)
    5.001132, 5.00268, 5.005971, 5.012604, 5.025155, 5.04725, 5.082956, 
    5.134978, 5.201641, 5.274235, 5.337543, 5.374701, 5.373543, 5.330182, 
    5.248117, 5.187968, 5.03577, 5.00039, 4.986063, 4.964749, 4.923753, 
    4.857672, 4.777114, 4.68915, 4.603427, 4.527005, 4.473067, 4.454343, 
    4.479911, 4.545097, 4.638662, 4.751842, 4.87722, 5.008308, 5.14009, 
    5.268059, 5.38738, 5.492204, 5.575282, 5.62822, 5.642832, 5.613966, 
    5.543258, 5.441728, 5.32815, 5.222465, 5.138189, 5.079276, 5.042429, 
    5.021496,
  // momentumX(5,20, 0-49)
    5.000885, 5.002056, 5.004517, 5.009397, 5.018436, 5.033949, 5.05833, 
    5.092862, 5.13604, 5.182454, 5.22361, 5.251111, 5.26051, 5.253445, 
    5.236856, 0, 4.882641, 4.890296, 4.897371, 4.893323, 4.87047, 4.819962, 
    4.758723, 4.686413, 4.605082, 4.517176, 4.437809, 4.388928, 4.388727, 
    4.437592, 4.525457, 4.634996, 4.760348, 4.894176, 5.031245, 5.167237, 
    5.297763, 5.417573, 5.519956, 5.596563, 5.638118, 5.636558, 5.588799, 
    5.500793, 5.388714, 5.274365, 5.176466, 5.104169, 5.057017, 5.029309,
  // momentumX(5,21, 0-49)
    5.000641, 5.001482, 5.003266, 5.006831, 5.013499, 5.025104, 5.043731, 
    5.070997, 5.106867, 5.148563, 5.190476, 5.225755, 5.249031, 5.258772, 
    5.257997, 0, 4.74108, 4.76133, 4.784954, 4.801523, 4.801844, 4.771854, 
    4.732392, 4.676557, 4.600542, 4.503641, 4.402691, 4.328095, 4.306149, 
    4.341571, 4.42612, 4.532413, 4.657756, 4.794104, 4.93592, 5.078889, 
    5.218863, 5.351027, 5.469194, 5.565336, 5.629769, 5.652613, 5.627135, 
    5.554501, 5.447219, 5.327146, 5.217059, 5.131421, 5.073335, 5.038131,
  // momentumX(5,22, 0-49)
    5.000444, 5.00103, 5.002293, 5.004852, 5.009718, 5.018359, 5.0326, 
    5.054197, 5.084013, 5.121048, 5.161894, 5.201262, 5.233709, 5.255754, 
    5.267343, 0, 4.627163, 4.653697, 4.689208, 4.723159, 4.745467, 4.737381, 
    4.725026, 4.694858, 4.635277, 4.538174, 4.417841, 4.312981, 4.261384, 
    4.275565, 4.351222, 4.44836, 4.569024, 4.704297, 4.848145, 4.995989, 
    5.143591, 5.286217, 5.41789, 5.530775, 5.614996, 5.659525, 5.65497, 
    5.598444, 5.498568, 5.375984, 5.256189, 5.158487, 5.089858, 5.047126,
  // momentumX(5,23, 0-49)
    5.000326, 5.000756, 5.0017, 5.003643, 5.007394, 5.014186, 5.025643, 
    5.043532, 5.069174, 5.102598, 5.141809, 5.182737, 5.220225, 5.249777, 
    5.26927, 0, 4.542715, 4.572813, 4.616893, 4.664588, 4.705509, 4.716725, 
    4.729808, 4.725214, 4.68426, 4.591591, 4.457345, 4.326142, 4.246144, 
    4.238336, 4.303779, 4.389193, 4.502711, 4.634574, 4.778222, 4.928749, 
    5.081713, 5.232281, 5.374473, 5.500473, 5.600245, 5.662012, 5.674566, 
    5.632014, 5.539653, 5.416502, 5.289604, 5.182093, 5.104459, 5.055098,
  // momentumX(5,24, 0-49)
    5.000295, 5.00068, 5.00153, 5.00328, 5.006674, 5.012842, 5.023315, 
    5.039814, 5.063758, 5.095514, 5.133634, 5.174624, 5.213623, 5.245886, 
    5.268474, 0, 4.488168, 4.520331, 4.569875, 4.626774, 4.680708, 4.705749, 
    4.737486, 4.751808, 4.725004, 4.637198, 4.495549, 4.347715, 4.248083, 
    4.223984, 4.28151, 4.357102, 4.464386, 4.592849, 4.73542, 4.886861, 
    5.042512, 5.19742, 5.345583, 5.479222, 5.588269, 5.660618, 5.684098, 
    5.651032, 5.564503, 5.442098, 5.311407, 5.19786, 5.114362, 5.060548,
  // momentumX(5,25, 0-49)
    5.000359, 5.000815, 5.001808, 5.003817, 5.007643, 5.014476, 5.025854, 
    5.043424, 5.068394, 5.100799, 5.138853, 5.178908, 5.216267, 5.246636, 
    5.267615, 0, 4.464517, 4.497284, 4.548565, 4.608568, 4.667108, 4.6971, 
    4.73595, 4.757792, 4.737058, 4.652288, 4.509429, 4.356791, 4.250607, 
    4.22062, 4.27515, 4.34684, 4.451613, 4.57867, 4.72073, 4.872409, 
    5.028946, 5.185324, 5.335518, 5.471749, 5.583937, 5.659878, 5.6871, 
    5.657343, 5.572935, 5.450924, 5.319024, 5.203423, 5.117879, 5.062491,
  // momentumX(5,26, 0-49)
    5.000526, 5.001181, 5.002566, 5.005302, 5.010374, 5.01916, 5.033297, 
    5.054275, 5.082738, 5.117734, 5.156352, 5.194211, 5.226768, 5.250868, 
    5.265858, 0, 4.47485, 4.506453, 4.555189, 4.611245, 4.664432, 4.688535, 
    4.720223, 4.735377, 4.710451, 4.625587, 4.487513, 4.343034, 4.245784, 
    4.222999, 4.281123, 4.356955, 4.46433, 4.592826, 4.735413, 4.886859, 
    5.042512, 5.19742, 5.345583, 5.479222, 5.588269, 5.660618, 5.684098, 
    5.651031, 5.564503, 5.442098, 5.311407, 5.19786, 5.114362, 5.060548,
  // momentumX(5,27, 0-49)
    5.000805, 5.001794, 5.003833, 5.007775, 5.014898, 5.026875, 5.045452, 
    5.071789, 5.105519, 5.144054, 5.182762, 5.21631, 5.240609, 5.254356, 
    5.259472, 0, 4.523546, 4.551486, 4.592946, 4.637959, 4.676403, 4.684864, 
    4.697034, 4.693454, 4.655822, 4.568797, 4.441556, 4.316923, 4.241585, 
    4.236356, 4.302987, 4.388885, 4.502593, 4.634529, 4.778204, 4.928742, 
    5.081711, 5.232281, 5.374472, 5.500473, 5.600244, 5.662012, 5.674566, 
    5.632014, 5.539653, 5.416502, 5.289604, 5.182093, 5.104459, 5.055098,
  // momentumX(5,28, 0-49)
    5.001189, 5.002643, 5.005589, 5.011191, 5.021119, 5.037401, 5.061837, 
    5.094956, 5.134828, 5.176611, 5.213614, 5.239749, 5.252041, 5.251792, 
    5.243953, 0, 4.61626, 4.63638, 4.665257, 4.692745, 4.709127, 4.695071, 
    4.679724, 4.649843, 4.594497, 4.505446, 4.395233, 4.299756, 4.254767, 
    4.27263, 4.350018, 4.447882, 4.568835, 4.704223, 4.848115, 4.995977, 
    5.143586, 5.286216, 5.417889, 5.530774, 5.614996, 5.659525, 5.65497, 
    5.598445, 5.498568, 5.375984, 5.256189, 5.158487, 5.089858, 5.047126,
  // momentumX(5,29, 0-49)
    5.001638, 5.003657, 5.007708, 5.01534, 5.02871, 5.05025, 5.081713, 
    5.122604, 5.168763, 5.212454, 5.244812, 5.259601, 5.255975, 5.238696, 
    5.215979, 0, 4.757369, 4.761571, 4.770969, 4.774717, 4.763777, 4.723468, 
    4.678093, 4.621346, 4.550265, 4.463518, 4.37518, 4.311992, 4.297986, 
    4.337866, 4.424553, 4.531772, 4.657499, 4.794, 4.935878, 5.078872, 
    5.218856, 5.351024, 5.469192, 5.565335, 5.629769, 5.652613, 5.627135, 
    5.554501, 5.447219, 5.327146, 5.217059, 5.131421, 5.073335, 5.038131,
  // momentumX(5,30, 0-49)
    5.002085, 5.004748, 5.010147, 5.020489, 5.03899, 5.069524, 5.115261, 
    5.176115, 5.24598, 5.31214, 5.358694, 5.372374, 5.346906, 5.283526, 
    5.188242, 5.105539, 4.913468, 4.864236, 4.846265, 4.829531, 4.79874, 
    4.743309, 4.680916, 4.612876, 4.541994, 4.469274, 4.40619, 4.370837, 
    4.379624, 4.433442, 4.523681, 4.634262, 4.760047, 4.894053, 5.031196, 
    5.167217, 5.297757, 5.417571, 5.519956, 5.596563, 5.638118, 5.636558, 
    5.588799, 5.500793, 5.388714, 5.274365, 5.176466, 5.104169, 5.057017, 
    5.029309,
  // momentumX(5,31, 0-49)
    5.002143, 5.004889, 5.010488, 5.021266, 5.040632, 5.072723, 5.12099, 
    5.185519, 5.260214, 5.332315, 5.385979, 5.407974, 5.391459, 5.335916, 
    5.244624, 5.177097, 5.096328, 5.048657, 5.011378, 4.966193, 4.904812, 
    4.824902, 4.735695, 4.645541, 4.563855, 4.495916, 4.451912, 4.441776, 
    4.473276, 4.541901, 4.637214, 4.751214, 4.876952, 5.008195, 5.140043, 
    5.268041, 5.387373, 5.492201, 5.575282, 5.62822, 5.642832, 5.613966, 
    5.543258, 5.441728, 5.328151, 5.222465, 5.138189, 5.079276, 5.042429, 
    5.021496,
  // momentumX(5,32, 0-49)
    5.001922, 5.004405, 5.009535, 5.019537, 5.037773, 5.068523, 5.115789, 
    5.180799, 5.258986, 5.338832, 5.40467, 5.442245, 5.443079, 5.405014, 
    5.329818, 5.271312, 5.264867, 5.214771, 5.161846, 5.095674, 5.012313, 
    4.915738, 4.80939, 4.706865, 4.621886, 4.561248, 4.53286, 4.540988, 
    4.588072, 4.666042, 4.76333, 4.877868, 5.000745, 5.126377, 5.249983, 
    5.366829, 5.471562, 5.557727, 5.617737, 5.643708, 5.629536, 5.574101, 
    5.484294, 5.375281, 5.266214, 5.1731, 5.103745, 5.057774, 5.03019, 
    5.015046,
  // momentumX(5,33, 0-49)
    5.00155, 5.003578, 5.007845, 5.01632, 5.032094, 5.059364, 5.102615, 
    5.16453, 5.242973, 5.328912, 5.40777, 5.464293, 5.487687, 5.473557, 
    5.422353, 5.376557, 5.412996, 5.361646, 5.298301, 5.217968, 5.119894, 
    5.013451, 4.898541, 4.791826, 4.709034, 4.656785, 4.640617, 4.661203, 
    4.717844, 4.800365, 4.89677, 5.009197, 5.126649, 5.243997, 5.35644, 
    5.458851, 5.545294, 5.608843, 5.642066, 5.638551, 5.595541, 5.5169, 
    5.414419, 5.305392, 5.206675, 5.128885, 5.074537, 5.040285, 5.020535, 
    5.010053,
  // momentumX(5,34, 0-49)
    5.001143, 5.002663, 5.005934, 5.012573, 5.025232, 5.04776, 5.084791, 
    5.14025, 5.21467, 5.302464, 5.391526, 5.466604, 5.514605, 5.528172, 
    5.505728, 5.478414, 5.53635, 5.487955, 5.419987, 5.331903, 5.225847, 
    5.115927, 5, 4.895658, 4.818719, 4.774924, 4.767848, 4.796153, 4.857343, 
    4.940302, 5.033179, 5.140856, 5.250273, 5.356515, 5.454584, 5.538877, 
    5.60298, 5.639935, 5.643376, 5.609665, 5.5406, 5.445177, 5.338465, 
    5.237003, 5.153089, 5.091654, 5.05119, 5.026856, 5.013346, 5.006411,
  // momentumX(5,35, 0-49)
    5.000779, 5.001836, 5.004165, 5.009008, 5.018488, 5.035882, 5.065555, 
    5.112102, 5.1783, 5.262308, 5.355819, 5.445318, 5.51646, 5.558745, 
    5.567586, 5.563785, 5.631766, 5.591699, 5.525231, 5.435889, 5.328604, 
    5.221323, 5.110783, 5.013813, 4.944966, 4.909076, 4.90834, 4.940494, 
    5.002017, 5.0818, 5.168562, 5.26862, 5.367057, 5.45893, 5.538898, 
    5.600948, 5.638573, 5.645639, 5.618137, 5.556546, 5.467717, 5.364568, 
    5.262632, 5.174875, 5.10799, 5.062179, 5.033578, 5.017106, 5.008286, 
    5.003901,
  // momentumX(5,36, 0-49)
    5.000493, 5.00118, 5.002732, 5.006036, 5.012685, 5.025267, 5.047535, 
    5.084073, 5.139023, 5.213765, 5.304395, 5.400975, 5.489923, 5.558537, 
    5.598734, 5.621789, 5.695973, 5.669862, 5.611474, 5.527821, 5.42626, 
    5.327377, 5.227425, 5.141449, 5.081936, 5.053137, 5.056394, 5.089209, 
    5.147419, 5.22072, 5.298621, 5.387753, 5.471721, 5.545353, 5.603, 
    5.638578, 5.646291, 5.622087, 5.565695, 5.482424, 5.383308, 5.282547, 
    5.193025, 5.122472, 5.072483, 5.040219, 5.021027, 5.010407, 5.004912, 
    5.002266,
  // momentumX(5,37, 0-49)
    5.000292, 5.00071, 5.00168, 5.003798, 5.008177, 5.016725, 5.032395, 
    5.059221, 5.101714, 5.163327, 5.244109, 5.338745, 5.436703, 5.525202, 
    5.5934, 5.644053, 5.725108, 5.718331, 5.675017, 5.604451, 5.51567, 
    5.430519, 5.345299, 5.272915, 5.223416, 5.200871, 5.206166, 5.236938, 
    5.288577, 5.352169, 5.418102, 5.492436, 5.557827, 5.608882, 5.639949, 
    5.645644, 5.622088, 5.568674, 5.489669, 5.39456, 5.296116, 5.20661, 
    5.134175, 5.081369, 5.046282, 5.0248, 5.012568, 5.006046, 5.00278, 
    5.001256,
  // momentumX(5,38, 0-49)
    5.000163, 5.000402, 5.000972, 5.002252, 5.004967, 5.01043, 5.02079, 
    5.039236, 5.069869, 5.116913, 5.18307, 5.267374, 5.363808, 5.462077, 
    5.550688, 5.62586, 5.715589, 5.73241, 5.710911, 5.660795, 5.591628, 
    5.525109, 5.458025, 5.401213, 5.362216, 5.345235, 5.350946, 5.377285, 
    5.419301, 5.469871, 5.520268, 5.57542, 5.617796, 5.642089, 5.643384, 
    5.61814, 5.565695, 5.489669, 5.398307, 5.302978, 5.215004, 5.142382, 
    5.088205, 5.051301, 5.028121, 5.014579, 5.007169, 5.003353, 5.001502, 
    5.000663,
  // momentumX(5,39, 0-49)
    5.000086, 5.000216, 5.000532, 5.00126, 5.002849, 5.006141, 5.012588, 
    5.024494, 5.045127, 5.078468, 5.128332, 5.196746, 5.282134, 5.37842, 
    5.476128, 5.568144, 5.666311, 5.708275, 5.713571, 5.690119, 5.646567, 
    5.603043, 5.557014, 5.517471, 5.489532, 5.477641, 5.482416, 5.502121, 
    5.53159, 5.565724, 5.596741, 5.628298, 5.64374, 5.638564, 5.60967, 
    5.556547, 5.482424, 5.39456, 5.302978, 5.217841, 5.146606, 5.092508, 
    5.054886, 5.030718, 5.016266, 5.008171, 5.003901, 5.001774, 5.000774, 
    5.000335,
  // momentumX(5,40, 0-49)
    5.000043, 5.00011, 5.000275, 5.000667, 5.001546, 5.00342, 5.007205, 
    5.014437, 5.02746, 5.049472, 5.084197, 5.134979, 5.203325, 5.287435, 
    5.381662, 5.479102, 5.581413, 5.64549, 5.67866, 5.685199, 5.671315, 
    5.65408, 5.631466, 5.610655, 5.594442, 5.587394, 5.59011, 5.601179, 
    5.615451, 5.629982, 5.638213, 5.642873, 5.629552, 5.595548, 5.540603, 
    5.467717, 5.383308, 5.296116, 5.215004, 5.146606, 5.093976, 5.056751, 
    5.03237, 5.017484, 5.008961, 5.004367, 5.002027, 5.000896, 5.000381, 
    5.000162,
  // momentumX(5,41, 0-49)
    5.000021, 5.000053, 5.000136, 5.000334, 5.000796, 5.001806, 5.003906, 
    5.008049, 5.015777, 5.029372, 5.051832, 5.086515, 5.136288, 5.202295, 
    5.282791, 5.373473, 5.471925, 5.54978, 5.606205, 5.641187, 5.657415, 
    5.667536, 5.669413, 5.668134, 5.664176, 5.661833, 5.66164, 5.662522, 
    5.65977, 5.652724, 5.636606, 5.613986, 5.57411, 5.516902, 5.445177, 
    5.364569, 5.282547, 5.20661, 5.142382, 5.092508, 5.056751, 5.032938, 
    5.018123, 5.009469, 5.004705, 5.002228, 5.001004, 5.000433, 5.00018, 
    5.000075,
  // momentumX(5,42, 0-49)
    5.00001, 5.000026, 5.000064, 5.00016, 5.000389, 5.000905, 5.002008, 
    5.004252, 5.008577, 5.016464, 5.030032, 5.051978, 5.08522, 5.132163, 
    5.193682, 5.268489, 5.354282, 5.43411, 5.503586, 5.559516, 5.601096, 
    5.635793, 5.660614, 5.678005, 5.686062, 5.688162, 5.684644, 5.674834, 
    5.655095, 5.62719, 5.588821, 5.543266, 5.484297, 5.41442, 5.338465, 
    5.262631, 5.193025, 5.134175, 5.088205, 5.054886, 5.03237, 5.018123, 
    5.009644, 5.004883, 5.002356, 5.001084, 5.000476, 5.000201, 5.000082, 
    5.000034,
  // momentumX(5,43, 0-49)
    5.000005, 5.000013, 5.00003, 5.000073, 5.000181, 5.000431, 5.000981, 
    5.002132, 5.00442, 5.008735, 5.016428, 5.029381, 5.049916, 5.080473, 
    5.122991, 5.178202, 5.245416, 5.316042, 5.385835, 5.450653, 5.507519, 
    5.559199, 5.60148, 5.633844, 5.652066, 5.657897, 5.651314, 5.632151, 
    5.598507, 5.554525, 5.500799, 5.441729, 5.37528, 5.30539, 5.237002, 
    5.174874, 5.122472, 5.081368, 5.051301, 5.030718, 5.017484, 5.009469, 
    5.004883, 5.002399, 5.001125, 5.000504, 5.000216, 5.000089, 5.000036, 
    5.000016,
  // momentumX(5,44, 0-49)
    5.000001, 5.000006, 5.000015, 5.000033, 5.000081, 5.000196, 5.000456, 
    5.001016, 5.002163, 5.004395, 5.008506, 5.01568, 5.027507, 5.045893, 
    5.072774, 5.109653, 5.157123, 5.211867, 5.271431, 5.332604, 5.392085, 
    5.449572, 5.500086, 5.540573, 5.56503, 5.573226, 5.564657, 5.539729, 
    5.498598, 5.447226, 5.38871, 5.328142, 5.266205, 5.206667, 5.153083, 
    5.107986, 5.07248, 5.046281, 5.028121, 5.016266, 5.008961, 5.004705, 
    5.002356, 5.001125, 5.000514, 5.000224, 5.000093, 5.000038, 5.000018, 
    5.000008,
  // momentumX(5,45, 0-49)
    5, 5.000002, 5.000007, 5.000016, 5.000035, 5.000085, 5.000203, 5.000461, 
    5.001007, 5.002101, 5.004179, 5.007924, 5.014315, 5.024631, 5.040349, 
    5.062917, 5.093406, 5.131166, 5.175416, 5.224458, 5.275883, 5.328215, 
    5.376691, 5.416956, 5.442389, 5.451115, 5.442218, 5.416569, 5.376009, 
    5.327141, 5.274342, 5.222435, 5.173072, 5.128863, 5.091638, 5.062168, 
    5.040212, 5.024796, 5.014577, 5.00817, 5.004367, 5.002228, 5.001084, 
    5.000504, 5.000224, 5.000095, 5.00004, 5.000018, 5.000009, 5.000004,
  // momentumX(5,46, 0-49)
    5, 5, 5.000003, 5.000008, 5.000017, 5.000037, 5.000086, 5.0002, 5.000446, 
    5.000955, 5.001951, 5.0038, 5.007055, 5.012488, 5.021063, 5.033856, 
    5.051858, 5.075415, 5.104631, 5.138946, 5.177042, 5.217485, 5.256517, 
    5.289888, 5.311668, 5.319259, 5.311596, 5.289727, 5.256232, 5.217037, 
    5.176403, 5.138111, 5.10367, 5.074477, 5.051146, 5.033548, 5.021009, 
    5.012557, 5.007162, 5.003898, 5.002025, 5.001004, 5.000476, 5.000216, 
    5.000093, 5.00004, 5.000018, 5.00001, 5.000005, 5,
  // momentumX(5,47, 0-49)
    5, 5, 5, 5.000004, 5.00001, 5.000017, 5.000035, 5.000082, 5.000188, 
    5.000413, 5.000865, 5.001729, 5.003295, 5.005988, 5.010376, 5.017145, 
    5.027009, 5.040486, 5.057955, 5.079401, 5.10426, 5.131539, 5.158699, 
    5.182441, 5.198313, 5.203908, 5.198285, 5.182379, 5.15859, 5.131369, 
    5.104017, 5.079085, 5.057591, 5.040131, 5.026741, 5.017027, 5.010357, 
    5.006016, 5.003337, 5.001766, 5.000893, 5.000431, 5.000199, 5.000088, 
    5.000038, 5.000018, 5.00001, 5.000006, 5.000001, 5,
  // momentumX(5,48, 0-49)
    5, 5, 5, 5, 5.000005, 5.000009, 5.000016, 5.000033, 5.000074, 5.000168, 
    5.00036, 5.000737, 5.001443, 5.002692, 5.004791, 5.008132, 5.013163, 
    5.020295, 5.029888, 5.0421, 5.056754, 5.073282, 5.09015, 5.105158, 
    5.115366, 5.118993, 5.115357, 5.105136, 5.090113, 5.073223, 5.056668, 
    5.041988, 5.029758, 5.020169, 5.013067, 5.00809, 5.004785, 5.002703, 
    5.001458, 5.00075, 5.000369, 5.000174, 5.000078, 5.000034, 5.000016, 
    5.000009, 5.000005, 5.000001, 5, 5,
  // momentumX(5,49, 0-49)
    5, 5, 5, 5, 5, 5.000002, 5.000004, 5.00001, 5.000021, 5.000049, 5.00011, 
    5.000237, 5.000488, 5.000957, 5.001791, 5.003193, 5.005428, 5.008776, 
    5.013537, 5.019944, 5.02806, 5.037715, 5.048037, 5.057581, 5.064183, 
    5.06655, 5.064181, 5.057576, 5.048025, 5.037696, 5.028031, 5.019907, 
    5.013492, 5.008731, 5.005393, 5.003181, 5.001791, 5.000962, 5.000493, 
    5.000242, 5.000113, 5.000051, 5.000022, 5.00001, 5.000005, 5.000002, 5, 
    5, 5, 5,
  // momentumX(6,0, 0-49)
    5.000001, 5.000006, 5.00001, 5.000018, 5.000034, 5.000072, 5.000154, 
    5.000316, 5.000631, 5.001208, 5.002222, 5.003925, 5.006657, 5.010836, 
    5.01693, 5.025394, 5.036568, 5.050474, 5.066961, 5.08557, 5.105506, 
    5.125745, 5.144631, 5.160282, 5.170508, 5.174044, 5.170405, 5.160065, 
    5.144283, 5.12525, 5.104868, 5.084815, 5.066161, 5.049734, 5.036002, 
    5.025083, 5.016811, 5.010836, 5.006715, 5.003999, 5.002289, 5.00126, 
    5.000666, 5.00034, 5.000166, 5.000079, 5.000038, 5.000019, 5.000011, 
    5.000007,
  // momentumX(6,1, 0-49)
    5.000005, 5.00001, 5.000018, 5.000033, 5.00007, 5.000151, 5.00032, 
    5.000653, 5.001278, 5.002406, 5.004348, 5.007544, 5.012561, 5.020073, 
    5.030783, 5.045307, 5.064008, 5.086517, 5.11232, 5.140503, 5.169809, 
    5.198979, 5.225753, 5.247741, 5.261885, 5.266718, 5.261647, 5.247239, 
    5.224946, 5.197832, 5.168324, 5.13874, 5.110439, 5.084771, 5.062673, 
    5.044592, 5.030516, 5.020079, 5.012699, 5.007718, 5.004508, 5.002532, 
    5.001365, 5.000708, 5.000353, 5.00017, 5.00008, 5.000038, 5.000021, 
    5.000012,
  // momentumX(6,2, 0-49)
    5.000009, 5.000016, 5.000031, 5.000069, 5.000152, 5.000327, 5.000679, 
    5.001356, 5.002598, 5.004784, 5.008452, 5.014331, 5.023312, 5.036367, 
    5.054408, 5.078065, 5.107471, 5.141197, 5.177971, 5.216177, 5.254053, 
    5.290477, 5.322897, 5.349, 5.365357, 5.37082, 5.364851, 5.347931, 
    5.321181, 5.288037, 5.250886, 5.212396, 5.173913, 5.137403, 5.104555, 
    5.076529, 5.053838, 5.036386, 5.023619, 5.014725, 5.008818, 5.005071, 
    5.002802, 5.001487, 5.000758, 5.000372, 5.000178, 5.000082, 5.000039, 
    5.000021,
  // momentumX(6,3, 0-49)
    5.000015, 5.000031, 5.000066, 5.000148, 5.000325, 5.000685, 5.001394, 
    5.002722, 5.005103, 5.009176, 5.015826, 5.026171, 5.041471, 5.06295, 
    5.091514, 5.127439, 5.170224, 5.216258, 5.26322, 5.308789, 5.351055, 
    5.389846, 5.422889, 5.44876, 5.464318, 5.469281, 5.463325, 5.446671, 
    5.41954, 5.385091, 5.344875, 5.301375, 5.2552, 5.208684, 5.164347, 
    5.124405, 5.090402, 5.063021, 5.042137, 5.027025, 5.016627, 5.009819, 
    5.005565, 5.003028, 5.001583, 5.000794, 5.000385, 5.00018, 5.000083, 
    5.00004,
  // momentumX(6,4, 0-49)
    5.000029, 5.000062, 5.00014, 5.00031, 5.000668, 5.001381, 5.002748, 
    5.005244, 5.009598, 5.016839, 5.0283, 5.045533, 5.070081, 5.103135, 
    5.145094, 5.195261, 5.252154, 5.308517, 5.361249, 5.407907, 5.447248, 
    5.481152, 5.508186, 5.528504, 5.5398, 5.542978, 5.537997, 5.524723, 
    5.502158, 5.472632, 5.436204, 5.394633, 5.346801, 5.294731, 5.241333, 
    5.189841, 5.143176, 5.103406, 5.07149, 5.047315, 5.029989, 5.018214, 
    5.010605, 5.005923, 5.003174, 5.001634, 5.000808, 5.000386, 5.00018, 
    5.000086,
  // momentumX(6,5, 0-49)
    5.000058, 5.000128, 5.000286, 5.000626, 5.001318, 5.002669, 5.005185, 
    5.009661, 5.017243, 5.029462, 5.048134, 5.075124, 5.1119, 5.158987, 
    5.215483, 5.279093, 5.347617, 5.408614, 5.459496, 5.498811, 5.526948, 
    5.548717, 5.563705, 5.573915, 5.578139, 5.578449, 5.57507, 5.567517, 
    5.553593, 5.534558, 5.508757, 5.477044, 5.435779, 5.385819, 5.329535, 
    5.270462, 5.212655, 5.159855, 5.114769, 5.078687, 5.051541, 5.032279, 
    5.019346, 5.011106, 5.006111, 5.003226, 5.001635, 5.000797, 5.000378, 
    5.000181,
  // momentumX(6,6, 0-49)
    5.000115, 5.000255, 5.000564, 5.001209, 5.002492, 5.00493, 5.009352, 
    5.016989, 5.029522, 5.049008, 5.077607, 5.11707, 5.168053, 5.229499, 
    5.298431, 5.370821, 5.445284, 5.502716, 5.543248, 5.567499, 5.578008, 
    5.582731, 5.581964, 5.579405, 5.574989, 5.571723, 5.570034, 5.569163, 
    5.56598, 5.56068, 5.55012, 5.534544, 5.507586, 5.468422, 5.417926, 
    5.358761, 5.295095, 5.231841, 5.173631, 5.123855, 5.084163, 5.05453, 
    5.033725, 5.019936, 5.011277, 5.006112, 5.003177, 5.001587, 5.000769, 
    5.000376,
  // momentumX(6,7, 0-49)
    5.000226, 5.000491, 5.001064, 5.002233, 5.004501, 5.008698, 5.016093, 
    5.028466, 5.048059, 5.0773, 5.118228, 5.171681, 5.236503, 5.309232, 
    5.384604, 5.457738, 5.530963, 5.576744, 5.600434, 5.605077, 5.595113, 
    5.581197, 5.563703, 5.547695, 5.534246, 5.527015, 5.526596, 5.532055, 
    5.539679, 5.548707, 5.554925, 5.558561, 5.5509, 5.529508, 5.493343, 
    5.443217, 5.382048, 5.31462, 5.246725, 5.183888, 5.130181, 5.087585, 
    5.056075, 5.034219, 5.019936, 5.011107, 5.005926, 5.003036, 5.001507, 
    5.000752,
  // momentumX(6,8, 0-49)
    5.000422, 5.000904, 5.001921, 5.003942, 5.007765, 5.014642, 5.026388, 
    5.045363, 5.074217, 5.115291, 5.169679, 5.236262, 5.311226, 5.388562, 
    5.461514, 5.526134, 5.591987, 5.620574, 5.624623, 5.609064, 5.579417, 
    5.548193, 5.515173, 5.486481, 5.46438, 5.452968, 5.453032, 5.463569, 
    5.480635, 5.502585, 5.524538, 5.547294, 5.560452, 5.560471, 5.544627, 
    5.511597, 5.462111, 5.399347, 5.328711, 5.256863, 5.190205, 5.133425, 
    5.088749, 5.056075, 5.033725, 5.019349, 5.010611, 5.00558, 5.002838, 
    5.001445,
  // momentumX(6,9, 0-49)
    5.000753, 5.001589, 5.003309, 5.006641, 5.012774, 5.023482, 5.041159, 
    5.068617, 5.108491, 5.162234, 5.228955, 5.304729, 5.382974, 5.456024, 
    5.5172, 5.565434, 5.620588, 5.629872, 5.615059, 5.581898, 5.535974, 
    5.490709, 5.444725, 5.404984, 5.375036, 5.359287, 5.358814, 5.372686, 
    5.397056, 5.429439, 5.464555, 5.504181, 5.536883, 5.558599, 5.565522, 
    5.554592, 5.52423, 5.475126, 5.410761, 5.337203, 5.261992, 5.192336, 
    5.133425, 5.087586, 5.054531, 5.032286, 5.018225, 5.009846, 5.005136, 
    5.00267,
  // momentumX(6,10, 0-49)
    5.001282, 5.002665, 5.005434, 5.010663, 5.020015, 5.035825, 5.060974, 
    5.098361, 5.149876, 5.215099, 5.290311, 5.368649, 5.441668, 5.501667, 
    5.54359, 5.570598, 5.614685, 5.605386, 5.574833, 5.52846, 5.471034, 
    5.416002, 5.360381, 5.31177, 5.275041, 5.254829, 5.25267, 5.267902, 
    5.297109, 5.337039, 5.382149, 5.435371, 5.484737, 5.526087, 5.55515, 
    5.567821, 5.560739, 5.532126, 5.482728, 5.416425, 5.34004, 5.261992, 
    5.190205, 5.130182, 5.084167, 5.051551, 5.03001, 5.016677, 5.008926, 
    5.004739,
  // momentumX(6,11, 0-49)
    5.002078, 5.004252, 5.008497, 5.016294, 5.029826, 5.051929, 5.085682, 
    5.133456, 5.195515, 5.268737, 5.346379, 5.41946, 5.479264, 5.519618, 
    5.53792, 5.542086, 5.576544, 5.550974, 5.508726, 5.454051, 5.390294, 
    5.330138, 5.268671, 5.213834, 5.171679, 5.146977, 5.141926, 5.156423, 
    5.187869, 5.232409, 5.284306, 5.34762, 5.410196, 5.467977, 5.516637, 
    5.551656, 5.568658, 5.564036, 5.535913, 5.485223, 5.416424, 5.337204, 
    5.256864, 5.183889, 5.12386, 5.078702, 5.04735, 5.027104, 5.014899, 
    5.008082,
  // momentumX(6,12, 0-49)
    5.003199, 5.006451, 5.012627, 5.023664, 5.042225, 5.071439, 5.11411, 
    5.171338, 5.240982, 5.31694, 5.390095, 5.450813, 5.491652, 5.508848, 
    5.502183, 5.484329, 5.5107, 5.471681, 5.42171, 5.363332, 5.298191, 
    5.237552, 5.174379, 5.116498, 5.070714, 5.04173, 5.032598, 5.044168, 
    5.075143, 5.121388, 5.177038, 5.247113, 5.3195, 5.390254, 5.455167, 
    5.509714, 5.549153, 5.568865, 5.565066, 5.535909, 5.482724, 5.41076, 
    5.328711, 5.246729, 5.17364, 5.114793, 5.071546, 5.042262, 5.023884, 
    5.013244,
  // momentumX(6,13, 0-49)
    5.004665, 5.00928, 5.017808, 5.032618, 5.056721, 5.093204, 5.144015, 
    5.208309, 5.2812, 5.354035, 5.416568, 5.459991, 5.479059, 5.472442, 
    5.441646, 5.404009, 5.422162, 5.372473, 5.318215, 5.260051, 5.197939, 
    5.141232, 5.080792, 5.023685, 4.976696, 4.944057, 4.92978, 4.936145, 
    4.963764, 5.008761, 5.065294, 5.139062, 5.21817, 5.298661, 5.376439, 
    5.447134, 5.506054, 5.548239, 5.568853, 5.564024, 5.532117, 5.475121, 
    5.399345, 5.314625, 5.231855, 5.159892, 5.10349, 5.063205, 5.036771, 
    5.020852,
  // momentumX(6,14, 0-49)
    5.006432, 5.012634, 5.023786, 5.042606, 5.072232, 5.115298, 5.172375, 
    5.240322, 5.311727, 5.376356, 5.424157, 5.448103, 5.445302, 5.416306, 
    5.363493, 5.308928, 5.315402, 5.257618, 5.201933, 5.147207, 5.091923, 
    5.043219, 4.99018, 4.938323, 4.893336, 4.858306, 4.838092, 4.836915, 
    4.85803, 4.898629, 4.953203, 5.027792, 5.110849, 5.19822, 5.285783, 
    5.369319, 5.444354, 5.506011, 5.549108, 5.568622, 5.560715, 5.524216, 
    5.462107, 5.382053, 5.295115, 5.212708, 5.143295, 5.09066, 5.054367, 
    5.031552,
  // momentumX(6,15, 0-49)
    5.008353, 5.01623, 5.03002, 5.052654, 5.087132, 5.135281, 5.196004, 
    5.263953, 5.329874, 5.383046, 5.414553, 5.419429, 5.396732, 5.348141, 
    5.276179, 5.207609, 5.194048, 5.130501, 5.075865, 5.027326, 4.982164, 
    4.945155, 4.904314, 4.862773, 4.823861, 4.788546, 4.762092, 4.751051, 
    4.762189, 4.794866, 4.844478, 4.917047, 5.001487, 5.09321, 5.187871, 
    5.281279, 5.369182, 5.446979, 5.509586, 5.551565, 5.567762, 5.554559, 
    5.511582, 5.443219, 5.358788, 5.270534, 5.190001, 5.124745, 5.077209, 
    5.045891,
  // momentumX(6,16, 0-49)
    5.010181, 5.019599, 5.035693, 5.061436, 5.099479, 5.150658, 5.212265, 
    5.277219, 5.335279, 5.376088, 5.392232, 5.380555, 5.341426, 5.277007, 
    5.189547, 5.10928, 5.061175, 4.993652, 4.942364, 4.902635, 4.870674, 
    4.848741, 4.82494, 4.799216, 4.771264, 4.738774, 4.706534, 4.683522, 
    4.680879, 4.701571, 4.742841, 4.810379, 4.893664, 4.987398, 5.086774, 
    5.187449, 5.285298, 5.376024, 5.45486, 5.516427, 5.555016, 5.565443, 
    5.544588, 5.493336, 5.417953, 5.329622, 5.241532, 5.164762, 5.10537, 
    5.064186,
  // momentumX(6,17, 0-49)
    5.011572, 5.022128, 5.039799, 5.067472, 5.107347, 5.159363, 5.219592, 
    5.279918, 5.329862, 5.35982, 5.363729, 5.339694, 5.288814, 5.213394, 
    5.115401, 5.023416, 4.91982, 4.848852, 4.803052, 4.775018, 4.75953, 
    4.755941, 4.754036, 4.749845, 4.738373, 4.712875, 4.676379, 4.639837, 
    4.619423, 4.623429, 4.652407, 4.711521, 4.790933, 4.884343, 4.986193, 
    5.091783, 5.19697, 5.297701, 5.389572, 5.46752, 5.525795, 5.558423, 
    5.560376, 5.529471, 5.46844, 5.385913, 5.294955, 5.209147, 5.138294, 
    5.086379,
  // momentumX(6,18, 0-49)
    5.012167, 5.023161, 5.04132, 5.069361, 5.109135, 5.160046, 5.217618, 
    5.273468, 5.317338, 5.340284, 5.337028, 5.306277, 5.249497, 5.169226, 
    5.067511, 4.957667, 4.773083, 4.697157, 4.658534, 4.645606, 4.650552, 
    4.668773, 4.693651, 4.71667, 4.727506, 4.714119, 4.676271, 4.625728, 
    4.583766, 4.56583, 4.577911, 4.624625, 4.69708, 4.787639, 4.889681, 
    4.997922, 5.108042, 5.21612, 5.318082, 5.409255, 5.484136, 5.536518, 
    5.560242, 5.550798, 5.507571, 5.435857, 5.34702, 5.255654, 5.174771, 
    5.111942,
  // momentumX(6,19, 0-49)
    5.011673, 5.022164, 5.039426, 5.06602, 5.103715, 5.152024, 5.206848, 
    5.260324, 5.302584, 5.324714, 5.321186, 5.290559, 5.234613, 5.15659, 
    5.058802, 4.913702, 4.622737, 4.538507, 4.507798, 4.513911, 4.544353, 
    4.588445, 4.64507, 4.700685, 4.73955, 4.744065, 4.709301, 4.645968, 
    4.579593, 4.53436, 4.524497, 4.554203, 4.616135, 4.700994, 4.800754, 
    4.909312, 5.022017, 5.134962, 5.244314, 5.345772, 5.434191, 5.503454, 
    5.546865, 5.558331, 5.534452, 5.477069, 5.394795, 5.301735, 5.213065, 
    5.139863,
  // momentumX(6,20, 0-49)
    5.009789, 5.018234, 5.032057, 5.053111, 5.08257, 5.119898, 5.161999, 
    5.20331, 5.237241, 5.258398, 5.264359, 5.256173, 5.237612, 5.213781, 
    5.189564, 0, 4.351584, 4.34895, 4.370693, 4.414233, 4.476791, 4.54938, 
    4.639208, 4.728305, 4.795688, 4.818511, 4.786697, 4.708689, 4.613272, 
    4.53438, 4.497091, 4.504663, 4.552106, 4.628093, 4.722847, 4.829231, 
    4.942132, 5.057541, 5.171772, 5.280826, 5.379914, 5.463161, 5.523698, 
    5.554443, 5.54987, 5.508664, 5.436234, 5.345024, 5.251167, 5.168735,
  // momentumX(6,21, 0-49)
    5.008009, 5.014865, 5.026288, 5.044007, 5.069425, 5.102808, 5.142482, 
    5.184568, 5.223716, 5.254673, 5.273949, 5.280734, 5.276828, 5.265878, 
    5.252289, 0, 4.170659, 4.190443, 4.237646, 4.309671, 4.403232, 4.505134, 
    4.625941, 4.743216, 4.833209, 4.872109, 4.84777, 4.765993, 4.654385, 
    4.551601, 4.492404, 4.478347, 4.510312, 4.576025, 4.664337, 4.767112, 
    4.878688, 4.994842, 5.111915, 5.226116, 5.33296, 5.426864, 5.501005, 
    5.547768, 5.560138, 5.534248, 5.47243, 5.384887, 5.287694, 5.197131,
  // momentumX(6,22, 0-49)
    5.006531, 5.012131, 5.021671, 5.036806, 5.059116, 5.089477, 5.127281, 
    5.16994, 5.2131, 5.25171, 5.281518, 5.300305, 5.308352, 5.308174, 
    5.303796, 0, 4.030805, 4.065196, 4.131796, 4.227709, 4.348972, 4.477757, 
    4.627515, 4.771355, 4.883232, 4.939029, 4.924598, 4.842271, 4.716929, 
    4.590865, 4.509266, 4.470721, 4.484496, 4.53761, 4.617585, 4.715239, 
    4.824254, 4.940064, 5.058887, 5.17696, 5.289956, 5.392478, 5.47778, 
    5.537942, 5.564931, 5.552924, 5.501613, 5.41886, 5.320036, 5.22286,
  // momentumX(6,23, 0-49)
    5.005608, 5.010423, 5.018781, 5.032283, 5.052613, 5.081013, 5.117546, 
    5.160475, 5.206153, 5.249742, 5.28655, 5.313443, 5.329684, 5.337036, 
    5.339309, 0, 3.936208, 3.979444, 4.05963, 4.173486, 4.31631, 4.465572, 
    4.636799, 4.799335, 4.926097, 4.994142, 4.988685, 4.909207, 4.776904, 
    4.635037, 4.536873, 4.476786, 4.473642, 4.514404, 4.585753, 4.677729, 
    4.783483, 4.898127, 5.017705, 5.138398, 5.255899, 5.364881, 5.458617, 
    5.528984, 5.567272, 5.566283, 5.52371, 5.445437, 5.345931, 5.243716,
  // momentumX(6,24, 0-49)
    5.005395, 5.009989, 5.017999, 5.030992, 5.050661, 5.078343, 5.114321, 
    5.157181, 5.203599, 5.248916, 5.288375, 5.318546, 5.338296, 5.349046, 
    5.354481, 0, 3.885182, 3.932935, 4.020948, 4.145664, 4.301788, 4.463101, 
    4.646461, 4.818689, 4.952569, 5.026831, 5.027077, 4.951261, 4.817554, 
    4.668488, 4.561754, 4.487683, 4.472909, 4.504726, 4.569493, 4.656837, 
    4.759587, 4.872656, 4.991975, 5.113683, 5.233487, 5.346098, 5.444815, 
    5.521412, 5.566805, 5.572984, 5.536391, 5.461555, 5.362166, 5.257078,
  // momentumX(6,25, 0-49)
    5.005977, 5.010957, 5.019516, 5.033198, 5.053604, 5.081876, 5.118042, 
    5.160445, 5.205666, 5.249183, 5.286569, 5.314772, 5.332943, 5.342594, 
    5.347287, 0, 3.875384, 3.92374, 4.013379, 4.140702, 4.30019, 4.464015, 
    4.64996, 4.823952, 4.9589, 5.034354, 5.036249, 4.962126, 4.829005, 
    4.67878, 4.570251, 4.491889, 4.473286, 4.501997, 4.564393, 4.650023, 
    4.75163, 4.864066, 4.983222, 5.105221, 5.225766, 5.339579, 5.439962, 
    5.518659, 5.566463, 5.575105, 5.5406, 5.46701, 5.367731, 5.261695,
  // momentumX(6,26, 0-49)
    5.007358, 5.013331, 5.023318, 5.038845, 5.061301, 5.09135, 5.128307, 
    5.169772, 5.211891, 5.250265, 5.281169, 5.302535, 5.31439, 5.318717, 
    5.319005, 0, 3.907399, 3.952108, 4.036621, 4.157588, 4.309739, 4.466147, 
    4.645107, 4.813356, 4.943969, 5.016002, 5.015329, 4.94009, 4.808348, 
    4.662022, 4.557912, 4.485681, 4.471959, 4.5043, 4.569307, 4.656758, 
    4.759554, 4.872642, 4.991968, 5.113681, 5.233484, 5.346098, 5.444815, 
    5.521413, 5.566805, 5.572984, 5.53639, 5.461555, 5.362166, 5.257078,
  // momentumX(6,27, 0-49)
    5.009464, 5.016989, 5.029191, 5.047569, 5.07317, 5.105905, 5.143998, 
    5.18394, 5.221245, 5.251712, 5.272612, 5.283283, 5.285047, 5.280668, 
    5.273688, 0, 3.984281, 4.020194, 4.092436, 4.198112, 4.332588, 4.472099, 
    4.634583, 4.789214, 4.909461, 4.973031, 4.965724, 4.887423, 4.759062, 
    4.622608, 4.529527, 4.472963, 4.471822, 4.513583, 4.585392, 4.677572, 
    4.783415, 4.898097, 5.017692, 5.138393, 5.255897, 5.36488, 5.458617, 
    5.528984, 5.567272, 5.566283, 5.52371, 5.445437, 5.345931, 5.243716,
  // momentumX(6,28, 0-49)
    5.012121, 5.021662, 5.036722, 5.058746, 5.08832, 5.12436, 5.163691, 
    5.201473, 5.232535, 5.253003, 5.261386, 5.258695, 5.247797, 5.232471, 
    5.216447, 0, 4.109945, 4.130611, 4.183319, 4.265604, 4.37358, 4.487952, 
    4.624791, 4.757003, 4.859302, 4.908553, 4.891548, 4.811182, 4.691791, 
    4.573579, 4.499115, 4.465442, 4.481968, 4.536459, 4.617074, 4.715014, 
    4.824155, 4.940021, 5.058867, 5.176952, 5.289953, 5.392476, 5.477779, 
    5.537941, 5.564931, 5.552924, 5.501613, 5.41886, 5.320036, 5.22286,
  // momentumX(6,29, 0-49)
    5.01504, 5.026921, 5.045306, 5.071594, 5.1058, 5.145628, 5.186234, 
    5.221255, 5.244844, 5.253647, 5.247667, 5.229831, 5.204763, 5.177385, 
    5.151611, 0, 4.284205, 4.28185, 4.307784, 4.359859, 4.434813, 4.518023, 
    4.622173, 4.724629, 4.802577, 4.8335, 4.806474, 4.727848, 4.624166, 
    4.531176, 4.480493, 4.472147, 4.507318, 4.574645, 4.663714, 4.766834, 
    4.878564, 4.994786, 5.11189, 5.226105, 5.332955, 5.426862, 5.501004, 
    5.547768, 5.560138, 5.534248, 5.47243, 5.384888, 5.287694, 5.197131,
  // momentumX(6,30, 0-49)
    5.01805, 5.03292, 5.056044, 5.089447, 5.133391, 5.184988, 5.237677, 
    5.28241, 5.310273, 5.315083, 5.294526, 5.249707, 5.183735, 5.100007, 
    5.000019, 4.8457, 4.545903, 4.460265, 4.430046, 4.441324, 4.48198, 
    4.537408, 4.612211, 4.688424, 4.746189, 4.764202, 4.733611, 4.662929, 
    4.579001, 4.51218, 4.48446, 4.498162, 4.54897, 4.626636, 4.722182, 
    4.82893, 4.941996, 5.057481, 5.171744, 5.280814, 5.379909, 5.463158, 
    5.523697, 5.554443, 5.54987, 5.508664, 5.436234, 5.345024, 5.251167, 
    5.168735,
  // momentumX(6,31, 0-49)
    5.019023, 5.03479, 5.059389, 5.094986, 5.141794, 5.196579, 5.252171, 
    5.298905, 5.32757, 5.332101, 5.310494, 5.263934, 5.195178, 5.107091, 
    5.00141, 4.883553, 4.684901, 4.605775, 4.566805, 4.557559, 4.570552, 
    4.598731, 4.639916, 4.681739, 4.709561, 4.707233, 4.671093, 4.611933, 
    4.553517, 4.517052, 4.514324, 4.54877, 4.613411, 4.699682, 4.800136, 
    4.909025, 5.021885, 5.134902, 5.244286, 5.345759, 5.434185, 5.503451, 
    5.546865, 5.558331, 5.534452, 5.477069, 5.394795, 5.301735, 5.213065, 
    5.139863,
  // momentumX(6,32, 0-49)
    5.018395, 5.033809, 5.058214, 5.094069, 5.14203, 5.199332, 5.259036, 
    5.311258, 5.346146, 5.356833, 5.340679, 5.298523, 5.232965, 5.146788, 
    5.041823, 4.942011, 4.822749, 4.747123, 4.69965, 4.673524, 4.664025, 
    4.668962, 4.681037, 4.693107, 4.696065, 4.679071, 4.64244, 4.597218, 
    4.562731, 4.552108, 4.569833, 4.620241, 4.694829, 4.786526, 4.889145, 
    4.997667, 5.107924, 5.216065, 5.318056, 5.409244, 5.484132, 5.536515, 
    5.560241, 5.550798, 5.507571, 5.435857, 5.34702, 5.255654, 5.174771, 
    5.111942,
  // momentumX(6,33, 0-49)
    5.016522, 5.030602, 5.0534, 5.087697, 5.134883, 5.193241, 5.256811, 
    5.316042, 5.360482, 5.382006, 5.376657, 5.344406, 5.287577, 5.209101, 
    5.111249, 5.021931, 4.958303, 4.88466, 4.830286, 4.790932, 4.763344, 
    4.748603, 4.736362, 4.723997, 4.707599, 4.681181, 4.647666, 4.616824, 
    4.603018, 4.612907, 4.64622, 4.708125, 4.789161, 4.883449, 4.985752, 
    5.091572, 5.196871, 5.297654, 5.389551, 5.46751, 5.525791, 5.558421, 
    5.560375, 5.529471, 5.46844, 5.385913, 5.294955, 5.209147, 5.138294, 
    5.086379,
  // momentumX(6,34, 0-49)
    5.013892, 5.025993, 5.046119, 5.077284, 5.121665, 5.178928, 5.244718, 
    5.310551, 5.365828, 5.401097, 5.410602, 5.392849, 5.349452, 5.283387, 
    5.197491, 5.117618, 5.088926, 5.017687, 4.958633, 4.909221, 4.867121, 
    4.835982, 4.804241, 4.772992, 4.742702, 4.71132, 4.683036, 4.66551, 
    4.668421, 4.693704, 4.738229, 4.807829, 4.892317, 4.98671, 5.086431, 
    5.187284, 5.285219, 5.375988, 5.454842, 5.516418, 5.555013, 5.565441, 
    5.544586, 5.493335, 5.417953, 5.329622, 5.241532, 5.164762, 5.10537, 
    5.064186,
  // momentumX(6,35, 0-49)
    5.010988, 5.020812, 5.037631, 5.064511, 5.10425, 5.157928, 5.223202, 
    5.293424, 5.358673, 5.408595, 5.435466, 5.43575, 5.409719, 5.359928, 
    5.289591, 5.220821, 5.212025, 5.144827, 5.083393, 5.026625, 4.973094, 
    4.928782, 4.882309, 4.837645, 4.798489, 4.765621, 4.743443, 4.737309, 
    4.752937, 4.789107, 4.841118, 4.915183, 5.000496, 5.092699, 5.187614, 
    5.281154, 5.369122, 5.446951, 5.509573, 5.55156, 5.56776, 5.554558, 
    5.511581, 5.443218, 5.358788, 5.270534, 5.190001, 5.124745, 5.077209, 
    5.045891,
  // momentumX(6,36, 0-49)
    5.008206, 5.015754, 5.029075, 5.051062, 5.084832, 5.132618, 5.194133, 
    5.265147, 5.33742, 5.400627, 5.445424, 5.465913, 5.46032, 5.430084, 
    5.378282, 5.323157, 5.325123, 5.264044, 5.202501, 5.140908, 5.078958, 
    5.024843, 4.968314, 4.915356, 4.871645, 4.839771, 4.823688, 4.826664, 
    4.851294, 4.894493, 4.950805, 5.026462, 5.110141, 5.197854, 5.285599, 
    5.369229, 5.444311, 5.505991, 5.549098, 5.568619, 5.560713, 5.524215, 
    5.462106, 5.382053, 5.295115, 5.212708, 5.143295, 5.09066, 5.054367, 
    5.031552,
  // momentumX(6,37, 0-49)
    5.005801, 5.011303, 5.021308, 5.038361, 5.065549, 5.105801, 5.160549, 
    5.228139, 5.302862, 5.375661, 5.436546, 5.477478, 5.494156, 5.486094, 
    5.455472, 5.416793, 5.425346, 5.372597, 5.313364, 5.249673, 5.182581, 
    5.122284, 5.060222, 5.003567, 4.958797, 4.929513, 4.918928, 4.928662, 
    4.958955, 5.005849, 5.063618, 5.138137, 5.217677, 5.298407, 5.37631, 
    5.447072, 5.506024, 5.548225, 5.568847, 5.564021, 5.532116, 5.475121, 
    5.399345, 5.314625, 5.231855, 5.159892, 5.10349, 5.063205, 5.036771, 
    5.020852,
  // momentumX(6,38, 0-49)
    5.003891, 5.007699, 5.014834, 5.027377, 5.048105, 5.080132, 5.126007, 
    5.186297, 5.258187, 5.335034, 5.407619, 5.466704, 5.505548, 5.521119, 
    5.513827, 5.494351, 5.508985, 5.466975, 5.412887, 5.350326, 5.281836, 
    5.219258, 5.155951, 5.099565, 5.056434, 5.03064, 5.024622, 5.038822, 
    5.071777, 5.119378, 5.175891, 5.246482, 5.319166, 5.390081, 5.455081, 
    5.509673, 5.549134, 5.568857, 5.565062, 5.535907, 5.482723, 5.41076, 
    5.32871, 5.246728, 5.17364, 5.114793, 5.071546, 5.042262, 5.023884, 
    5.013244,
  // momentumX(6,39, 0-49)
    5.002481, 5.004988, 5.009824, 5.01858, 5.03355, 5.057617, 5.093771, 
    5.144087, 5.20835, 5.282921, 5.360754, 5.432937, 5.491165, 5.529831, 
    5.546874, 5.548873, 5.571401, 5.542856, 5.497346, 5.439801, 5.37418, 
    5.313456, 5.252906, 5.200124, 5.160659, 5.138759, 5.136208, 5.152687, 
    5.185562, 5.231051, 5.283538, 5.347201, 5.409976, 5.467864, 5.516581, 
    5.55163, 5.568645, 5.56403, 5.53591, 5.485222, 5.416424, 5.337203, 
    5.256864, 5.183889, 5.12386, 5.078702, 5.04735, 5.027104, 5.014899, 
    5.008082,
  // momentumX(6,40, 0-49)
    5.001506, 5.003077, 5.006195, 5.012006, 5.022259, 5.039356, 5.066173, 
    5.105471, 5.158852, 5.225492, 5.301316, 5.379313, 5.451182, 5.50957, 
    5.549834, 5.574276, 5.607434, 5.595249, 5.56227, 5.514218, 5.45616, 
    5.401567, 5.34748, 5.301089, 5.266817, 5.248916, 5.24868, 5.265357, 
    5.295565, 5.336142, 5.381646, 5.435097, 5.484591, 5.526011, 5.555113, 
    5.567804, 5.56073, 5.532122, 5.482724, 5.416423, 5.340039, 5.261992, 
    5.190205, 5.130182, 5.084167, 5.051551, 5.03001, 5.016677, 5.008926, 
    5.004739,
  // momentumX(6,41, 0-49)
    5.000872, 5.001811, 5.003726, 5.007394, 5.014062, 5.025565, 5.044321, 
    5.073099, 5.114377, 5.169344, 5.236801, 5.312582, 5.390053, 5.461687, 
    5.521057, 5.566554, 5.612437, 5.619046, 5.602568, 5.568698, 5.523036, 
    5.478834, 5.434624, 5.396982, 5.369114, 5.355171, 5.356116, 5.371006, 
    5.396053, 5.428863, 5.464231, 5.504002, 5.536785, 5.558545, 5.565493, 
    5.554577, 5.524221, 5.475122, 5.410758, 5.337202, 5.261991, 5.192336, 
    5.133424, 5.087586, 5.054531, 5.032286, 5.018225, 5.009846, 5.005136, 
    5.00267,
  // momentumX(6,42, 0-49)
    5.000481, 5.001017, 5.00214, 5.004345, 5.008471, 5.015812, 5.028213, 
    5.048029, 5.077842, 5.119837, 5.174886, 5.241633, 5.316115, 5.392297, 
    5.463521, 5.525497, 5.583997, 5.61024, 5.613234, 5.597641, 5.568791, 
    5.538901, 5.507612, 5.480733, 5.460288, 5.450224, 5.451291, 5.462511, 
    5.480014, 5.502224, 5.524326, 5.547166, 5.560371, 5.560421, 5.544595, 
    5.511576, 5.462096, 5.399337, 5.328705, 5.25686, 5.190202, 5.133424, 
    5.088748, 5.056075, 5.033725, 5.019349, 5.010611, 5.00558, 5.002838, 
    5.001445,
  // momentumX(6,43, 0-49)
    5.000254, 5.000546, 5.001174, 5.002439, 5.00487, 5.009325, 5.017095, 
    5.029969, 5.050164, 5.080025, 5.121449, 5.175093, 5.239628, 5.311485, 
    5.385376, 5.456191, 5.523962, 5.567801, 5.590858, 5.595832, 5.586867, 
    5.574288, 5.558316, 5.543778, 5.53159, 5.525327, 5.525582, 5.531467, 
    5.539334, 5.548489, 5.55477, 5.558441, 5.550801, 5.52943, 5.493284, 
    5.443173, 5.382017, 5.3146, 5.246713, 5.18388, 5.130176, 5.087583, 
    5.056074, 5.034219, 5.019936, 5.011107, 5.005926, 5.003036, 5.001507, 
    5.000752,
  // momentumX(6,44, 0-49)
    5.000128, 5.000281, 5.000617, 5.00131, 5.002675, 5.005249, 5.009875, 
    5.017793, 5.030678, 5.050543, 5.079468, 5.119081, 5.169894, 5.230724, 
    5.298507, 5.369052, 5.439737, 5.495649, 5.53579, 5.560483, 5.571956, 
    5.577868, 5.578365, 5.576972, 5.573505, 5.570918, 5.569647, 5.568985, 
    5.565864, 5.560555, 5.549966, 5.534374, 5.507415, 5.468267, 5.417797, 
    5.358663, 5.295023, 5.231793, 5.1736, 5.123836, 5.084153, 5.054524, 
    5.033722, 5.019935, 5.011277, 5.006111, 5.003177, 5.001587, 5.000769, 
    5.000376,
  // momentumX(6,45, 0-49)
    5.000063, 5.000138, 5.000311, 5.000674, 5.001407, 5.002824, 5.005446, 
    5.010069, 5.017841, 5.03027, 5.049132, 5.07621, 5.112875, 5.159539, 
    5.21521, 5.277477, 5.343553, 5.403429, 5.454043, 5.493758, 5.522719, 
    5.545506, 5.561567, 5.57276, 5.57775, 5.578548, 5.575379, 5.567812, 
    5.55373, 5.5345, 5.508538, 5.476731, 5.435433, 5.385492, 5.329256, 
    5.270243, 5.212493, 5.159744, 5.114697, 5.078644, 5.051517, 5.032265, 
    5.019338, 5.011102, 5.00611, 5.003224, 5.001634, 5.000797, 5.000378, 
    5.000181,
  // momentumX(6,46, 0-49)
    5.000031, 5.000067, 5.00015, 5.000331, 5.000709, 5.001454, 5.002869, 
    5.005435, 5.009881, 5.017223, 5.02877, 5.046025, 5.070468, 5.103213, 
    5.144585, 5.193819, 5.249195, 5.304764, 5.3573, 5.404286, 5.444343, 
    5.479204, 5.507306, 5.528643, 5.540705, 5.544287, 5.539324, 5.525741, 
    5.502674, 5.472641, 5.435821, 5.39402, 5.3461, 5.29405, 5.24074, 
    5.189366, 5.142821, 5.103158, 5.071325, 5.047211, 5.029928, 5.018178, 
    5.010585, 5.005913, 5.00317, 5.001631, 5.000807, 5.000385, 5.000178, 
    5.000086,
  // momentumX(6,47, 0-49)
    5.000016, 5.000032, 5.000071, 5.000156, 5.000339, 5.000712, 5.00144, 
    5.002793, 5.0052, 5.009297, 5.015947, 5.026236, 5.041384, 5.062566, 
    5.090646, 5.125872, 5.167685, 5.213145, 5.259974, 5.305874, 5.348906, 
    5.388846, 5.423281, 5.450551, 5.467137, 5.472547, 5.466381, 5.448959, 
    5.420728, 5.385215, 5.34418, 5.300195, 5.253817, 5.207319, 5.163136, 
    5.123419, 5.089652, 5.062486, 5.041776, 5.026793, 5.016487, 5.009737, 
    5.005519, 5.003005, 5.001571, 5.000789, 5.000381, 5.000178, 5.000082, 
    5.00004,
  // momentumX(6,48, 0-49)
    5.00001, 5.000016, 5.000032, 5.00007, 5.000153, 5.000327, 5.000675, 
    5.00134, 5.002559, 5.004692, 5.008262, 5.013968, 5.022671, 5.035318, 
    5.052807, 5.075786, 5.104437, 5.137691, 5.174414, 5.213105, 5.252073, 
    5.290257, 5.324902, 5.35331, 5.371335, 5.377446, 5.370953, 5.352503, 
    5.323604, 5.288409, 5.249669, 5.210224, 5.171314, 5.134784, 5.102191, 
    5.074564, 5.052313, 5.035273, 5.022853, 5.014224, 5.008505, 5.004887, 
    5.002697, 5.001432, 5.000731, 5.000358, 5.00017, 5.000078, 5.000036, 
    5.000019,
  // momentumX(6,49, 0-49)
    5.000003, 5.000005, 5.00001, 5.000021, 5.000048, 5.000105, 5.000226, 
    5.000469, 5.000938, 5.001801, 5.003329, 5.005904, 5.010058, 5.016455, 
    5.025851, 5.039001, 5.056527, 5.078323, 5.104247, 5.133745, 5.165843, 
    5.199856, 5.232936, 5.261728, 5.280608, 5.287194, 5.280442, 5.261369, 
    5.232347, 5.199001, 5.164706, 5.132356, 5.102732, 5.076899, 5.055445, 
    5.038478, 5.025686, 5.016487, 5.010173, 5.006035, 5.00344, 5.001884, 
    5.000993, 5.000504, 5.000246, 5.000115, 5.000053, 5.000024, 5.000012, 
    5.000007,
  // momentumX(7,0, 0-49)
    5.000065, 5.000127, 5.000259, 5.000518, 5.001007, 5.001891, 5.003428, 
    5.005995, 5.010108, 5.016434, 5.025755, 5.038896, 5.056596, 5.079338, 
    5.107157, 5.139503, 5.175241, 5.211763, 5.247095, 5.279533, 5.307879, 
    5.331899, 5.350907, 5.364714, 5.372608, 5.374767, 5.371186, 5.361848, 
    5.346594, 5.326201, 5.300992, 5.271825, 5.239199, 5.204507, 5.169468, 
    5.135854, 5.105211, 5.078644, 5.05671, 5.039443, 5.026458, 5.017118, 
    5.010684, 5.006434, 5.003739, 5.002098, 5.001138, 5.000597, 5.000308, 
    5.000164,
  // momentumX(7,1, 0-49)
    5.000121, 5.000238, 5.00048, 5.000947, 5.001812, 5.003347, 5.005964, 
    5.010249, 5.016973, 5.027078, 5.041602, 5.061525, 5.087564, 5.119916, 
    5.158052, 5.20067, 5.245986, 5.289452, 5.328742, 5.362245, 5.389309, 
    5.411021, 5.42722, 5.438537, 5.444373, 5.445482, 5.441986, 5.433731, 
    5.419994, 5.40147, 5.377745, 5.349227, 5.315303, 5.277005, 5.236064, 
    5.194644, 5.154975, 5.118989, 5.08803, 5.062733, 5.043062, 5.028478, 
    5.018152, 5.011154, 5.00661, 5.003779, 5.002086, 5.001116, 5.000584, 
    5.000315,
  // momentumX(7,2, 0-49)
    5.000235, 5.000459, 5.00091, 5.001763, 5.003306, 5.005982, 5.010434, 
    5.017533, 5.028368, 5.04416, 5.066104, 5.095097, 5.131435, 5.174539, 
    5.222845, 5.274029, 5.325931, 5.371635, 5.409235, 5.437857, 5.457925, 
    5.47228, 5.481415, 5.48696, 5.488639, 5.487854, 5.484875, 5.479411, 
    5.470135, 5.457471, 5.440103, 5.41785, 5.388554, 5.352391, 5.310528, 
    5.264997, 5.218402, 5.17348, 5.132623, 5.097514, 5.068947, 5.046889, 
    5.030686, 5.019336, 5.011737, 5.006867, 5.003877, 5.00212, 5.001133, 
    5.000619,
  // momentumX(7,3, 0-49)
    5.000447, 5.000865, 5.001686, 5.003202, 5.005878, 5.010405, 5.017734, 
    5.029084, 5.045851, 5.069425, 5.100871, 5.14055, 5.18778, 5.240693, 
    5.296419, 5.351787, 5.405229, 5.447082, 5.476982, 5.495352, 5.503921, 
    5.507381, 5.506683, 5.504385, 5.500591, 5.497306, 5.494962, 5.493176, 
    5.490098, 5.485869, 5.478354, 5.466926, 5.447763, 5.419919, 5.383484, 
    5.339691, 5.290837, 5.239985, 5.190429, 5.145115, 5.106135, 5.074507, 
    5.050228, 5.032541, 5.020276, 5.012163, 5.007035, 5.003933, 5.00215, 
    5.001194,
  // momentumX(7,4, 0-49)
    5.00083, 5.001577, 5.003015, 5.005607, 5.010071, 5.01742, 5.028973, 
    5.046284, 5.070925, 5.104134, 5.146344, 5.196767, 5.253208, 5.312281, 
    5.370041, 5.423226, 5.472451, 5.504696, 5.522296, 5.52714, 5.522073, 
    5.513369, 5.501997, 5.491229, 5.481532, 5.475423, 5.473501, 5.47537, 
    5.478836, 5.483813, 5.487583, 5.489424, 5.484031, 5.469409, 5.444396, 
    5.408932, 5.364272, 5.312967, 5.258545, 5.204911, 5.155597, 5.11315, 
    5.078824, 5.052646, 5.033748, 5.020789, 5.012327, 5.007061, 5.003947, 
    5.002234,
  // momentumX(7,5, 0-49)
    5.00148, 5.002769, 5.005187, 5.009442, 5.016574, 5.027974, 5.045319, 
    5.070355, 5.104497, 5.148292, 5.200894, 5.259817, 5.321171, 5.380404, 
    5.433293, 5.477595, 5.517872, 5.536584, 5.539735, 5.53039, 5.512024, 
    5.492009, 5.470812, 5.452157, 5.436851, 5.427817, 5.425859, 5.430663, 
    5.439898, 5.453335, 5.467922, 5.483245, 5.492867, 5.494058, 5.484577, 
    5.462999, 5.429098, 5.384137, 5.330914, 5.273443, 5.216244, 5.163455, 
    5.118066, 5.081542, 5.053911, 5.034173, 5.020812, 5.012223, 5.006996, 
    5.004036,
  // momentumX(7,6, 0-49)
    5.002537, 5.004672, 5.008571, 5.015256, 5.026145, 5.042995, 5.067703, 
    5.101876, 5.146226, 5.199944, 5.260352, 5.323129, 5.38313, 5.435542, 
    5.476911, 5.507005, 5.535779, 5.539415, 5.528361, 5.50633, 5.476847, 
    5.447856, 5.418829, 5.393694, 5.373574, 5.361693, 5.35911, 5.365716, 
    5.379266, 5.39945, 5.423106, 5.450462, 5.474294, 5.491517, 5.499191, 
    5.494801, 5.476672, 5.444415, 5.399313, 5.344433, 5.284281, 5.224, 
    5.16831, 5.120595, 5.082476, 5.053929, 5.033796, 5.020385, 5.011956, 
    5.007038,
  // momentumX(7,7, 0-49)
    5.004174, 5.007567, 5.013592, 5.023635, 5.039485, 5.063149, 5.09643, 
    5.140269, 5.194015, 5.254954, 5.318458, 5.378851, 5.430717, 5.47008, 
    5.495052, 5.507923, 5.524962, 5.513952, 5.490565, 5.458614, 5.421184, 
    5.386325, 5.352101, 5.322395, 5.298602, 5.284111, 5.280297, 5.287394, 
    5.303493, 5.328266, 5.358603, 5.39561, 5.431551, 5.463284, 5.487547, 
    5.501169, 5.501382, 5.486283, 5.455358, 5.409954, 5.353441, 5.290848, 
    5.227934, 5.169954, 5.120609, 5.081582, 5.052734, 5.032722, 5.019694, 
    5.011834,
  // momentumX(7,8, 0-49)
    5.006591, 5.011756, 5.020663, 5.035065, 5.057024, 5.088521, 5.130782, 
    5.183451, 5.243975, 5.307598, 5.368227, 5.41984, 5.457864, 5.479952, 
    5.486041, 5.480951, 5.487695, 5.463608, 5.430469, 5.391768, 5.349826, 
    5.31244, 5.275925, 5.243874, 5.217835, 5.201171, 5.195599, 5.201853, 
    5.21865, 5.245731, 5.280169, 5.3241, 5.369467, 5.413232, 5.452092, 
    5.482594, 5.501349, 5.505374, 5.492573, 5.462371, 5.416243, 5.357937, 
    5.29305, 5.227945, 5.16834, 5.118135, 5.078969, 5.050519, 5.031245, 
    5.019186,
  // momentumX(7,9, 0-49)
    5.009975, 5.017505, 5.030089, 5.049776, 5.078679, 5.118333, 5.168806, 
    5.227921, 5.291047, 5.351834, 5.403693, 5.44137, 5.461924, 5.464885, 
    5.451752, 5.429615, 5.428216, 5.392973, 5.352669, 5.310205, 5.26699, 
    5.230297, 5.194464, 5.162518, 5.135951, 5.117805, 5.110119, 5.114284, 
    5.12995, 5.157085, 5.193079, 5.241197, 5.293196, 5.346199, 5.396987, 
    5.442087, 5.477869, 5.500757, 5.507577, 5.49611, 5.465787, 5.418324, 
    5.357944, 5.290869, 5.224051, 5.163567, 5.113378, 5.074952, 5.047724, 
    5.029982,
  // momentumX(7,10, 0-49)
    5.01446, 5.02496, 5.041936, 5.067563, 5.103665, 5.150827, 5.207461, 
    5.269351, 5.330144, 5.382782, 5.421267, 5.441902, 5.443639, 5.42762, 
    5.396376, 5.358976, 5.351389, 5.30677, 5.26151, 5.217797, 5.176116, 
    5.143035, 5.110799, 5.081596, 5.056532, 5.03793, 5.028039, 5.029017, 
    5.041786, 5.066779, 5.101882, 5.151564, 5.207518, 5.267011, 5.326935, 
    5.383892, 5.434252, 5.474237, 5.500106, 5.508534, 5.497243, 5.465786, 
    5.416254, 5.353475, 5.284362, 5.216415, 5.155936, 5.106784, 5.070136, 
    5.045145,
  // momentumX(7,11, 0-49)
    5.020058, 5.034059, 5.055914, 5.087668, 5.130448, 5.183438, 5.24315, 
    5.303562, 5.357356, 5.397788, 5.420244, 5.422883, 5.40632, 5.37279, 
    5.325267, 5.274648, 5.261842, 5.209301, 5.160816, 5.117825, 5.079991, 
    5.053068, 5.027225, 5.003541, 4.982328, 4.9647, 4.952865, 4.949788, 
    4.957981, 4.978666, 5.010483, 5.059205, 5.116598, 5.180028, 5.246441, 
    5.312511, 5.374698, 5.429252, 5.472255, 5.499822, 5.50852, 5.4961, 
    5.46238, 5.410001, 5.344549, 5.27369, 5.205394, 5.146018, 5.099126, 
    5.065478,
  // momentumX(7,12, 0-49)
    5.026608, 5.044453, 5.071303, 5.108771, 5.156913, 5.213257, 5.272523, 
    5.327488, 5.37078, 5.396759, 5.402548, 5.387994, 5.354888, 5.305989, 
    5.244225, 5.182299, 5.163545, 5.104256, 5.053853, 5.013101, 4.980991, 
    4.962399, 4.945583, 4.930279, 4.915555, 4.900771, 4.887709, 4.880032, 
    4.882082, 4.896287, 4.922391, 4.967634, 5.024047, 5.089039, 5.159525, 
    5.232173, 5.303509, 5.369896, 5.427476, 5.472199, 5.500046, 5.507537, 
    5.492572, 5.455415, 5.399471, 5.33125, 5.259198, 5.191624, 5.134699, 
    5.091459,
  // momentumX(7,13, 0-49)
    5.033735, 5.05548, 5.086987, 5.129162, 5.180753, 5.237656, 5.293234, 
    5.339825, 5.370763, 5.381915, 5.372065, 5.342326, 5.295123, 5.233254, 
    5.159248, 5.08756, 5.059693, 4.994692, 4.943421, 4.906126, 4.881305, 
    4.872905, 4.867583, 4.863523, 4.858131, 4.848498, 4.835467, 4.823103, 
    4.817653, 4.823181, 4.841021, 4.880143, 4.933115, 4.997382, 5.069714, 
    5.146647, 5.224686, 5.300283, 5.36973, 5.429057, 5.474072, 5.500647, 
    5.505333, 5.486337, 5.44461, 5.384568, 5.313798, 5.241476, 5.176003, 
    5.123024,
  // momentumX(7,14, 0-49)
    5.040861, 5.066214, 5.101596, 5.147029, 5.199935, 5.254867, 5.304424, 
    5.34119, 5.35965, 5.357197, 5.333939, 5.29176, 5.233256, 5.160916, 
    5.076638, 4.99614, 4.952772, 4.88308, 4.831912, 4.799187, 4.783082, 
    4.786512, 4.794985, 4.804932, 4.811784, 4.809976, 4.798848, 4.782353, 
    4.768427, 4.763132, 4.769983, 4.80008, 4.846959, 4.908147, 4.980169, 
    5.059281, 5.141819, 5.224236, 5.302959, 5.374205, 5.433871, 5.477612, 
    5.501223, 5.501401, 5.476885, 5.429611, 5.365265, 5.292587, 5.221282, 
    5.159416,
  // momentumX(7,15, 0-49)
    5.04727, 5.075588, 5.113734, 5.160819, 5.213135, 5.26433, 5.306828, 
    5.333897, 5.341276, 5.327645, 5.294003, 5.242578, 5.175807, 5.095669, 
    5.003297, 4.913842, 4.844732, 4.771318, 4.721283, 4.694343, 4.688432, 
    4.705205, 4.729593, 4.756072, 4.777933, 4.786829, 4.780121, 4.760928, 
    4.738266, 4.720271, 4.713288, 4.731091, 4.768864, 4.824393, 4.893883, 
    4.973128, 5.058129, 5.145205, 5.230836, 5.311429, 5.383089, 5.441543, 
    5.482284, 5.501088, 5.494987, 5.46355, 5.410028, 5.341596, 5.268045, 
    5.19916,
  // momentumX(7,16, 0-49)
    5.052221, 5.082582, 5.122238, 5.169528, 5.219952, 5.266737, 5.302544, 
    5.321485, 5.320392, 5.298859, 5.258375, 5.201202, 5.129457, 5.044556, 
    4.946846, 4.846074, 4.737124, 4.660678, 4.612901, 4.593229, 4.599227, 
    4.630776, 4.672967, 4.718068, 4.757268, 4.779699, 4.780499, 4.761142, 
    4.730637, 4.698801, 4.675304, 4.677201, 4.702387, 4.749299, 4.813816, 
    4.891094, 4.976588, 5.066315, 5.156695, 5.244262, 5.325356, 5.395911, 
    5.45143, 5.487248, 5.499257, 5.485078, 5.445483, 5.385374, 5.313462, 
    5.240213,
  // momentumX(7,17, 0-49)
    5.055084, 5.086399, 5.126359, 5.172816, 5.22089, 5.263784, 5.294598, 
    5.308188, 5.302143, 5.27656, 5.233084, 5.173849, 5.100662, 5.014484, 
    4.914962, 4.796424, 4.630887, 4.5516, 4.507199, 4.496636, 4.516641, 
    4.564325, 4.625845, 4.690973, 4.749099, 4.787496, 4.799221, 4.783396, 
    4.747558, 4.702156, 4.66026, 4.64256, 4.651261, 4.686162, 4.742951, 
    4.81599, 4.899972, 4.990417, 5.083542, 5.175914, 5.264064, 5.344178, 
    5.411934, 5.462564, 5.491307, 5.494365, 5.470315, 5.421548, 5.354854, 
    5.280277,
  // momentumX(7,18, 0-49)
    5.055455, 5.086561, 5.125804, 5.170914, 5.217056, 5.257705, 5.286389, 
    5.298403, 5.291608, 5.26616, 5.223593, 5.165879, 5.094666, 5.010685, 
    4.912883, 4.764289, 4.52522, 4.443193, 4.403152, 4.403866, 4.440429, 
    4.50552, 4.587378, 4.673081, 4.750764, 4.806866, 4.832855, 4.825094, 
    4.788147, 4.731499, 4.671028, 4.630623, 4.61889, 4.638094, 4.684124, 
    4.750472, 4.830854, 4.920098, 5.014065, 5.109241, 5.202271, 5.289577, 
    5.367074, 5.430085, 5.473558, 5.492756, 5.484509, 5.448822, 5.390132, 
    5.31718,
  // momentumX(7,19, 0-49)
    5.053221, 5.082938, 5.120615, 5.164308, 5.209677, 5.250699, 5.281166, 
    5.296271, 5.293453, 5.272348, 5.234126, 5.180676, 5.113756, 5.033909, 
    4.938658, 4.742922, 4.415196, 4.33217, 4.297563, 4.311978, 4.368104, 
    4.45188, 4.554541, 4.660558, 4.75763, 4.832474, 4.875569, 4.880461, 
    4.847667, 4.784114, 4.707324, 4.64267, 4.607326, 4.607371, 4.639596, 
    4.696743, 4.771411, 4.857562, 4.950556, 5.046688, 5.142635, 5.234991, 
    5.319911, 5.392896, 5.448824, 5.4824, 5.489161, 5.467055, 5.418115, 
    5.349228,
  // momentumX(7,20, 0-49)
    5.047519, 5.072911, 5.105344, 5.143125, 5.182673, 5.219129, 5.247638, 
    5.264693, 5.268921, 5.261077, 5.243481, 5.219299, 5.191885, 5.164235, 
    5.138397, 0, 4.114454, 4.114334, 4.146542, 4.211831, 4.306983, 4.4182, 
    4.544752, 4.671088, 4.786033, 4.877743, 4.936459, 4.953573, 4.925799, 
    4.857228, 4.766321, 4.677095, 4.616313, 4.594654, 4.610526, 4.65621, 
    4.723191, 4.804475, 4.894822, 4.990243, 5.087366, 5.182891, 5.273173, 
    5.353907, 5.420018, 5.465905, 5.486187, 5.477157, 5.438637, 5.375458,
  // momentumX(7,21, 0-49)
    5.042906, 5.065928, 5.096264, 5.132921, 5.173195, 5.212954, 5.247571, 
    5.273136, 5.287375, 5.289968, 5.282302, 5.266943, 5.247061, 5.225951, 
    5.206573, 0, 3.960332, 3.978011, 4.033281, 4.12433, 4.2451, 4.375662, 
    4.518851, 4.658369, 4.784651, 4.88853, 4.961393, 4.993842, 4.979385, 
    4.918301, 4.827318, 4.723927, 4.643672, 4.602317, 4.601614, 4.634759, 
    4.692778, 4.76789, 4.85425, 4.947518, 5.044199, 5.141039, 5.234534, 
    5.320562, 5.394155, 5.449563, 5.480793, 5.482881, 5.453789, 5.39637,
  // momentumX(7,22, 0-49)
    5.039219, 5.060489, 5.089365, 5.125412, 5.166588, 5.209273, 5.24895, 
    5.281309, 5.303318, 5.313817, 5.313527, 5.304658, 5.290368, 5.274252, 
    5.259961, 0, 3.835406, 3.868202, 3.942687, 4.05515, 4.197188, 4.343217, 
    4.499814, 4.650155, 4.786009, 4.900363, 4.985329, 5.030774, 5.027747, 
    4.973923, 4.885179, 4.770913, 4.6747, 4.616134, 4.600175, 4.62134, 
    4.670562, 4.739481, 4.821707, 4.912546, 5.008337, 5.105797, 5.201505, 
    5.291459, 5.370781, 5.433647, 5.473652, 5.484908, 5.46392, 5.41185,
  // momentumX(7,23, 0-49)
    5.037024, 5.057234, 5.085255, 5.120999, 5.162849, 5.207517, 5.250546, 
    5.287356, 5.314402, 5.329967, 5.334363, 5.329612, 5.318913, 5.30611, 
    5.295335, 0, 3.75083, 3.794178, 3.882296, 4.009888, 4.166729, 4.322514, 
    4.487185, 4.643687, 4.784962, 4.90581, 4.999001, 5.054017, 5.060269, 
    5.013733, 4.929824, 4.809685, 4.70313, 4.632049, 4.604081, 4.615284, 
    4.656912, 4.720334, 4.798786, 4.887294, 4.982037, 5.079676, 5.176805, 
    5.269478, 5.352865, 5.421083, 5.467453, 5.485446, 5.470525, 5.42257,
  // momentumX(7,24, 0-49)
    5.036716, 5.05663, 5.084397, 5.120026, 5.162042, 5.207297, 5.25141, 
    5.289758, 5.318656, 5.336201, 5.342546, 5.339622, 5.330624, 5.319474, 
    5.310493, 0, 3.710093, 3.758837, 3.854186, 3.98978, 4.154303, 4.314251, 
    4.482039, 4.640524, 4.783451, 4.906882, 5.004126, 5.064573, 5.076762, 
    5.03577, 4.956805, 4.834767, 4.72329, 4.645191, 4.609799, 4.614413, 
    4.65074, 4.710127, 4.785641, 4.872161, 4.96578, 5.063129, 5.160812, 
    5.254916, 5.340633, 5.41205, 5.462324, 5.484553, 5.473571, 5.428463,
  // momentumX(7,25, 0-49)
    5.038471, 5.058876, 5.086976, 5.122606, 5.164133, 5.208367, 5.251034, 
    5.287758, 5.315138, 5.33149, 5.337061, 5.33376, 5.324667, 5.313553, 
    5.304569, 0, 3.712392, 3.76137, 3.857336, 3.993675, 4.158824, 4.318006, 
    4.484923, 4.642324, 4.784227, 4.907133, 5.004549, 5.065886, 5.079467, 
    5.040195, 4.963305, 4.841302, 4.72898, 4.649186, 4.611698, 4.614275, 
    4.648862, 4.706868, 4.781345, 4.867144, 4.960334, 5.057543, 5.155376, 
    5.249931, 5.336409, 5.408885, 5.460465, 5.484119, 5.474478, 5.430358,
  // momentumX(7,26, 0-49)
    5.042217, 5.063863, 5.092844, 5.128556, 5.168951, 5.210625, 5.24946, 
    5.281579, 5.304241, 5.31635, 5.31849, 5.312615, 5.301614, 5.288908, 
    5.278151, 0, 3.755883, 3.80003, 3.890133, 4.020155, 4.179138, 4.333121, 
    4.495686, 4.649438, 4.788105, 4.907743, 5.001677, 5.059398, 5.069646, 
    5.02778, 4.949212, 4.828493, 4.718805, 4.642381, 4.608218, 4.613591, 
    4.650334, 4.709931, 4.785549, 4.872119, 4.96576, 5.06312, 5.160808, 
    5.254914, 5.340632, 5.412049, 5.462324, 5.484553, 5.473571, 5.428463,
  // momentumX(7,27, 0-49)
    5.047648, 5.071205, 5.101556, 5.137453, 5.176219, 5.214128, 5.247229, 
    5.272307, 5.287539, 5.292675, 5.288845, 5.278172, 5.26337, 5.247412, 
    5.233242, 0, 3.837907, 3.872372, 3.950503, 4.067498, 4.213774, 4.358329, 
    4.513062, 4.660518, 4.793601, 4.907108, 4.993864, 5.043576, 5.046104, 
    4.997985, 4.914999, 4.797587, 4.69459, 4.626752, 4.60112, 4.613746, 
    4.65615, 4.719967, 4.798612, 4.887213, 4.981999, 5.079659, 5.176796, 
    5.269475, 5.352864, 5.421082, 5.467452, 5.485446, 5.470524, 5.42257,
  // momentumX(7,28, 0-49)
    5.054279, 5.08032, 5.1125, 5.148775, 5.185695, 5.219107, 5.245215, 
    5.261521, 5.267226, 5.263089, 5.25097, 5.233331, 5.212831, 5.192018, 
    5.172996, 0, 3.95486, 3.975625, 4.036456, 4.134297, 4.261631, 4.392307, 
    4.535101, 4.672795, 4.797129, 4.90109, 4.976916, 5.014869, 5.006731, 
    4.951005, 4.863965, 4.753953, 4.662951, 4.608952, 4.596192, 4.619275, 
    4.669537, 4.738986, 4.821471, 4.912435, 5.008284, 5.105772, 5.201493, 
    5.291453, 5.370779, 5.433645, 5.473652, 5.484908, 5.46392, 5.41185,
  // momentumX(7,29, 0-49)
    5.061519, 5.090569, 5.125088, 5.162135, 5.197347, 5.22602, 5.244443, 
    5.250815, 5.245413, 5.230116, 5.207698, 5.181172, 5.153317, 5.126302, 
    5.101217, 0, 4.100039, 4.105047, 4.144559, 4.218102, 4.320959, 4.433148, 
    4.559563, 4.683653, 4.795854, 4.887011, 4.948723, 4.97219, 4.951942, 
    4.889277, 4.801144, 4.70358, 4.629909, 4.594042, 4.597061, 4.6324, 
    4.6916, 4.767314, 4.853972, 4.947385, 5.044137, 5.141009, 5.23452, 
    5.320555, 5.394152, 5.449561, 5.480793, 5.482881, 5.453789, 5.396369,
  // momentumX(7,30, 0-49)
    5.069942, 5.104444, 5.145037, 5.188226, 5.228665, 5.260446, 5.278681, 
    5.280539, 5.265384, 5.23421, 5.188872, 5.131349, 5.06307, 4.983942, 
    4.890614, 4.694397, 4.378685, 4.306954, 4.281877, 4.30549, 4.370964, 
    4.459809, 4.568273, 4.679267, 4.780853, 4.860884, 4.909776, 4.919673, 
    4.888474, 4.82117, 4.735869, 4.654694, 4.601761, 4.586124, 4.605887, 
    4.653808, 4.721985, 4.803879, 4.89453, 4.990101, 5.087297, 5.182858, 
    5.273158, 5.353899, 5.420014, 5.465903, 5.486187, 5.477157, 5.438637, 
    5.375458,
  // momentumX(7,31, 0-49)
    5.073872, 5.110393, 5.153061, 5.197888, 5.238931, 5.269813, 5.28551, 
    5.283435, 5.26344, 5.227028, 5.17638, 5.113566, 5.040033, 4.956133, 
    4.860312, 4.711382, 4.476999, 4.403505, 4.371749, 4.381316, 4.427418, 
    4.499416, 4.589086, 4.681817, 4.765648, 4.827684, 4.859194, 4.855018, 
    4.817186, 4.75356, 4.681082, 4.623222, 4.59458, 4.599795, 4.6354, 
    4.694525, 4.770272, 4.856986, 4.950268, 5.046546, 5.142564, 5.234956, 
    5.319895, 5.392888, 5.448821, 5.482398, 5.48916, 5.467055, 5.418115, 
    5.349227,
  // momentumX(7,32, 0-49)
    5.074563, 5.111968, 5.156186, 5.203183, 5.24673, 5.279979, 5.297396, 
    5.296023, 5.275575, 5.23764, 5.184599, 5.118748, 5.041742, 4.954269, 
    4.855663, 4.736937, 4.571723, 4.498174, 4.459996, 4.456672, 4.485158, 
    4.540483, 4.610906, 4.684608, 4.750361, 4.79529, 4.81181, 4.797491, 
    4.758013, 4.70317, 4.647774, 4.613843, 4.608014, 4.631615, 4.680494, 
    4.748522, 4.829835, 4.919573, 5.013799, 5.109106, 5.202204, 5.289543, 
    5.367058, 5.430077, 5.473555, 5.492754, 5.484507, 5.448821, 5.390131, 
    5.31718,
  // momentumX(7,33, 0-49)
    5.072055, 5.109157, 5.154137, 5.203316, 5.250513, 5.288494, 5.311002, 
    5.31429, 5.297483, 5.261912, 5.210007, 5.14432, 5.066876, 4.978845, 
    4.880323, 4.778907, 4.66792, 4.594558, 4.550687, 4.536237, 4.549191, 
    4.588276, 4.639575, 4.693966, 4.741624, 4.770691, 4.775239, 4.755387, 
    4.719284, 4.677091, 4.640542, 4.628673, 4.642346, 4.680838, 4.739939, 
    4.814349, 4.8991, 4.989961, 5.083307, 5.175795, 5.264003, 5.344147, 
    5.411918, 5.462556, 5.491303, 5.494362, 5.470314, 5.421547, 5.354854, 
    5.280277,
  // momentumX(7,34, 0-49)
    5.066685, 5.102252, 5.146866, 5.197575, 5.248649, 5.292713, 5.322759, 
    5.333969, 5.324487, 5.295034, 5.247876, 5.185752, 5.11112, 5.025746, 
    4.930516, 4.839296, 4.766814, 4.694075, 4.645786, 4.622183, 4.62171, 
    4.645421, 4.67846, 4.714131, 4.744484, 4.759594, 4.755527, 4.734432, 
    4.705405, 4.677551, 4.65919, 4.666082, 4.695303, 4.745059, 4.811397, 
    4.889759, 4.975869, 5.065935, 5.156497, 5.244161, 5.325305, 5.395886, 
    5.451417, 5.487242, 5.499254, 5.485077, 5.445483, 5.385374, 5.313462, 
    5.240213,
  // momentumX(7,35, 0-49)
    5.059091, 5.091941, 5.134801, 5.18574, 5.23992, 5.290249, 5.329171, 
    5.350695, 5.351656, 5.331776, 5.292833, 5.237574, 5.16882, 5.088939, 
    4.999584, 4.915709, 4.867932, 4.796804, 4.745568, 4.71463, 4.70265, 
    4.712214, 4.728501, 4.746943, 4.761694, 4.765309, 4.755863, 4.73676, 
    4.716686, 4.702873, 4.700494, 4.722412, 4.763369, 4.821098, 4.89199, 
    4.972076, 5.057559, 5.144899, 5.230677, 5.311346, 5.383048, 5.441524, 
    5.482273, 5.501082, 5.494984, 5.463549, 5.410028, 5.341596, 5.268045, 
    5.19916,
  // momentumX(7,36, 0-49)
    5.050116, 5.079262, 5.118917, 5.168323, 5.223925, 5.279467, 5.327296, 
    5.360398, 5.374112, 5.366771, 5.339256, 5.293997, 5.233984, 5.162076, 
    5.080613, 5.003589, 4.970191, 4.901921, 4.849092, 4.81234, 4.790542, 
    4.787408, 4.788884, 4.792263, 4.793777, 4.788606, 4.776517, 4.761394, 
    4.750595, 4.749277, 4.760054, 4.793442, 4.842779, 4.90564, 4.978724, 
    5.058472, 5.141376, 5.223999, 5.302834, 5.37414, 5.433838, 5.477597, 
    5.501214, 5.501397, 5.476884, 5.429609, 5.365265, 5.292587, 5.221282, 
    5.159416,
  // momentumX(7,37, 0-49)
    5.040674, 5.065457, 5.100637, 5.146596, 5.201307, 5.259878, 5.315217, 
    5.359754, 5.387404, 5.394824, 5.381534, 5.34921, 5.300679, 5.239072, 
    5.167283, 5.097776, 5.072126, 5.007897, 4.954634, 4.913358, 4.883272, 
    4.869039, 4.857895, 4.848771, 4.839742, 4.828416, 4.815767, 4.805543, 
    4.803319, 4.812391, 4.833456, 4.87515, 4.92999, 4.995509, 5.06863, 
    5.146039, 5.224351, 5.300103, 5.369635, 5.429007, 5.474048, 5.500636, 
    5.505328, 5.486333, 5.444608, 5.384567, 5.313798, 5.241476, 5.176003, 
    5.123024,
  // momentumX(7,38, 0-49)
    5.031587, 5.051754, 5.081593, 5.122414, 5.173713, 5.232343, 5.292474, 
    5.346719, 5.387997, 5.411265, 5.414304, 5.39752, 5.363111, 5.314147, 
    5.253855, 5.193147, 5.17178, 5.112633, 5.059998, 5.015416, 4.978568, 
    4.954986, 4.933573, 4.914676, 4.897844, 4.882706, 4.870935, 4.86574, 
    4.870833, 4.888049, 4.916724, 4.963934, 5.021742, 5.087658, 5.158724, 
    5.231721, 5.303259, 5.369761, 5.427405, 5.472163, 5.500027, 5.507529, 
    5.492567, 5.455412, 5.39947, 5.33125, 5.259198, 5.191624, 5.134699, 
    5.091459,
  // momentumX(7,39, 0-49)
    5.023478, 5.03917, 5.063326, 5.09785, 5.143517, 5.198998, 5.260269, 
    5.32098, 5.373845, 5.412485, 5.432821, 5.433532, 5.415639, 5.38168, 
    5.334877, 5.284673, 5.266556, 5.213517, 5.162659, 5.11611, 5.074186, 
    5.043216, 5.01401, 4.988095, 4.966056, 4.949053, 4.939028, 4.938462, 
    4.949347, 4.97249, 5.0063, 5.056495, 5.114914, 5.179015, 5.245848, 
    5.312171, 5.374506, 5.429146, 5.472199, 5.499791, 5.508503, 5.496091, 
    5.462376, 5.409999, 5.344549, 5.273689, 5.205394, 5.146018, 5.099126, 
    5.065478,
  // momentumX(7,40, 0-49)
    5.01671, 5.028383, 5.047037, 5.074806, 5.113331, 5.162851, 5.22134, 
    5.284199, 5.344914, 5.396571, 5.433529, 5.452536, 5.452931, 5.436152, 
    5.404949, 5.367265, 5.35313, 5.307418, 5.259766, 5.2129, 5.167883, 
    5.131764, 5.097353, 5.067103, 5.04221, 5.024868, 5.016986, 5.020291, 
    5.035318, 5.062237, 5.098837, 5.149593, 5.206281, 5.266251, 5.326477, 
    5.383618, 5.434089, 5.474142, 5.500051, 5.508503, 5.497226, 5.465776, 
    5.416249, 5.353471, 5.28436, 5.216414, 5.155935, 5.106784, 5.070136, 
    5.045145,
  // momentumX(7,41, 0-49)
    5.011393, 5.019699, 5.033443, 5.054687, 5.08547, 5.127131, 5.179427, 
    5.239829, 5.303455, 5.363914, 5.414792, 5.451157, 5.470404, 5.472347, 
    5.458686, 5.435668, 5.427438, 5.390626, 5.348041, 5.302955, 5.257243, 
    5.218533, 5.181604, 5.149585, 5.123898, 5.107349, 5.101637, 5.107809, 
    5.125257, 5.153823, 5.190883, 5.239744, 5.292246, 5.345578, 5.396583, 
    5.44182, 5.477694, 5.500643, 5.507504, 5.496064, 5.465759, 5.418307, 
    5.357935, 5.290864, 5.224049, 5.163566, 5.113376, 5.074951, 5.047723, 
    5.029982,
  // momentumX(7,42, 0-49)
    5.007448, 5.013103, 5.022773, 5.03824, 5.061559, 5.094617, 5.138445, 
    5.192428, 5.253744, 5.317492, 5.377594, 5.428209, 5.465016, 5.485915, 
    5.491031, 5.484582, 5.484806, 5.458848, 5.423669, 5.382972, 5.339408, 
    5.300989, 5.264325, 5.232959, 5.208259, 5.193301, 5.189502, 5.197357, 
    5.215441, 5.243477, 5.278582, 5.322964, 5.368637, 5.412613, 5.451626, 
    5.482244, 5.501094, 5.50519, 5.492446, 5.462286, 5.416188, 5.357902, 
    5.293029, 5.227933, 5.168333, 5.118133, 5.078968, 5.050518, 5.031245, 
    5.019185,
  // momentumX(7,43, 0-49)
    5.004671, 5.00836, 5.014862, 5.025596, 5.042367, 5.06715, 5.101645, 
    5.146619, 5.201205, 5.262506, 5.325803, 5.385471, 5.436242, 5.474329, 
    5.498009, 5.509168, 5.520347, 5.507353, 5.482279, 5.449014, 5.41083, 
    5.375861, 5.342307, 5.313881, 5.291713, 5.278893, 5.276544, 5.284764, 
    5.301612, 5.326838, 5.35743, 5.394591, 5.430645, 5.462481, 5.486856, 
    5.500595, 5.500926, 5.485937, 5.455106, 5.409778, 5.353324, 5.290773, 
    5.22789, 5.169929, 5.120594, 5.081575, 5.05273, 5.03272, 5.019693, 
    5.011834,
  // momentumX(7,44, 0-49)
    5.002813, 5.005119, 5.009302, 5.016413, 5.027887, 5.045482, 5.071043, 
    5.106079, 5.151144, 5.205262, 5.265625, 5.327862, 5.386883, 5.437991, 
    5.477863, 5.506032, 5.529777, 5.531497, 5.519186, 5.496544, 5.467158, 
    5.438933, 5.411334, 5.388013, 5.36974, 5.359428, 5.357933, 5.365097, 
    5.378753, 5.398783, 5.422194, 5.449341, 5.473051, 5.490255, 5.498004, 
    5.493757, 5.475805, 5.443734, 5.398806, 5.344073, 5.284039, 5.223843, 
    5.168211, 5.120537, 5.082442, 5.053911, 5.033787, 5.020379, 5.011954, 
    5.007036,
  // momentumX(7,45, 0-49)
    5.001627, 5.00301, 5.005588, 5.010087, 5.017568, 5.029425, 5.047313, 
    5.072919, 5.10756, 5.151648, 5.204203, 5.262649, 5.32308, 5.380993, 
    5.432267, 5.474555, 5.510695, 5.527712, 5.530097, 5.520863, 5.503451, 
    5.485116, 5.466168, 5.449955, 5.436787, 5.429237, 5.42793, 5.432586, 
    5.441073, 5.453529, 5.467171, 5.481771, 5.49093, 5.491922, 5.482465, 
    5.461075, 5.427461, 5.382823, 5.329916, 5.272722, 5.215748, 5.163129, 
    5.11786, 5.081418, 5.053839, 5.034134, 5.020792, 5.012212, 5.00699, 
    5.004033,
  // momentumX(7,46, 0-49)
    5.000904, 5.001698, 5.003219, 5.005941, 5.01059, 5.018181, 5.030026, 
    5.047634, 5.072513, 5.105799, 5.147814, 5.197673, 5.25313, 5.310821, 
    5.366889, 5.418075, 5.464053, 5.494967, 5.512374, 5.518117, 5.514961, 
    5.509031, 5.500986, 5.493574, 5.486524, 5.481907, 5.480128, 5.480912, 
    5.48242, 5.485212, 5.486995, 5.487328, 5.480935, 5.465807, 5.440713, 
    5.405491, 5.361278, 5.310514, 5.256648, 5.203514, 5.154617, 5.112494, 
    5.078404, 5.052387, 5.033595, 5.020703, 5.01228, 5.007036, 5.003934, 
    5.002227,
  // momentumX(7,47, 0-49)
    5.000479, 5.000916, 5.001769, 5.003335, 5.006079, 5.010685, 5.018091, 
    5.029477, 5.046185, 5.069523, 5.100471, 5.139313, 5.185328, 5.236683, 
    5.29062, 5.344086, 5.395159, 5.436237, 5.466683, 5.48693, 5.498612, 
    5.506318, 5.510494, 5.51297, 5.512695, 5.511067, 5.508265, 5.504123, 
    5.497348, 5.489172, 5.47811, 5.463986, 5.442956, 5.414068, 5.377319, 
    5.333785, 5.285583, 5.235593, 5.186958, 5.142507, 5.104268, 5.07323, 
    5.049392, 5.032015, 5.019961, 5.011981, 5.006932, 5.003879, 5.00212, 
    5.001179,
  // momentumX(7,48, 0-49)
    5.000237, 5.00046, 5.000906, 5.001745, 5.003255, 5.005858, 5.010167, 
    5.017009, 5.027408, 5.04252, 5.063472, 5.091123, 5.125785, 5.16698, 
    5.213346, 5.262811, 5.313305, 5.359091, 5.398305, 5.430139, 5.45493, 
    5.475578, 5.491802, 5.50423, 5.510761, 5.511994, 5.507837, 5.49834, 
    5.482945, 5.46386, 5.440705, 5.414022, 5.381519, 5.343398, 5.300726, 
    5.255343, 5.209594, 5.165942, 5.126526, 5.092831, 5.06552, 5.044494, 
    5.029083, 5.018308, 5.011105, 5.006493, 5.003665, 5.002002, 5.00107, 
    5.000583,
  // momentumX(7,49, 0-49)
    5.000078, 5.000158, 5.000323, 5.000648, 5.001265, 5.002378, 5.004317, 
    5.007565, 5.012781, 5.020815, 5.032668, 5.049388, 5.071904, 5.100811, 
    5.136148, 5.177304, 5.223419, 5.26947, 5.313471, 5.353898, 5.39002, 
    5.424407, 5.454918, 5.480593, 5.49589, 5.500593, 5.494115, 5.476953, 
    5.449314, 5.416775, 5.380487, 5.34278, 5.30167, 5.258408, 5.214767, 
    5.172745, 5.1342, 5.100561, 5.072627, 5.050539, 5.033884, 5.021892, 
    5.013636, 5.008191, 5.004746, 5.002652, 5.001432, 5.00075, 5.000383, 
    5.000201,
  // momentumX(8,0, 0-49)
    5.001369, 5.00236, 5.004135, 5.007111, 5.011874, 5.019187, 5.02997, 
    5.045208, 5.065813, 5.092411, 5.125103, 5.163265, 5.205472, 5.249606, 
    5.293155, 5.333694, 5.369721, 5.397316, 5.416229, 5.42692, 5.430637, 
    5.429839, 5.425939, 5.420931, 5.415915, 5.412307, 5.410614, 5.410615, 
    5.41119, 5.411488, 5.409767, 5.404738, 5.39423, 5.377171, 5.353137, 
    5.322467, 5.286308, 5.246513, 5.205389, 5.165338, 5.128472, 5.096318, 
    5.069674, 5.048647, 5.032804, 5.021383, 5.013495, 5.008281, 5.005001, 
    5.003084,
  // momentumX(8,1, 0-49)
    5.002229, 5.003803, 5.006566, 5.011106, 5.018226, 5.028921, 5.044301, 
    5.065442, 5.093146, 5.127659, 5.168413, 5.213895, 5.261753, 5.309123, 
    5.353121, 5.391528, 5.424201, 5.445468, 5.456513, 5.458668, 5.453891, 
    5.445782, 5.435674, 5.425931, 5.417472, 5.412071, 5.410341, 5.412109, 
    5.416037, 5.421542, 5.426564, 5.429821, 5.428074, 5.419613, 5.403261, 
    5.378569, 5.345982, 5.306887, 5.263489, 5.218513, 5.174774, 5.134702, 
    5.100015, 5.071559, 5.049369, 5.032875, 5.021171, 5.013241, 5.008139, 
    5.005085,
  // momentumX(8,2, 0-49)
    5.003713, 5.006243, 5.010573, 5.017516, 5.028118, 5.043579, 5.065092, 
    5.093582, 5.12938, 5.171907, 5.219525, 5.269629, 5.319023, 5.3645, 
    5.403409, 5.434417, 5.459604, 5.47129, 5.472511, 5.465329, 5.452096, 
    5.437172, 5.421472, 5.407487, 5.395916, 5.388781, 5.386798, 5.389922, 
    5.39677, 5.407083, 5.418703, 5.430604, 5.438771, 5.441057, 5.435635, 
    5.421216, 5.397282, 5.364281, 5.323711, 5.278013, 5.230247, 5.183597, 
    5.140839, 5.103923, 5.073798, 5.050491, 5.033351, 5.021364, 5.013425, 
    5.008539,
  // momentumX(8,3, 0-49)
    5.006076, 5.010056, 5.016683, 5.027022, 5.042336, 5.063916, 5.092799, 
    5.129389, 5.173098, 5.222139, 5.273632, 5.324032, 5.36979, 5.408006, 
    5.436888, 5.456504, 5.471837, 5.472431, 5.463517, 5.447612, 5.427128, 
    5.40682, 5.386859, 5.369648, 5.355633, 5.346969, 5.344492, 5.348353, 
    5.357283, 5.371386, 5.388593, 5.408371, 5.426187, 5.439701, 5.446662, 
    5.445097, 5.433551, 5.411355, 5.378881, 5.337667, 5.290347, 5.24031, 
    5.191145, 5.146004, 5.107107, 5.075537, 5.051323, 5.033752, 5.021726, 
    5.014085,
  // momentumX(8,4, 0-49)
    5.009637, 5.015692, 5.025481, 5.040294, 5.061502, 5.09025, 5.127049, 
    5.171336, 5.221224, 5.273581, 5.324505, 5.370071, 5.407087, 5.433594, 
    5.449055, 5.455122, 5.460109, 5.449643, 5.431532, 5.408463, 5.382619, 
    5.358882, 5.336395, 5.317299, 5.301744, 5.291907, 5.288743, 5.292657, 
    5.302639, 5.319189, 5.340461, 5.366611, 5.392787, 5.416655, 5.435787, 
    5.447778, 5.450466, 5.442185, 5.42209, 5.39045, 5.348847, 5.300132, 
    5.24806, 5.196651, 5.149448, 5.108942, 5.07633, 5.051642, 5.034104, 
    5.022564,
  // momentumX(8,5, 0-49)
    5.01475, 5.023616, 5.037497, 5.057807, 5.085801, 5.12212, 5.166306, 
    5.216456, 5.269265, 5.320505, 5.365861, 5.401783, 5.426079, 5.438101, 
    5.438597, 5.430701, 5.42629, 5.4058, 5.380095, 5.351824, 5.322756, 
    5.297715, 5.274599, 5.255134, 5.239125, 5.228632, 5.224696, 5.228026, 
    5.237998, 5.255537, 5.279135, 5.309788, 5.342454, 5.374955, 5.404862, 
    5.429592, 5.446565, 5.453413, 5.448264, 5.430104, 5.399138, 5.357038, 
    5.306925, 5.252957, 5.199602, 5.15078, 5.109215, 5.07619, 5.051716, 
    5.034968,
  // momentumX(8,6, 0-49)
    5.021751, 5.034218, 5.053062, 5.079626, 5.114713, 5.158042, 5.207815, 
    5.260664, 5.312117, 5.35747, 5.39277, 5.415498, 5.424806, 5.421356, 
    5.406937, 5.385913, 5.373868, 5.3448, 5.313278, 5.281764, 5.251529, 
    5.227237, 5.205383, 5.187147, 5.171925, 5.161469, 5.156841, 5.159067, 
    5.168033, 5.185125, 5.209272, 5.242446, 5.279513, 5.318528, 5.357177, 
    5.392874, 5.422873, 5.444416, 5.454944, 5.452408, 5.435674, 5.404944, 
    5.362053, 5.310448, 5.254735, 5.199829, 5.15, 5.108155, 5.075609, 5.052327,
  // momentumX(8,7, 0-49)
    5.03087, 5.047679, 5.07213, 5.105202, 5.146861, 5.19554, 5.247961, 
    5.299513, 5.345158, 5.38049, 5.402569, 5.410242, 5.403994, 5.385534, 
    5.357308, 5.324667, 5.306974, 5.270771, 5.235045, 5.202008, 5.172415, 
    5.150715, 5.131906, 5.116521, 5.103456, 5.093926, 5.088892, 5.089666, 
    5.096759, 5.112054, 5.135026, 5.168761, 5.208121, 5.251438, 5.296572, 
    5.341026, 5.38205, 5.416742, 5.442186, 5.45566, 5.454984, 5.438967, 
    5.407883, 5.363819, 5.310629, 5.253408, 5.197519, 5.147527, 5.106443, 
    5.075536,
  // momentumX(8,8, 0-49)
    5.042141, 5.063857, 5.094147, 5.13329, 5.180078, 5.231492, 5.282947, 
    5.329145, 5.365218, 5.387711, 5.395039, 5.387403, 5.366355, 5.334259, 
    5.293848, 5.251297, 5.229727, 5.187588, 5.148976, 5.115803, 5.088339, 
    5.070806, 5.056664, 5.045733, 5.036299, 5.028781, 5.023865, 5.023066, 
    5.027584, 5.039847, 5.060001, 5.092403, 5.132013, 5.177479, 5.226856, 
    5.277767, 5.32753, 5.373251, 5.411896, 5.440407, 5.455941, 5.456232, 
    5.440107, 5.408016, 5.362398, 5.307615, 5.249297, 5.193226, 5.14417, 
    5.105097,
  // momentumX(8,9, 0-49)
    5.055322, 5.08219, 5.118004, 5.162039, 5.21173, 5.262723, 5.309602, 
    5.347069, 5.371074, 5.379469, 5.372033, 5.35006, 5.315778, 5.271844, 
    5.22097, 5.170115, 5.145872, 5.098701, 5.058197, 5.025952, 5.0018, 
    4.989735, 4.981704, 4.976761, 4.972498, 4.968266, 4.964252, 4.962024, 
    4.963476, 4.971612, 4.987387, 5.016612, 5.05449, 5.100041, 5.151529, 
    5.206686, 5.262909, 5.317366, 5.367041, 5.408783, 5.439424, 5.456029, 
    5.456311, 5.439203, 5.405454, 5.357993, 5.301782, 5.243008, 5.187781, 
    5.140861,
  // momentumX(8,10, 0-49)
    5.069841, 5.101693, 5.142138, 5.189268, 5.239218, 5.286673, 5.326009, 
    5.352551, 5.363453, 5.357918, 5.336849, 5.30226, 5.256696, 5.202795, 
    5.143048, 5.085224, 5.058656, 5.007109, 4.965445, 4.934928, 4.915015, 
    4.909478, 4.908812, 4.911294, 4.913756, 4.914239, 4.912184, 4.908985, 
    4.907153, 4.910244, 4.920147, 4.944366, 4.97854, 5.022159, 5.07372, 
    5.131052, 5.191589, 5.252552, 5.310984, 5.363772, 5.407672, 5.439425, 
    5.456047, 5.4553, 5.436343, 5.400368, 5.35093, 5.293661, 5.235225, 
    5.181823,
  // momentumX(8,11, 0-49)
    5.084838, 5.121063, 5.164775, 5.212887, 5.260504, 5.301888, 5.331789, 
    5.346568, 5.34467, 5.326456, 5.293612, 5.248514, 5.193708, 5.13161, 
    5.064352, 5.000533, 4.970798, 4.915408, 4.873148, 4.844985, 4.83006, 
    4.831906, 4.839677, 4.850883, 4.861561, 4.868284, 4.869509, 4.866175, 
    4.861197, 4.858579, 4.861226, 4.878594, 4.907023, 4.946648, 4.996276, 
    5.053806, 5.116663, 5.182054, 5.247064, 5.308654, 5.363636, 5.408683, 
    5.44047, 5.45601, 5.453212, 5.431593, 5.392934, 5.341518, 5.283602, 
    5.226091,
  // momentumX(8,12, 0-49)
    5.099267, 5.138888, 5.184268, 5.231308, 5.274516, 5.308251, 5.328059, 
    5.331479, 5.318122, 5.289199, 5.246833, 5.19346, 5.131418, 5.062748, 
    4.989133, 4.919843, 4.884488, 4.825829, 4.783488, 4.758223, 4.748928, 
    4.758839, 4.775925, 4.796943, 4.817178, 4.831673, 4.837736, 4.835538, 
    4.828052, 4.819459, 4.813668, 4.822335, 4.842855, 4.876289, 4.92189, 
    4.977654, 5.040928, 5.108822, 5.178389, 5.246644, 5.310491, 5.366675, 
    5.411796, 5.442484, 5.455814, 5.449941, 5.424872, 5.383087, 5.32959, 
    5.271071,
  // momentumX(8,13, 0-49)
    5.112081, 5.153917, 5.199409, 5.243758, 5.281303, 5.306915, 5.317125, 
    5.310584, 5.287816, 5.250561, 5.201094, 5.141697, 5.07436, 5.000659, 
    4.921747, 4.846888, 4.801401, 4.740222, 4.698379, 4.676562, 4.673483, 
    4.691962, 4.719002, 4.750622, 4.781459, 4.80514, 4.817774, 4.818466, 
    4.809773, 4.795585, 4.780596, 4.77881, 4.789131, 4.813954, 4.853247, 
    4.905177, 4.966969, 5.035536, 5.107794, 5.180731, 5.25133, 5.316455, 
    5.372781, 5.41683, 5.445218, 5.455135, 5.445074, 5.415627, 5.37001, 
    5.313847,
  // momentumX(8,14, 0-49)
    5.122416, 5.165294, 5.209671, 5.250387, 5.28198, 5.300036, 5.302077, 
    5.287667, 5.25795, 5.214927, 5.160814, 5.097618, 5.026911, 4.949761, 
    4.8667, 4.785186, 4.722669, 4.659978, 4.619365, 4.601606, 4.605288, 
    4.632604, 4.669907, 4.712483, 4.754512, 4.788497, 4.809477, 4.815284, 
    4.807504, 4.789055, 4.764913, 4.75128, 4.749103, 4.762674, 4.793109, 
    4.838937, 4.897255, 4.964674, 5.037851, 5.11364, 5.18903, 5.260995, 
    5.326344, 5.381658, 5.423375, 5.448099, 5.453174, 5.437504, 5.402347, 
    5.351675,
  // momentumX(8,15, 0-49)
    5.129766, 5.172712, 5.215269, 5.252206, 5.278469, 5.290407, 5.286373, 
    5.266594, 5.232567, 5.18635, 5.129982, 5.065152, 4.993019, 4.914148, 
    4.828405, 4.73751, 4.64882, 4.585863, 4.547379, 4.534361, 4.545287, 
    4.581367, 4.628794, 4.682116, 4.735318, 4.780255, 4.811194, 4.824649, 
    4.820728, 4.800571, 4.768612, 4.74255, 4.725894, 4.725502, 4.744281, 
    4.781486, 4.83417, 4.898561, 4.970917, 5.047832, 5.126202, 5.203052, 
    5.275322, 5.339731, 5.392716, 5.430585, 5.449921, 5.448276, 5.425073, 
    5.382407,
  // momentumX(8,16, 0-49)
    5.134052, 5.176439, 5.217067, 5.250836, 5.273164, 5.281045, 5.27343, 
    5.250941, 5.215213, 5.16822, 5.111789, 5.047322, 4.975654, 4.896925, 
    4.81037, 4.704902, 4.579583, 4.517775, 4.48243, 4.474857, 4.49339, 
    4.537728, 4.59462, 4.65787, 4.721575, 4.777524, 4.819635, 4.843246, 
    4.846655, 4.828532, 4.791764, 4.754059, 4.721835, 4.705099, 4.70937, 
    4.735244, 4.779961, 4.839344, 4.909132, 4.985513, 5.065176, 5.145107, 
    5.222342, 5.293738, 5.355831, 5.404837, 5.436883, 5.448555, 5.437765, 
    5.404779,
  // momentumX(8,17, 0-49)
    5.13558, 5.177178, 5.216339, 5.248187, 5.268536, 5.274807, 5.266268, 
    5.243672, 5.208608, 5.162899, 5.108179, 5.045659, 4.975985, 4.899038, 
    4.813493, 4.685416, 4.513347, 4.454445, 4.423234, 4.421718, 4.448077, 
    4.499756, 4.565007, 4.636907, 4.70996, 4.776448, 4.830373, 4.866174, 
    4.880282, 4.868591, 4.831599, 4.784774, 4.737452, 4.702971, 4.690291, 
    4.702183, 4.736541, 4.78889, 4.854359, 4.928604, 5.007979, 5.08934, 
    5.169746, 5.246167, 5.315263, 5.37328, 5.416127, 5.43977, 5.440993, 
    5.418493,
  // momentumX(8,18, 0-49)
    5.134904, 5.175833, 5.214426, 5.246045, 5.266733, 5.274041, 5.267223, 
    5.246889, 5.214422, 5.171445, 5.119457, 5.059613, 4.99252, 4.917845, 
    4.833514, 4.673349, 4.446044, 4.392892, 4.366827, 4.371818, 4.406159, 
    4.46414, 4.53652, 4.615712, 4.696862, 4.773158, 4.838974, 4.888155, 
    4.915483, 4.914273, 4.88238, 4.830496, 4.7705, 4.718554, 4.687547, 
    4.683339, 4.705169, 4.748554, 4.808033, 4.878636, 4.956275, 5.037578, 
    5.119546, 5.199218, 5.273369, 5.338331, 5.389959, 5.423878, 5.43611, 
    5.42413,
  // momentumX(8,19, 0-49)
    5.132595, 5.173156, 5.21232, 5.245671, 5.269256, 5.280378, 5.277858, 
    5.261819, 5.23324, 5.193517, 5.144123, 5.086297, 5.020607, 4.946133, 
    4.858912, 4.659686, 4.369835, 4.327592, 4.308208, 4.320153, 4.362873, 
    4.426592, 4.505294, 4.590879, 4.679287, 4.764817, 4.84228, 4.905135, 
    4.946831, 4.958759, 4.936626, 4.884299, 4.815693, 4.74858, 4.699572, 
    4.678265, 4.686046, 4.71891, 4.770968, 4.836618, 4.91126, 4.991214, 
    5.073359, 5.154741, 5.232225, 5.30225, 5.360712, 5.4031, 5.424982, 
    5.422957,
  // momentumX(8,20, 0-49)
    5.126199, 5.16312, 5.199585, 5.231456, 5.255075, 5.268044, 5.269554, 
    5.260229, 5.241733, 5.216325, 5.186499, 5.154742, 5.123319, 5.093983, 
    5.067405, 0, 4.110707, 4.123703, 4.162252, 4.22343, 4.302578, 4.387699, 
    4.480834, 4.576489, 4.673163, 4.767192, 4.854263, 4.927924, 4.980938, 
    5.003913, 4.991771, 4.940973, 4.867107, 4.788014, 4.72289, 4.684924, 
    4.678152, 4.699588, 4.743227, 4.802933, 4.873587, 4.951164, 5.032368, 
    5.114204, 5.193589, 5.267064, 5.330619, 5.379736, 5.409759, 5.416706,
  // momentumX(8,21, 0-49)
    5.123293, 5.160292, 5.19839, 5.233569, 5.261959, 5.280674, 5.288291, 
    5.284894, 5.271763, 5.25098, 5.225037, 5.196559, 5.168098, 5.141923, 
    5.119676, 0, 4.030297, 4.047019, 4.093606, 4.164876, 4.254046, 4.343937, 
    4.441362, 4.540665, 4.641256, 4.74086, 4.835884, 4.920084, 4.985749, 
    5.023064, 5.026696, 4.98524, 4.915319, 4.832731, 4.757448, 4.705839, 
    4.685367, 4.695097, 4.729599, 4.782505, 4.848262, 4.922476, 5.001632, 
    5.082644, 5.162446, 5.237658, 5.304375, 5.358139, 5.394198, 5.408191,
  // momentumX(8,22, 0-49)
    5.121522, 5.158882, 5.19856, 5.236558, 5.268754, 5.291821, 5.30385, 
    5.304541, 5.29497, 5.277183, 5.253765, 5.227507, 5.201188, 5.177412, 
    5.158434, 0, 3.962537, 3.984438, 4.038232, 4.117738, 4.215069, 4.308348, 
    4.409274, 4.511858, 4.616008, 4.720365, 4.821665, 4.913651, 4.988194, 
    5.035557, 5.051208, 5.016985, 4.95165, 4.868662, 4.787441, 4.726087, 
    4.694775, 4.694649, 4.721154, 4.767963, 4.829233, 4.900268, 4.97734, 
    5.057264, 5.136958, 5.2131, 5.281876, 5.338915, 5.379454, 5.398909,
  // momentumX(8,23, 0-49)
    5.120916, 5.158588, 5.199337, 5.239162, 5.273767, 5.299524, 5.314222, 
    5.31733, 5.309831, 5.293787, 5.271873, 5.247006, 5.222109, 5.199984, 
    5.183231, 0, 3.917093, 3.943388, 4.002137, 4.086914, 4.189435, 4.283938, 
    4.386425, 4.49054, 4.59648, 4.703573, 4.808774, 4.905783, 4.986151, 
    5.040359, 5.064946, 5.036311, 4.975649, 4.894337, 4.810658, 4.743364, 
    4.704498, 4.696982, 4.71723, 4.759143, 4.816749, 4.885137, 4.960407, 
    5.039274, 5.118623, 5.195158, 5.265129, 5.324236, 5.367732, 5.390903,
  // momentumX(8,24, 0-49)
    5.121484, 5.15919, 5.200179, 5.240473, 5.275757, 5.302342, 5.317935, 
    5.321938, 5.315293, 5.30006, 5.278937, 5.254865, 5.230805, 5.209631, 
    5.194072, 0, 3.898081, 3.926662, 3.987599, 4.074533, 4.179204, 4.273223, 
    4.375597, 4.479658, 4.58575, 4.69365, 4.800478, 4.89992, 4.983319, 
    5.04135, 5.071414, 5.046269, 4.989053, 4.909707, 4.825484, 4.755218, 
    4.711973, 4.699844, 4.715989, 4.754571, 4.8096, 4.876063, 4.949962, 
    5.027952, 5.106898, 5.183519, 5.254107, 5.31441, 5.359709, 5.385231,
  // momentumX(8,25, 0-49)
    5.12319, 5.160546, 5.200797, 5.240048, 5.274151, 5.299625, 5.314344, 
    5.317798, 5.31093, 5.295742, 5.274842, 5.251086, 5.227356, 5.206459, 
    5.191058, 0, 3.905595, 3.934001, 3.99451, 4.080811, 4.184822, 4.277218, 
    4.378278, 4.481149, 4.586186, 4.693312, 4.799687, 4.89899, 4.982497, 
    5.040989, 5.072271, 5.047817, 4.991623, 4.913149, 4.829183, 4.758409, 
    4.714091, 4.70067, 4.715574, 4.753094, 4.807269, 4.873075, 4.946495, 
    5.024164, 5.102949, 5.179572, 5.250342, 5.311027, 5.356915, 5.383218,
  // momentumX(8,26, 0-49)
    5.125965, 5.16261, 5.201203, 5.237979, 5.269135, 5.291635, 5.303749, 
    5.305204, 5.296997, 5.28103, 5.259737, 5.235774, 5.211836, 5.190529, 
    5.174261, 0, 3.937386, 3.963501, 4.021425, 4.104737, 4.20558, 4.295581, 
    4.394385, 4.495152, 4.598157, 4.703125, 4.807133, 4.903847, 4.984638, 
    5.040278, 5.0684, 5.04177, 4.983876, 4.904703, 4.821317, 4.752176, 
    4.709991, 4.698662, 4.715331, 4.75422, 4.809419, 4.87597, 4.949917, 
    5.027929, 5.106887, 5.183514, 5.254105, 5.314409, 5.359708, 5.385231,
  // momentumX(8,27, 0-49)
    5.129717, 5.165435, 5.201689, 5.23486, 5.261594, 5.279465, 5.287314, 
    5.285252, 5.274403, 5.256595, 5.234052, 5.209174, 5.184377, 5.16194, 
    5.143804, 0, 3.989284, 4.01185, 4.065571, 4.143941, 4.239443, 4.326462, 
    4.422174, 4.519982, 4.619985, 4.72141, 4.821146, 4.912863, 4.98817, 
    5.037752, 5.058598, 5.027196, 4.965382, 4.884583, 4.802653, 4.737598, 
    4.700779, 4.694783, 4.716008, 4.758492, 4.81641, 4.884964, 4.96032, 
    5.03923, 5.118601, 5.195146, 5.265124, 5.324234, 5.36773, 5.390903,
  // momentumX(8,28, 0-49)
    5.134365, 5.169187, 5.202791, 5.231663, 5.252913, 5.264796, 5.266833, 
    5.25964, 5.244601, 5.223562, 5.198596, 5.171845, 5.145388, 5.121049, 
    5.100052, 0, 4.056873, 4.075941, 4.124346, 4.195992, 4.284093, 4.367258, 
    4.458745, 4.55243, 4.648153, 4.744445, 4.837958, 4.922404, 4.989758, 
    5.030591, 5.041007, 5.003144, 4.936561, 4.854705, 4.776264, 4.7182, 
    4.689766, 4.691714, 4.719532, 4.767098, 4.828782, 4.900036, 4.977222, 
    5.057204, 5.136929, 5.213084, 5.281867, 5.338911, 5.379453, 5.398908,
  // momentumX(8,29, 0-49)
    5.139871, 5.174164, 5.205247, 5.229603, 5.244735, 5.249564, 5.244349, 
    5.230343, 5.209353, 5.183419, 5.154596, 5.124834, 5.095839, 5.068839, 
    5.043989, 0, 4.134919, 4.152247, 4.194923, 4.258248, 4.336938, 4.414831, 
    4.500596, 4.588754, 4.67878, 4.768302, 4.853632, 4.928486, 4.985303, 
    5.014688, 5.012098, 4.966738, 4.896005, 4.815494, 4.744064, 4.696627, 
    4.679617, 4.691761, 4.727758, 4.781523, 4.847747, 4.922211, 5.001495, 
    5.082574, 5.16241, 5.23764, 5.304365, 5.358133, 5.394195, 5.408189,
  // momentumX(8,30, 0-49)
    5.149293, 5.187366, 5.220729, 5.245617, 5.259345, 5.260664, 5.249608, 
    5.227057, 5.194283, 5.152627, 5.103288, 5.047123, 4.984291, 4.913467, 
    4.830404, 4.635087, 4.366791, 4.33845, 4.330659, 4.350416, 4.397135, 
    4.457949, 4.533136, 4.614896, 4.700094, 4.78401, 4.861721, 4.926516, 
    4.971288, 4.987126, 4.969789, 4.916682, 4.843794, 4.76844, 4.708371, 
    4.675247, 4.67223, 4.696182, 4.74135, 4.801925, 4.873054, 4.950885, 
    5.032222, 5.114128, 5.19355, 5.267044, 5.330608, 5.37973, 5.409755, 
    5.416704,
  // momentumX(8,31, 0-49)
    5.154108, 5.192601, 5.225134, 5.247748, 5.25784, 5.254495, 5.238242, 
    5.21049, 5.172945, 5.127208, 5.074561, 5.015869, 4.951433, 4.880641, 
    4.801196, 4.644937, 4.432422, 4.392949, 4.379121, 4.393623, 4.43407, 
    4.491832, 4.56249, 4.638905, 4.717442, 4.792549, 4.859183, 4.911111, 
    4.942367, 4.945229, 4.916481, 4.861229, 4.793419, 4.729975, 4.685867, 
    4.669163, 4.680465, 4.715677, 4.769167, 4.835639, 4.910736, 4.990936, 
    5.073214, 5.154664, 5.232185, 5.30223, 5.360701, 5.403094, 5.424978, 
    5.422956,
  // momentumX(8,32, 0-49)
    5.157407, 5.197023, 5.230282, 5.252917, 5.262111, 5.256892, 5.237898, 
    5.206759, 5.165463, 5.115866, 5.059437, 4.997152, 4.929425, 4.855934, 
    4.775219, 4.651386, 4.489683, 4.443143, 4.423618, 4.431955, 4.465497, 
    4.519353, 4.584921, 4.655719, 4.727498, 4.793783, 4.849238, 4.888139, 
    4.905953, 4.896959, 4.860013, 4.806783, 4.748804, 4.70111, 4.675007, 
    4.67511, 4.700132, 4.745621, 4.806382, 4.877728, 4.955783, 5.037313, 
    5.119405, 5.199143, 5.273329, 5.33831, 5.389947, 5.423872, 5.436106, 
    5.424129,
  // momentumX(8,33, 0-49)
    5.158516, 5.199754, 5.23505, 5.259749, 5.270575, 5.266178, 5.24701, 
    5.214706, 5.171402, 5.119178, 5.05975, 4.994316, 4.923507, 4.847308, 
    4.764863, 4.663693, 4.545833, 4.494422, 4.469296, 4.470886, 4.496832, 
    4.54519, 4.604345, 4.668429, 4.732591, 4.78956, 4.833763, 4.860198, 
    4.866086, 4.848289, 4.808124, 4.76158, 4.717298, 4.687345, 4.679305, 
    4.695044, 4.732172, 4.786329, 4.852901, 4.927793, 5.007535, 5.089099, 
    5.169616, 5.246097, 5.315227, 5.37326, 5.416117, 5.439764, 5.44099, 
    5.418491,
  // momentumX(8,34, 0-49)
    5.156674, 5.199654, 5.237898, 5.26634, 5.281066, 5.280095, 5.263408, 
    5.232435, 5.189331, 5.136365, 5.075525, 5.008317, 4.935713, 4.858127, 
    4.77535, 4.688264, 4.605028, 4.550157, 4.519898, 4.514716, 4.532631, 
    4.573838, 4.625031, 4.68093, 4.736253, 4.78332, 4.816595, 4.832085, 
    4.828914, 4.806611, 4.768563, 4.732501, 4.703937, 4.691649, 4.700083, 
    4.72925, 4.776286, 4.837176, 4.907887, 4.984814, 5.064787, 5.144894, 
    5.222227, 5.293676, 5.355797, 5.404819, 5.436873, 5.448549, 5.437762, 
    5.404777,
  // momentumX(8,35, 0-49)
    5.151281, 5.195655, 5.237204, 5.270538, 5.291034, 5.29586, 5.284276, 
    5.257265, 5.216847, 5.165399, 5.10517, 5.038023, 4.965342, 4.888039, 
    4.806555, 4.727874, 4.66922, 4.612257, 4.577751, 4.566242, 4.576077, 
    4.608909, 4.650864, 4.69726, 4.742668, 4.779547, 4.802795, 4.809654, 
    4.800983, 4.778551, 4.746922, 4.72342, 4.710607, 4.714301, 4.736648, 
    4.776581, 4.831155, 4.89677, 4.969879, 5.047243, 5.125873, 5.202868, 
    5.275223, 5.339676, 5.392687, 5.430571, 5.449914, 5.448271, 5.425071, 
    5.382406,
  // momentumX(8,36, 0-49)
    5.142104, 5.187049, 5.231609, 5.270293, 5.297827, 5.310411, 5.306343, 
    5.285905, 5.250766, 5.203276, 5.145887, 5.080808, 5.009852, 4.934427, 
    4.85556, 4.782229, 4.739129, 4.681488, 4.643786, 4.626654, 4.628716, 
    4.652565, 4.684572, 4.720676, 4.75562, 4.782554, 4.797193, 4.798059, 
    4.787327, 4.768233, 4.745573, 4.734941, 4.736442, 4.753576, 4.786968, 
    4.834998, 4.894826, 4.963222, 5.037002, 5.113153, 5.188756, 5.260842, 
    5.326259, 5.381612, 5.423351, 5.448085, 5.453167, 5.4375, 5.402345, 
    5.351675,
  // momentumX(8,37, 0-49)
    5.129393, 5.173698, 5.220318, 5.263993, 5.299031, 5.320687, 5.326133, 
    5.314678, 5.287379, 5.246348, 5.194114, 5.133163, 5.065706, 4.993609, 
    4.918402, 4.849136, 4.814672, 4.757637, 4.717738, 4.695762, 4.690593, 
    4.705426, 4.727391, 4.753076, 4.777669, 4.795451, 4.803186, 4.800547, 
    4.790458, 4.776838, 4.763995, 4.765265, 4.778885, 4.806695, 4.848376, 
    4.902049, 4.965028, 5.034365, 5.107103, 5.18033, 5.251101, 5.316327, 
    5.372707, 5.41679, 5.445196, 5.455124, 5.445068, 5.415625, 5.370009, 
    5.313847,
  // momentumX(8,38, 0-49)
    5.113876, 5.156118, 5.203286, 5.250753, 5.292802, 5.323964, 5.340252, 
    5.339784, 5.322693, 5.290582, 5.245847, 5.191123, 5.128939, 5.06156, 
    4.990949, 4.92551, 4.895123, 4.839703, 4.798448, 4.772382, 4.760661, 
    4.766866, 4.779205, 4.794943, 4.809895, 4.819722, 4.822293, 4.81818, 
    4.810492, 4.803233, 4.799835, 4.811351, 4.83469, 4.870549, 4.918038, 
    4.975163, 5.039362, 5.107861, 5.17781, 5.2463, 5.31029, 5.36656, 
    5.411729, 5.442446, 5.455794, 5.449931, 5.424867, 5.383084, 5.329588, 
    5.27107,
  // momentumX(8,39, 0-49)
    5.096656, 5.135428, 5.181291, 5.230628, 5.278194, 5.318223, 5.345743, 
    5.35758, 5.352668, 5.331766, 5.29685, 5.250499, 5.195425, 5.134211, 
    5.069193, 5.00797, 4.979156, 4.926097, 4.884192, 4.854754, 4.837235, 
    4.835485, 4.838983, 4.845691, 4.852136, 4.855419, 4.85442, 4.850298, 
    4.845923, 4.844999, 4.849974, 4.869821, 4.900551, 4.94209, 4.99318, 
    5.051761, 5.115341, 5.181213, 5.246534, 5.308325, 5.363435, 5.408561, 
    5.440397, 5.455967, 5.453187, 5.43158, 5.392928, 5.341514, 5.283599, 
    5.22609,
  // momentumX(8,40, 0-49)
    5.079001, 5.113148, 5.155824, 5.20466, 5.255383, 5.302495, 5.340465, 
    5.364939, 5.373489, 5.365705, 5.342792, 5.306976, 5.260952, 5.2075, 
    5.149253, 5.093055, 5.064897, 5.0148, 4.972912, 4.940837, 4.918354, 
    4.909531, 4.905233, 4.904131, 4.903456, 4.901661, 4.898442, 4.895254, 
    4.894445, 4.899253, 4.911187, 4.93741, 4.973363, 5.018431, 5.071098, 
    5.129232, 5.190343, 5.251703, 5.310411, 5.363389, 5.407419, 5.439262, 
    5.455943, 5.455236, 5.436306, 5.400346, 5.350918, 5.293653, 5.235221, 
    5.181822,
  // momentumX(8,41, 0-49)
    5.062121, 5.090923, 5.128824, 5.174737, 5.225716, 5.277128, 5.323496, 
    5.359679, 5.381943, 5.388488, 5.379393, 5.356171, 5.321213, 5.27729, 
    5.227234, 5.177218, 5.149961, 5.103456, 5.062327, 5.028457, 5.001982, 
    4.98717, 4.976339, 4.968845, 4.962564, 4.957095, 4.952728, 4.950969, 
    4.953513, 4.963099, 4.980418, 5.011087, 5.050213, 5.096777, 5.149055, 
    5.204819, 5.261506, 5.316321, 5.366274, 5.40823, 5.439034, 5.455762, 
    5.456133, 5.439089, 5.405383, 5.35795, 5.301758, 5.242993, 5.187772, 
    5.140857,
  // momentumX(8,42, 0-49)
    5.046977, 5.07022, 5.102299, 5.143245, 5.191529, 5.243844, 5.29543, 
    5.341003, 5.375879, 5.396879, 5.402698, 5.393766, 5.371802, 5.339299, 
    5.299088, 5.256725, 5.231469, 5.189376, 5.149957, 5.115338, 5.086065, 
    5.066585, 5.050688, 5.038368, 5.028037, 5.02018, 5.015453, 5.015247, 
    5.020588, 5.033757, 5.054786, 5.087964, 5.128242, 5.174273, 5.224139, 
    5.275482, 5.32564, 5.371724, 5.410694, 5.439491, 5.455265, 5.455751, 
    5.439777, 5.407797, 5.36226, 5.307529, 5.249246, 5.193198, 5.144154, 
    5.105088,
  // momentumX(8,43, 0-49)
    5.034163, 5.052107, 5.077977, 5.1126, 5.155713, 5.205489, 5.25843, 
    5.309834, 5.354713, 5.388844, 5.409515, 5.415804, 5.408386, 5.389111, 
    5.360541, 5.327561, 5.306041, 5.269506, 5.233062, 5.199059, 5.168477, 
    5.145934, 5.126657, 5.111196, 5.098354, 5.089241, 5.084676, 5.085835, 
    5.093141, 5.108504, 5.131452, 5.165137, 5.204473, 5.247838, 5.293118, 
    5.337825, 5.379192, 5.41429, 5.440164, 5.454059, 5.453766, 5.438076, 
    5.407258, 5.363396, 5.310354, 5.253236, 5.197416, 5.147466, 5.106408, 
    5.075515,
  // momentumX(8,44, 0-49)
    5.023893, 5.037152, 5.057038, 5.08481, 5.121122, 5.165492, 5.215907, 
    5.268845, 5.319784, 5.364102, 5.398016, 5.419214, 5.427063, 5.422406, 
    5.407182, 5.385447, 5.369846, 5.3404, 5.308588, 5.276946, 5.246899, 
    5.223215, 5.202463, 5.185639, 5.171791, 5.162381, 5.15825, 5.160318, 
    5.168521, 5.184505, 5.207436, 5.239498, 5.275653, 5.314039, 5.352384, 
    5.388091, 5.418369, 5.440388, 5.451512, 5.449613, 5.433495, 5.403317, 
    5.360887, 5.309646, 5.254205, 5.199492, 5.149795, 5.108033, 5.075538, 
    5.052284,
  // momentumX(8,45, 0-49)
    5.016068, 5.025445, 5.040023, 5.06117, 5.090047, 5.127151, 5.171838, 
    5.22204, 5.274341, 5.324514, 5.368355, 5.402508, 5.425014, 5.435463, 
    5.434813, 5.426049, 5.418765, 5.398278, 5.373139, 5.345995, 5.318683, 
    5.296079, 5.275944, 5.259601, 5.246169, 5.237257, 5.233617, 5.23592, 
    5.243749, 5.258614, 5.279437, 5.307597, 5.338169, 5.369109, 5.398049, 
    5.4224, 5.439507, 5.446893, 5.442554, 5.425341, 5.395344, 5.354149, 
    5.304817, 5.251482, 5.198609, 5.150136, 5.108815, 5.075948, 5.051572, 
    5.034879,
  // momentumX(8,46, 0-49)
    5.010371, 5.016713, 5.026895, 5.042174, 5.063859, 5.092983, 5.129908, 
    5.173916, 5.222999, 5.273985, 5.323053, 5.366474, 5.401325, 5.425965, 
    5.440145, 5.44553, 5.448809, 5.439283, 5.423095, 5.402858, 5.380724, 
    5.361625, 5.344312, 5.33029, 5.318596, 5.310812, 5.307542, 5.309251, 
    5.315293, 5.327178, 5.343702, 5.365603, 5.388121, 5.409129, 5.4263, 
    5.437255, 5.439753, 5.431987, 5.41292, 5.382617, 5.342471, 5.295172, 
    5.244368, 5.194016, 5.147643, 5.107752, 5.075573, 5.051174, 5.03382, 
    5.022387,
  // momentumX(8,47, 0-49)
    5.006379, 5.010458, 5.017199, 5.027631, 5.042955, 5.064367, 5.092776, 
    5.128459, 5.170724, 5.217763, 5.2668, 5.314528, 5.357748, 5.393965, 
    5.421778, 5.441412, 5.456867, 5.46001, 5.454927, 5.44398, 5.429455, 
    5.416289, 5.403948, 5.393989, 5.385193, 5.379011, 5.375869, 5.37608, 
    5.378881, 5.385936, 5.396016, 5.409431, 5.421616, 5.430514, 5.434071, 
    5.430398, 5.418005, 5.396079, 5.364757, 5.325294, 5.280035, 5.23211, 
    5.184909, 5.141459, 5.10393, 5.073397, 5.049934, 5.032877, 5.021182, 
    5.013739,
  // momentumX(8,48, 0-49)
    5.003644, 5.006086, 5.010241, 5.016864, 5.02692, 5.041507, 5.061704, 
    5.088339, 5.121694, 5.161249, 5.20556, 5.252367, 5.298956, 5.342635, 
    5.381233, 5.413701, 5.441738, 5.458355, 5.465828, 5.466006, 5.46107, 
    5.455938, 5.450424, 5.446013, 5.441033, 5.436764, 5.433451, 5.431307, 
    5.42953, 5.430123, 5.431936, 5.435133, 5.435347, 5.430807, 5.42, 
    5.401847, 5.375895, 5.342507, 5.302944, 5.259302, 5.21424, 5.17055, 
    5.13068, 5.096348, 5.068379, 5.046762, 5.030877, 5.019772, 5.012416, 
    5.007883,
  // momentumX(8,49, 0-49)
    5.001472, 5.002565, 5.00451, 5.007768, 5.012981, 5.020984, 5.032765, 
    5.049376, 5.071753, 5.100489, 5.135601, 5.176348, 5.22122, 5.268123, 
    5.314735, 5.359285, 5.403051, 5.435205, 5.457379, 5.470873, 5.477746, 
    5.48514, 5.4914, 5.497845, 5.49962, 5.498258, 5.49363, 5.486034, 
    5.474223, 5.463232, 5.452115, 5.442515, 5.428285, 5.40822, 5.38172, 
    5.348891, 5.31062, 5.268536, 5.22482, 5.181884, 5.141978, 5.106841, 
    5.077487, 5.054176, 5.036537, 5.023789, 5.01498, 5.009157, 5.005493, 
    5.003342,
  // momentumX(9,0, 0-49)
    5.013042, 5.019694, 5.029954, 5.044734, 5.064919, 5.091146, 5.123545, 
    5.161498, 5.203522, 5.247341, 5.290179, 5.329203, 5.361989, 5.386886, 
    5.403194, 5.411325, 5.413615, 5.407965, 5.397056, 5.382667, 5.366389, 
    5.350346, 5.335258, 5.322433, 5.312547, 5.306667, 5.305348, 5.308775, 
    5.316498, 5.328191, 5.342663, 5.358954, 5.37482, 5.38847, 5.398046, 
    5.401766, 5.398109, 5.386037, 5.365193, 5.336077, 5.300086, 5.259408, 
    5.216734, 5.174833, 5.136135, 5.102393, 5.074556, 5.052821, 5.03683, 
    5.025922,
  // momentumX(9,1, 0-49)
    5.018539, 5.027684, 5.041417, 5.060682, 5.086233, 5.118349, 5.15655, 
    5.19942, 5.244636, 5.289235, 5.330095, 5.364451, 5.390327, 5.406764, 
    5.413841, 5.412899, 5.408258, 5.395083, 5.37753, 5.357601, 5.33689, 
    5.31798, 5.300873, 5.28678, 5.275898, 5.269395, 5.267859, 5.271605, 
    5.28021, 5.293866, 5.31147, 5.332596, 5.354544, 5.375515, 5.393538, 
    5.406585, 5.412741, 5.410409, 5.398545, 5.376884, 5.346107, 5.307889, 
    5.264752, 5.219728, 5.175877, 5.135812, 5.10137, 5.073483, 5.052285, 
    5.037354,
  // momentumX(9,2, 0-49)
    5.026684, 5.039216, 5.057403, 5.082047, 5.113499, 5.151348, 5.194202, 
    5.239692, 5.284729, 5.326012, 5.360569, 5.386237, 5.401902, 5.407519, 
    5.403984, 5.393466, 5.38223, 5.362339, 5.339471, 5.315671, 5.292365, 
    5.272373, 5.254879, 5.240854, 5.229998, 5.223449, 5.221773, 5.225418, 
    5.234077, 5.248452, 5.26766, 5.291913, 5.318253, 5.345037, 5.370354, 
    5.392126, 5.40825, 5.416761, 5.416035, 5.405025, 5.383495, 5.35221, 
    5.312987, 5.268557, 5.222194, 5.177207, 5.136419, 5.101797, 5.074339, 
    5.054193,
  // momentumX(9,3, 0-49)
    5.037796, 5.054545, 5.077931, 5.108358, 5.145469, 5.18788, 5.233158, 
    5.278073, 5.319133, 5.353187, 5.377922, 5.392138, 5.395739, 5.389587, 
    5.375238, 5.355539, 5.338708, 5.313167, 5.286374, 5.260293, 5.236083, 
    5.216662, 5.200305, 5.187636, 5.177845, 5.171894, 5.170265, 5.173514, 
    5.181518, 5.195473, 5.21482, 5.240509, 5.269487, 5.300368, 5.331426, 
    5.360679, 5.385998, 5.405237, 5.416381, 5.417744, 5.408212, 5.3875, 
    5.356378, 5.316756, 5.271558, 5.224334, 5.17869, 5.137706, 5.103526, 
    5.07722,
  // momentumX(9,4, 0-49)
    5.052035, 5.073641, 5.102532, 5.138441, 5.180034, 5.224841, 5.269492, 
    5.310276, 5.3438, 5.367561, 5.380238, 5.381697, 5.372798, 5.355103, 
    5.330607, 5.30267, 5.281563, 5.251438, 5.221951, 5.194925, 5.171211, 
    5.153751, 5.139843, 5.129701, 5.121983, 5.117336, 5.116074, 5.11881, 
    5.125641, 5.138234, 5.156425, 5.182015, 5.211965, 5.245227, 5.280334, 
    5.31548, 5.34862, 5.37757, 5.400111, 5.414134, 5.417838, 5.409997, 
    5.390258, 5.359409, 5.319504, 5.273733, 5.225988, 5.18022, 5.139762, 
    5.106874,
  // momentumX(9,5, 0-49)
    5.06927, 5.096024, 5.130133, 5.170412, 5.21444, 5.258764, 5.299453, 
    5.332823, 5.356091, 5.367723, 5.367478, 5.356185, 5.335419, 5.307194, 
    5.273708, 5.238726, 5.214715, 5.180921, 5.149723, 5.122785, 5.100636, 
    5.086227, 5.075836, 5.069233, 5.064543, 5.061961, 5.061525, 5.063834, 
    5.069201, 5.079716, 5.095667, 5.119814, 5.149218, 5.18323, 5.220694, 
    5.260019, 5.299302, 5.336403, 5.369049, 5.394906, 5.411742, 5.417627, 
    5.411244, 5.392218, 5.361438, 5.321201, 5.275047, 5.227249, 5.182064, 
    5.142961,
  // momentumX(9,6, 0-49)
    5.088974, 5.120697, 5.159075, 5.201886, 5.245714, 5.28647, 5.320168, 
    5.343662, 5.355105, 5.354039, 5.341181, 5.318075, 5.28674, 5.249392, 
    5.208251, 5.167442, 5.141766, 5.105011, 5.072841, 5.046739, 5.026933, 
    5.016384, 5.01034, 5.008129, 5.007359, 5.007643, 5.008629, 5.010802, 
    5.014644, 5.022597, 5.035425, 5.056958, 5.084433, 5.117664, 5.155847, 
    5.197634, 5.241279, 5.284737, 5.325753, 5.361929, 5.390816, 5.410064, 
    5.417652, 5.412226, 5.393486, 5.362525, 5.321963, 5.275724, 5.22841, 
    5.184418,
  // momentumX(9,7, 0-49)
    5.110209, 5.146196, 5.187303, 5.230341, 5.2712, 5.305634, 5.330105, 
    5.342353, 5.341588, 5.328314, 5.30397, 5.270539, 5.230231, 5.185272, 
    5.137776, 5.092242, 5.065883, 5.026673, 4.994061, 4.969322, 4.952398, 
    4.94629, 4.94522, 4.948102, 4.952066, 4.956038, 4.959166, 4.961686, 
    4.96418, 4.969313, 4.978322, 4.996211, 5.020468, 5.051454, 5.088767, 
    5.131334, 5.177573, 5.225541, 5.273042, 5.317697, 5.356995, 5.388387, 
    5.409444, 5.418111, 5.413079, 5.394205, 5.362855, 5.321998, 5.275874, 
    5.22923,
  // momentumX(9,8, 0-49)
    5.131696, 5.170769, 5.212703, 5.253581, 5.289032, 5.315145, 5.329186, 
    5.329929, 5.317555, 5.293313, 5.25909, 5.217057, 5.16942, 5.118283, 
    5.06558, 5.016235, 4.989789, 4.94848, 4.915803, 4.892795, 4.879127, 
    4.877858, 4.882214, 4.890742, 4.900167, 4.908644, 4.914731, 4.918277, 
    4.919837, 4.922133, 4.926813, 4.940151, 4.959956, 4.987245, 5.022112, 
    5.063804, 5.110915, 5.161597, 5.213713, 5.264927, 5.312754, 5.354599, 
    5.387856, 5.410053, 5.419156, 5.413955, 5.394502, 5.362439, 5.321009, 
    5.274606,
  // momentumX(9,9, 0-49)
    5.152001, 5.192673, 5.233472, 5.270114, 5.29842, 5.315174, 5.318628, 
    5.308538, 5.285864, 5.252336, 5.21005, 5.161165, 5.107756, 5.051719, 
    4.994766, 4.942291, 4.915819, 4.872682, 4.84023, 4.81922, 4.809059, 
    4.812881, 4.822952, 4.837524, 4.85301, 4.866771, 4.876707, 4.882144, 
    4.883457, 4.883184, 4.883249, 4.891264, 4.905428, 4.927546, 4.95835, 
    4.997493, 5.043778, 5.095445, 5.150386, 5.2063, 5.260748, 5.311169, 
    5.354927, 5.389367, 5.412012, 5.420855, 5.414785, 5.39402, 5.360405, 
    5.317352,
  // momentumX(9,10, 0-49)
    5.169785, 5.210491, 5.248452, 5.279398, 5.299693, 5.307023, 5.300615, 
    5.281043, 5.249805, 5.208882, 5.160379, 5.106323, 5.048559, 4.988734, 
    4.928304, 4.873112, 4.845929, 4.801261, 4.769295, 4.750492, 4.743991, 
    4.753007, 4.768904, 4.789725, 4.811697, 4.831421, 4.846126, 4.854508, 
    4.856575, 4.854371, 4.849869, 4.852006, 4.859412, 4.874855, 4.899894, 
    4.934735, 4.978467, 5.029416, 5.085478, 5.144336, 5.203576, 5.260691, 
    5.313084, 5.358071, 5.392953, 5.41521, 5.422825, 5.414724, 5.391241, 
    5.354405,
  // momentumX(9,11, 0-49)
    5.184051, 5.223395, 5.257313, 5.281863, 5.294163, 5.292828, 5.27793, 
    5.25065, 5.212797, 5.166412, 5.113485, 5.055821, 4.994998, 4.932372, 
    4.869107, 4.811265, 4.781673, 4.735917, 4.704734, 4.688303, 4.685516, 
    4.699636, 4.72124, 4.748251, 4.776879, 4.803067, 4.823434, 4.835981, 
    4.840165, 4.837159, 4.828632, 4.824708, 4.824437, 4.831717, 4.849192, 
    4.877854, 4.917208, 4.965708, 5.021219, 5.081358, 5.143673, 5.205681, 
    5.264839, 5.318503, 5.363908, 5.398248, 5.41888, 5.423704, 5.411665, 
    5.383304,
  // momentumX(9,12, 0-49)
    5.194335, 5.231282, 5.260574, 5.278791, 5.28386, 5.275225, 5.253618, 
    5.220604, 5.178126, 5.128154, 5.072487, 5.012671, 4.949991, 4.885493, 
    4.82, 4.759103, 4.724104, 4.677974, 4.647959, 4.634027, 4.634865, 
    4.653734, 4.680614, 4.713413, 4.74852, 4.781399, 4.808202, 4.826231, 
    4.834251, 4.832163, 4.82086, 4.811296, 4.802845, 4.800652, 4.808741, 
    4.829211, 4.862217, 4.906439, 4.959705, 5.019504, 5.083271, 5.148478, 
    5.212607, 5.273064, 5.327098, 5.371778, 5.404087, 5.421196, 5.420952, 
    5.402519,
  // momentumX(9,13, 0-49)
    5.20077, 5.234771, 5.259482, 5.27208, 5.271227, 5.25703, 5.230669, 
    5.19392, 5.148717, 5.09689, 5.04002, 4.97939, 4.916002, 4.850582, 
    4.783556, 4.718486, 4.673654, 4.628222, 4.599886, 4.588519, 4.592689, 
    4.615596, 4.646937, 4.684716, 4.725712, 4.765153, 4.798926, 4.823727, 
    4.837541, 4.838665, 4.826695, 4.812769, 4.796377, 4.783873, 4.780921, 
    4.791139, 4.815689, 4.853671, 4.902922, 4.960753, 5.024401, 5.091208, 
    5.158616, 5.22405, 5.284799, 5.337901, 5.380161, 5.408309, 5.419418, 
    5.411558,
  // momentumX(9,14, 0-49)
    5.204044, 5.235059, 5.255784, 5.26395, 5.258807, 5.240928, 5.211757, 
    5.173126, 5.126891, 5.074712, 5.01796, 4.9577, 4.894693, 4.829371, 
    4.761736, 4.690343, 4.630024, 4.586733, 4.560706, 4.551862, 4.558817, 
    4.584635, 4.619225, 4.660789, 4.706684, 4.75217, 4.793106, 4.82573, 
    4.84728, 4.85427, 4.84457, 4.828547, 4.805531, 4.782758, 4.767636, 
    4.765727, 4.779678, 4.809348, 4.852722, 4.90692, 4.968901, 5.035783, 
    5.104878, 5.173582, 5.2392, 5.2988, 5.349137, 5.386735, 5.408215, 5.410872,
  // momentumX(9,15, 0-49)
    5.205245, 5.233704, 5.251448, 5.256646, 5.248955, 5.229216, 5.198977, 
    5.160035, 5.114126, 5.062756, 5.007135, 4.948183, 4.886503, 4.822322, 
    4.75529, 4.674098, 4.592133, 4.552732, 4.529696, 4.523179, 4.532108, 
    4.559325, 4.595654, 4.639558, 4.689092, 4.739789, 4.787691, 4.828758, 
    4.859601, 4.875039, 4.871017, 4.856003, 4.828897, 4.797172, 4.769747, 
    4.754407, 4.755836, 4.775146, 4.810735, 4.859603, 4.918382, 4.983872, 
    5.053164, 5.123552, 5.192328, 5.2566, 5.31316, 5.358506, 5.389058, 5.40165,
  // momentumX(9,16, 0-49)
    5.205641, 5.232349, 5.248367, 5.25215, 5.243571, 5.223566, 5.193663, 
    5.155571, 5.1109, 5.061044, 5.007129, 4.950017, 4.890282, 4.828084, 
    4.762897, 4.667199, 4.558082, 4.524595, 4.505179, 4.500589, 4.510473, 
    4.537367, 4.573853, 4.618652, 4.670533, 4.725457, 4.779788, 4.82938, 
    4.870381, 4.896234, 4.90115, 4.890569, 4.862889, 4.82492, 4.786451, 
    4.75743, 4.745025, 4.7522, 4.7782, 4.820086, 4.874176, 4.936878, 
    5.004986, 5.075613, 5.145999, 5.21328, 5.274343, 5.325768, 5.363969, 
    5.385563,
  // momentumX(9,17, 0-49)
    5.206429, 5.23244, 5.24809, 5.25195, 5.243927, 5.22491, 5.196322, 
    5.159752, 5.116711, 5.068528, 5.016322, 4.960996, 4.903182, 4.84309, 
    4.780164, 4.665139, 4.525096, 4.499957, 4.484663, 4.481379, 4.491128, 
    4.516054, 4.551351, 4.595904, 4.649085, 4.707342, 4.767391, 4.825082, 
    4.876275, 4.913509, 4.929801, 4.926649, 4.902213, 4.861757, 4.814963, 
    4.77341, 4.746902, 4.740796, 4.755741, 4.789182, 4.837222, 4.895868, 
    4.96155, 5.03114, 5.101774, 5.170614, 5.234653, 5.290627, 5.335063, 
    5.36453,
  // momentumX(9,18, 0-49)
    5.208497, 5.234978, 5.251599, 5.256881, 5.250602, 5.233477, 5.206757, 
    5.171896, 5.13033, 5.083377, 5.032204, 4.977786, 4.920807, 4.861402, 
    4.798707, 4.662005, 4.489505, 4.475817, 4.465091, 4.462282, 4.47091, 
    4.492671, 4.525987, 4.569733, 4.623669, 4.684685, 4.74978, 4.814837, 
    4.875535, 4.924022, 4.952873, 4.959058, 4.941103, 4.902152, 4.850769, 
    4.799243, 4.759669, 4.740109, 4.743153, 4.767068, 4.80796, 4.861491, 
    4.9237, 4.991181, 5.060933, 5.130117, 5.195842, 5.255026, 5.304377, 
    5.340523,
  // momentumX(9,19, 0-49)
    5.212205, 5.240322, 5.25919, 5.267125, 5.263608, 5.249043, 5.224416, 
    5.191014, 5.150217, 5.103388, 5.051769, 4.996344, 4.937584, 4.874966, 
    4.806328, 4.651233, 4.447761, 4.448816, 4.443101, 4.439723, 4.446472, 
    4.464695, 4.496089, 4.539269, 4.594101, 4.657805, 4.727543, 4.799196, 
    4.868299, 4.927033, 4.968306, 4.984324, 4.974784, 4.940611, 4.888542, 
    4.830527, 4.780185, 4.748146, 4.739299, 4.753189, 4.786242, 4.833904, 
    4.891861, 4.956418, 5.024415, 5.092998, 5.159379, 5.220663, 5.273758, 
    5.315415,
  // momentumX(9,20, 0-49)
    5.212728, 5.239095, 5.257136, 5.265122, 5.262591, 5.250175, 5.229265, 
    5.201706, 5.169541, 5.134852, 5.099675, 5.065902, 5.035129, 5.008301, 
    4.984965, 0, 4.281867, 4.296238, 4.319592, 4.349007, 4.384036, 4.42006, 
    4.463272, 4.513869, 4.573604, 4.641306, 4.715052, 4.791258, 4.865699, 
    4.931174, 4.981727, 5.005177, 5.003088, 4.974547, 4.924257, 4.862964, 
    4.804741, 4.762134, 4.742292, 4.746347, 4.771365, 4.812787, 4.866036, 
    4.927151, 4.99281, 5.06013, 5.12641, 5.188928, 5.244792, 5.290888,
  // momentumX(9,21, 0-49)
    5.21802, 5.246518, 5.267158, 5.277958, 5.278198, 5.26831, 5.249588, 
    5.223853, 5.193182, 5.159711, 5.125531, 5.092601, 5.062645, 5.036921, 
    5.015751, 0, 4.280171, 4.286097, 4.301404, 4.32449, 4.355588, 4.38597, 
    4.42638, 4.475754, 4.535542, 4.604822, 4.681754, 4.762756, 4.84341, 
    4.91684, 4.978211, 5.011083, 5.019394, 5.000573, 4.957034, 4.897546, 
    4.835649, 4.785192, 4.75563, 4.750137, 4.766894, 4.801638, 4.849658, 
    4.906757, 4.969437, 5.034751, 5.100053, 5.162745, 5.22009, 5.269087,
  // momentumX(9,22, 0-49)
    5.22302, 5.253256, 5.275841, 5.288589, 5.290601, 5.282212, 5.264708, 
    5.239964, 5.210128, 5.177406, 5.143931, 5.111705, 5.082527, 5.057864, 
    5.038573, 0, 4.278119, 4.278525, 4.288034, 4.306596, 4.335303, 4.361061, 
    4.399333, 4.447818, 4.507654, 4.578084, 4.657235, 4.741405, 4.825919, 
    4.904216, 4.972783, 5.011243, 5.026633, 5.015471, 4.978484, 4.922526, 
    4.859972, 4.804983, 4.768548, 4.755605, 4.765541, 4.794574, 4.838022, 
    4.891535, 4.95148, 5.014856, 5.079045, 5.141546, 5.199745, 5.250741,
  // momentumX(9,23, 0-49)
    5.226744, 5.258028, 5.281734, 5.295559, 5.298512, 5.290893, 5.27401, 
    5.249787, 5.220436, 5.188205, 5.155255, 5.1236, 5.095076, 5.07127, 
    5.053352, 0, 4.279414, 4.276551, 4.281965, 4.297147, 4.32407, 4.345681, 
    4.381749, 4.428933, 4.488155, 4.558842, 4.639098, 4.725091, 4.811872, 
    4.893102, 4.966422, 5.00808, 5.028121, 5.022609, 4.991148, 4.939076, 
    4.877542, 4.820482, 4.779746, 4.76159, 4.766459, 4.791107, 4.830965, 
    4.881619, 4.93934, 5.001071, 5.064211, 5.126318, 5.184858, 5.237008,
  // momentumX(9,24, 0-49)
    5.228496, 5.259939, 5.283836, 5.297881, 5.301076, 5.293717, 5.277114, 
    5.253204, 5.224204, 5.192366, 5.159845, 5.128648, 5.100616, 5.077384, 
    5.060251, 0, 4.283651, 4.279233, 4.282315, 4.295458, 4.321284, 4.339952, 
    4.374256, 4.42016, 4.47849, 4.548845, 4.629343, 4.716074, 4.803885, 
    4.886553, 4.962506, 5.005624, 5.028133, 5.025902, 4.997901, 4.948527, 
    4.888073, 4.830173, 4.787071, 4.765799, 4.767502, 4.789327, 4.826833, 
    4.875592, 4.931826, 4.992456, 5.054884, 5.116711, 5.175456, 5.228333,
  // momentumX(9,25, 0-49)
    5.22796, 5.258594, 5.281716, 5.295139, 5.297939, 5.290426, 5.27388, 
    5.250185, 5.221498, 5.190021, 5.157872, 5.127028, 5.099308, 5.07633, 
    5.059365, 0, 4.289196, 4.284725, 4.287505, 4.300285, 4.325872, 4.343461, 
    4.376945, 4.422066, 4.479642, 4.549365, 4.629392, 4.715792, 4.803343, 
    4.885863, 4.962089, 5.004999, 5.027723, 5.026116, 4.998996, 4.950472, 
    4.89053, 4.832613, 4.789001, 4.766916, 4.767715, 4.788686, 4.825451, 
    4.87359, 4.929327, 4.989579, 5.051758, 5.113479, 5.17228, 5.22539,
  // momentumX(9,26, 0-49)
    5.225247, 5.254143, 5.275551, 5.287515, 5.289261, 5.281141, 5.26438, 
    5.240758, 5.21231, 5.18114, 5.149289, 5.11869, 5.091106, 5.068068, 
    5.050664, 0, 4.295433, 4.292458, 4.29705, 4.311205, 4.33739, 4.355901, 
    4.389616, 4.434559, 4.491645, 4.560555, 4.639478, 4.724538, 4.810594, 
    4.891437, 4.965577, 5.006762, 5.027511, 5.023829, 4.99484, 4.945057, 
    4.88476, 4.827417, 4.78503, 4.764428, 4.766649, 4.788824, 4.826549, 
    4.875436, 4.931742, 4.99241, 5.054859, 5.116698, 5.175449, 5.22833,
  // momentumX(9,27, 0-49)
    5.220861, 5.247246, 5.266091, 5.275759, 5.275703, 5.266364, 5.248924, 
    5.225036, 5.196589, 5.16555, 5.133861, 5.103376, 5.075775, 5.052415, 
    5.034029, 0, 4.302463, 4.302832, 4.311277, 4.328385, 4.355904, 4.377017, 
    4.411754, 4.456905, 4.513578, 4.58136, 4.658477, 4.741166, 4.824496, 
    4.902151, 4.97192, 5.009845, 5.026492, 5.018219, 4.984942, 4.932204, 
    4.871093, 4.815196, 4.775881, 4.759018, 4.764867, 4.790172, 4.830435, 
    4.881328, 4.939181, 5.000987, 5.064165, 5.126294, 5.184847, 5.237001,
  // momentumX(9,28, 0-49)
    5.215629, 5.238973, 5.254549, 5.261092, 5.258357, 5.246945, 5.228058, 
    5.203263, 5.174317, 5.143045, 5.111273, 5.080747, 5.053013, 5.029168, 
    5.009374, 0, 4.311146, 4.317119, 4.331298, 4.35264, 4.382026, 4.406691, 
    4.442622, 4.4878, 4.543655, 4.609676, 4.684156, 4.763472, 4.842965, 
    4.916097, 4.979532, 5.0127, 5.023324, 5.008373, 4.969041, 4.912435, 
    4.850762, 4.797608, 4.763256, 4.75213, 4.763408, 4.793327, 4.837316, 
    4.891145, 4.951268, 5.014741, 5.078983, 5.141513, 5.199726, 5.250731,
  // momentumX(9,29, 0-49)
    5.210575, 5.230656, 5.242446, 5.245065, 5.238635, 5.224026, 5.202578, 
    5.175876, 5.145615, 5.11352, 5.081297, 5.050559, 5.022669, 4.99836, 
    4.977002, 0, 4.32097, 4.335202, 4.357126, 4.384002, 4.415863, 4.444396, 
    4.481161, 4.525657, 4.579839, 4.643129, 4.713893, 4.78861, 4.862862, 
    4.929764, 4.984661, 5.011045, 5.013606, 4.990396, 4.944409, 4.88464, 
    4.824273, 4.776336, 4.749413, 4.746114, 4.764445, 4.80021, 4.84885, 
    4.906308, 4.96919, 5.034617, 5.099981, 5.162707, 5.22007, 5.269075,
  // momentumX(9,30, 0-49)
    5.211185, 5.232265, 5.243868, 5.245254, 5.236584, 5.218601, 5.192334, 
    5.158899, 5.119413, 5.074954, 5.0265, 4.974833, 4.92029, 4.862335, 
    4.799018, 4.650102, 4.46623, 4.474145, 4.474097, 4.474111, 4.482029, 
    4.496277, 4.523712, 4.562758, 4.613616, 4.67399, 4.741224, 4.811243, 
    4.879523, 4.938704, 4.982891, 5.000132, 4.992626, 4.960247, 4.908324, 
    4.847715, 4.791922, 4.752495, 4.735684, 4.742134, 4.768816, 4.811302, 
    4.865192, 4.926679, 4.992549, 5.059987, 5.126332, 5.188886, 5.244769, 
    5.290876,
  // momentumX(9,31, 0-49)
    5.20908, 5.227884, 5.236427, 5.234247, 5.221874, 5.200438, 5.171289, 
    5.135762, 5.095062, 5.050255, 5.002267, 4.951888, 4.899677, 4.845722, 
    4.789222, 4.658228, 4.501397, 4.496706, 4.493328, 4.495354, 4.506206, 
    4.525119, 4.554814, 4.594297, 4.643971, 4.701432, 4.764091, 4.828028, 
    4.888942, 4.939219, 4.972041, 4.980291, 4.964257, 4.925714, 4.87197, 
    4.814879, 4.767239, 4.738547, 4.732779, 4.749048, 4.783735, 4.832435, 
    4.89102, 4.955945, 5.024151, 5.092851, 5.159298, 5.220619, 5.273735, 
    5.315403,
  // momentumX(9,32, 0-49)
    5.209422, 5.227388, 5.234317, 5.229859, 5.214752, 5.190379, 5.15834, 
    5.120173, 5.077215, 5.030576, 4.981167, 4.929723, 4.876769, 4.822464, 
    4.766259, 4.657221, 4.530038, 4.515179, 4.508562, 4.511379, 4.524328, 
    4.547682, 4.579953, 4.620469, 4.669526, 4.724418, 4.782448, 4.839732, 
    4.892161, 4.932154, 4.95264, 4.951416, 4.927637, 4.885253, 4.833202, 
    4.783412, 4.747004, 4.730926, 4.736993, 4.76317, 4.805598, 4.860101, 
    4.922898, 4.990724, 5.060675, 5.129973, 5.195764, 5.254982, 5.304353, 
    5.340511,
  // momentumX(9,33, 0-49)
    5.211784, 5.230331, 5.23714, 5.231805, 5.215128, 5.188638, 5.154125, 
    5.113319, 5.067709, 5.018507, 4.966658, 4.912882, 4.857656, 4.801088, 
    4.742635, 4.653386, 4.555256, 4.532505, 4.522496, 4.524918, 4.538918, 
    4.565711, 4.600144, 4.641606, 4.68998, 4.742125, 4.795075, 4.84495, 
    4.887879, 4.916761, 4.925084, 4.915268, 4.8861, 4.843475, 4.797151, 
    4.758084, 4.735029, 4.73236, 4.75014, 4.785647, 4.835072, 4.894595, 
    4.960809, 5.030715, 5.101532, 5.170478, 5.234578, 5.290584, 5.33504, 
    5.364517,
  // momentumX(9,34, 0-49)
    5.215219, 5.235668, 5.243885, 5.23924, 5.222435, 5.195026, 5.158927, 
    5.11603, 5.067999, 5.016191, 4.961662, 4.905194, 4.847309, 4.788183, 
    4.727444, 4.6529, 4.580625, 4.55162, 4.538008, 4.538926, 4.552721, 
    4.581357, 4.616908, 4.658594, 4.70565, 4.754443, 4.80167, 4.843497, 
    4.87642, 4.894343, 4.89206, 4.875939, 4.844918, 4.806159, 4.769204, 
    4.743195, 4.734305, 4.744707, 4.773262, 4.816971, 4.872271, 4.935742, 
    5.004318, 5.075227, 5.145776, 5.213154, 5.274272, 5.325727, 5.363947, 
    5.38555,
  // momentumX(9,35, 0-49)
    5.218414, 5.241881, 5.252987, 5.250708, 5.235466, 5.208694, 5.172336, 
    5.12841, 5.078754, 5.02491, 4.968103, 4.90927, 4.849085, 4.787934, 
    4.725807, 4.660797, 4.609091, 4.575197, 4.557967, 4.556472, 4.56875, 
    4.597325, 4.632507, 4.673204, 4.717884, 4.762468, 4.803359, 4.83689, 
    4.860095, 4.868361, 4.85827, 4.839107, 4.810142, 4.778883, 4.753745, 
    4.741656, 4.746446, 4.768659, 4.806472, 4.856906, 4.916722, 4.98287, 
    5.052571, 5.123204, 5.192127, 5.256485, 5.313095, 5.358469, 5.389037, 
    5.401639,
  // momentumX(9,36, 0-49)
    5.219895, 5.247176, 5.262488, 5.264244, 5.252396, 5.228087, 5.193159, 
    5.149686, 5.099665, 5.044836, 4.98664, 4.926233, 4.864524, 4.80219, 
    4.739642, 4.680242, 4.642906, 4.605454, 4.584847, 4.580313, 4.589905, 
    4.616549, 4.649711, 4.687962, 4.729007, 4.768494, 4.802673, 4.828212, 
    4.842849, 4.843726, 4.829322, 4.810611, 4.787079, 4.765726, 4.753314, 
    4.754615, 4.771617, 4.803811, 4.849074, 4.904593, 4.967452, 5.034897, 
    5.104344, 5.173264, 5.239013, 5.29869, 5.349073, 5.3867, 5.408195, 
    5.410862,
  // momentumX(9,37, 0-49)
    5.218255, 5.249717, 5.27024, 5.277552, 5.270936, 5.25105, 5.219474, 
    5.178236, 5.129437, 5.075015, 5.016646, 4.955743, 4.893483, 4.830852, 
    4.76865, 4.712382, 4.683611, 4.643882, 4.620321, 4.612436, 4.618487, 
    4.641649, 4.671282, 4.705679, 4.741915, 4.775605, 4.803057, 4.82145, 
    4.829312, 4.825551, 4.810279, 4.794975, 4.779095, 4.768571, 4.768416, 
    4.7816, 4.808813, 4.848932, 4.899767, 4.958707, 5.023099, 5.090394, 
    5.158112, 5.223743, 5.284613, 5.33779, 5.380095, 5.408271, 5.419396, 
    5.411546,
  // momentumX(9,38, 0-49)
    5.212383, 5.247881, 5.274166, 5.288225, 5.288517, 5.274992, 5.248788, 
    5.21174, 5.165967, 5.113562, 5.056436, 4.996264, 4.934503, 4.87243, 
    4.811168, 4.756728, 4.73197, 4.691082, 4.665075, 4.653807, 4.65584, 
    4.674464, 4.699435, 4.72888, 4.759443, 4.786973, 4.808064, 4.820529, 
    4.823663, 4.81791, 4.804527, 4.794577, 4.787253, 4.787226, 4.797941, 
    4.821002, 4.856258, 4.902263, 4.956853, 5.017594, 5.082009, 5.147655, 
    5.212077, 5.272727, 5.326886, 5.371646, 5.404006, 5.421148, 5.420925, 
    5.402503,
  // momentumX(9,39, 0-49)
    5.20167, 5.240501, 5.272511, 5.294001, 5.302503, 5.297089, 5.278226, 
    5.247378, 5.20655, 5.157911, 5.103568, 5.045445, 4.985273, 4.924599, 
    4.864816, 4.811718, 4.787943, 4.746778, 4.718848, 4.70439, 4.702281, 
    4.715828, 4.73548, 4.759322, 4.783782, 4.805178, 4.82057, 4.828451, 
    4.828772, 4.823126, 4.813404, 4.809672, 4.810735, 4.820044, 4.839785, 
    4.870599, 4.911798, 4.96177, 5.018401, 5.079369, 5.142285, 5.204723, 
    5.264188, 5.318067, 5.363621, 5.398062, 5.418763, 5.423631, 5.411623, 
    5.383276,
  // momentumX(9,40, 0-49)
    5.186132, 5.22708, 5.264103, 5.293013, 5.310456, 5.314495, 5.304725, 
    5.282016, 5.248078, 5.205032, 5.155106, 5.100437, 5.043005, 4.984615, 
    4.926899, 4.87519, 4.850765, 4.809989, 4.780656, 4.763356, 4.757268, 
    4.765635, 4.779768, 4.797813, 4.816178, 4.8318, 4.84232, 4.846885, 
    4.845916, 4.841768, 4.836526, 4.838995, 4.847562, 4.864634, 4.891436, 
    4.927948, 4.973135, 5.025293, 5.082327, 5.141959, 5.201804, 5.259393, 
    5.312152, 5.357416, 5.392503, 5.414909, 5.422629, 5.414599, 5.391162, 
    5.354355,
  // momentumX(9,41, 0-49)
    5.166451, 5.207902, 5.248558, 5.28407, 5.310394, 5.324593, 5.325236, 
    5.312375, 5.287194, 5.251593, 5.207793, 5.158082, 5.10465, 5.049539, 
    4.994611, 4.944724, 4.91911, 4.879265, 4.849064, 4.829385, 4.819679, 
    4.823095, 4.831874, 4.844314, 4.856938, 4.867391, 4.873917, 4.876226, 
    4.875024, 4.873092, 4.872416, 4.880478, 4.895287, 4.918398, 4.950332, 
    4.990605, 5.037953, 5.090587, 5.146398, 5.203084, 5.258206, 5.309211, 
    5.353455, 5.388292, 5.41125, 5.42033, 5.414435, 5.393792, 5.360259, 
    5.317256,
  // momentumX(9,42, 0-49)
    5.143857, 5.184021, 5.226386, 5.266863, 5.301079, 5.325276, 5.336976, 
    5.335222, 5.320437, 5.294066, 5.258155, 5.215016, 5.166993, 5.116336, 
    5.06512, 5.017797, 4.99126, 4.952888, 4.922406, 4.90091, 4.888094, 
    4.887012, 4.890862, 4.898168, 4.905657, 4.911681, 4.915056, 4.915931, 
    4.915131, 4.915613, 4.919096, 4.931798, 4.951411, 4.978819, 5.014019, 
    5.056201, 5.103926, 5.155319, 5.208214, 5.260242, 5.308877, 5.35149, 
    5.38544, 5.408236, 5.417833, 5.413025, 5.393868, 5.362019, 5.320735, 
    5.274421,
  // momentumX(9,43, 0-49)
    5.119925, 5.157089, 5.198948, 5.24208, 5.282256, 5.315266, 5.337736, 
    5.347641, 5.344442, 5.32887, 5.302574, 5.267717, 5.226689, 5.18188, 
    5.135561, 5.09184, 5.065246, 5.028996, 4.998917, 4.976262, 4.960958, 
    4.95599, 4.955519, 4.958347, 4.961455, 4.963848, 4.964833, 4.96487, 
    4.964771, 4.967505, 4.974444, 4.990649, 5.013561, 5.043531, 5.080167, 
    5.122412, 5.168684, 5.217022, 5.265179, 5.3107, 5.350989, 5.383418, 
    5.405475, 5.415052, 5.410805, 5.392574, 5.361722, 5.321233, 5.275365, 
    5.228883,
  // momentumX(9,44, 0-49)
    5.096272, 5.129057, 5.168241, 5.211352, 5.254784, 5.29438, 5.326228, 
    5.34737, 5.35621, 5.352563, 5.337418, 5.312571, 5.280278, 5.24296, 
    5.203005, 5.164229, 5.138921, 5.105624, 5.076772, 5.053725, 5.036647, 
    5.028522, 5.024458, 5.023581, 5.023133, 5.022689, 5.021945, 5.021548, 
    5.022201, 5.026792, 5.036315, 5.054803, 5.079486, 5.110286, 5.146511, 
    5.186906, 5.22978, 5.273088, 5.314514, 5.351556, 5.381634, 5.402251, 
    5.411257, 5.407187, 5.389662, 5.359727, 5.319985, 5.274365, 5.22749, 
    5.183779,
  // momentumX(9,45, 0-49)
    5.074281, 5.101814, 5.136524, 5.17699, 5.220571, 5.263685, 5.302406, 
    5.333194, 5.353523, 5.36219, 5.359307, 5.346044, 5.324288, 5.296298, 
    5.264447, 5.232249, 5.209951, 5.180675, 5.154027, 5.131465, 5.113417, 
    5.102954, 5.096113, 5.092372, 5.089212, 5.08668, 5.084756, 5.084169, 
    5.085434, 5.091334, 5.102482, 5.122004, 5.14693, 5.17682, 5.210737, 
    5.247275, 5.284656, 5.320791, 5.353364, 5.379928, 5.39808, 5.405691, 
    5.401236, 5.384155, 5.355194, 5.316544, 5.271692, 5.224903, 5.180446, 
    5.141823,
  // momentumX(9,46, 0-49)
    5.0549, 5.07686, 5.105901, 5.141548, 5.18226, 5.22542, 5.26764, 5.305339, 
    5.335418, 5.355771, 5.36553, 5.365007, 5.355437, 5.338662, 5.316822, 
    5.293051, 5.275785, 5.251806, 5.228491, 5.207395, 5.189259, 5.177374, 
    5.168643, 5.162926, 5.157879, 5.153938, 5.151259, 5.150574, 5.152169, 
    5.158724, 5.17048, 5.189789, 5.213448, 5.240694, 5.270373, 5.30097, 
    5.330666, 5.357411, 5.379015, 5.393284, 5.398237, 5.392398, 5.375129, 
    5.346938, 5.309633, 5.26622, 5.22047, 5.176284, 5.136996, 5.104896,
  // momentumX(9,47, 0-49)
    5.038558, 5.055104, 5.07795, 5.107332, 5.142719, 5.182619, 5.224613, 
    5.265657, 5.302625, 5.332863, 5.354623, 5.367231, 5.371015, 5.367095, 
    5.3571, 5.343633, 5.333583, 5.316318, 5.297566, 5.279008, 5.261748, 
    5.249465, 5.23981, 5.233042, 5.226902, 5.222136, 5.219, 5.218166, 
    5.219665, 5.226124, 5.237422, 5.255292, 5.276211, 5.299119, 5.322676, 
    5.345291, 5.365184, 5.380476, 5.389296, 5.389965, 5.381234, 5.362558, 
    5.334355, 5.298147, 5.256485, 5.212605, 5.169889, 5.131297, 5.098928, 
    5.073874,
  // momentumX(9,48, 0-49)
    5.025191, 5.036808, 5.053524, 5.076003, 5.104483, 5.138533, 5.17689, 
    5.217495, 5.257764, 5.295023, 5.326963, 5.351994, 5.369394, 5.379289, 
    5.382505, 5.380936, 5.380241, 5.371087, 5.358146, 5.343263, 5.327931, 
    5.316406, 5.306894, 5.300048, 5.293569, 5.288468, 5.285032, 5.28385, 
    5.284679, 5.29018, 5.29989, 5.31511, 5.331882, 5.348882, 5.364614, 
    5.377472, 5.385822, 5.388123, 5.38307, 5.369785, 5.348024, 5.318344, 
    5.282197, 5.241826, 5.199984, 5.1595, 5.122818, 5.091662, 5.06691, 
    5.048687,
  // momentumX(9,49, 0-49)
    5.012385, 5.018913, 5.028864, 5.043107, 5.062448, 5.087427, 5.118075, 
    5.153737, 5.193004, 5.233839, 5.273879, 5.31083, 5.342823, 5.368688, 
    5.388059, 5.402215, 5.418763, 5.421006, 5.415788, 5.405649, 5.392869, 
    5.385442, 5.379874, 5.377387, 5.372908, 5.368307, 5.363704, 5.359727, 
    5.355256, 5.355647, 5.359989, 5.371101, 5.38187, 5.390671, 5.395897, 
    5.396035, 5.389802, 5.3763, 5.355184, 5.326793, 5.292233, 5.253324, 
    5.212403, 5.171985, 5.134371, 5.101318, 5.073847, 5.052252, 5.036246, 
    5.025198,
  // momentumX(10,0, 0-49)
    5.063582, 5.085031, 5.112928, 5.146696, 5.184947, 5.225497, 5.265574, 
    5.302221, 5.332746, 5.355133, 5.368267, 5.371976, 5.366912, 5.354355, 
    5.335983, 5.3139, 5.291661, 5.267425, 5.244224, 5.223267, 5.205225, 
    5.190944, 5.179907, 5.172104, 5.167113, 5.164995, 5.165788, 5.169702, 
    5.176876, 5.187829, 5.202584, 5.221438, 5.243492, 5.268015, 5.293913, 
    5.31977, 5.34392, 5.364543, 5.379786, 5.387915, 5.38752, 5.377726, 
    5.358419, 5.3304, 5.295416, 5.256012, 5.215207, 5.176044, 5.141145, 
    5.112394,
  // momentumX(10,1, 0-49)
    5.079928, 5.105417, 5.137311, 5.174423, 5.214681, 5.255301, 5.293159, 
    5.325284, 5.349298, 5.363727, 5.368092, 5.362825, 5.349079, 5.32849, 
    5.302971, 5.274961, 5.249591, 5.22163, 5.19565, 5.1729, 5.153946, 
    5.139993, 5.129792, 5.123188, 5.119247, 5.117973, 5.119292, 5.123413, 
    5.130458, 5.141384, 5.156361, 5.176321, 5.200119, 5.227235, 5.256737, 
    5.287312, 5.31734, 5.344975, 5.368256, 5.385231, 5.394138, 5.393606, 
    5.382902, 5.362143, 5.332445, 5.295923, 5.255486, 5.214435, 5.175961, 
    5.142664,
  // momentumX(10,2, 0-49)
    5.100276, 5.12977, 5.1649, 5.203756, 5.243615, 5.281312, 5.313743, 
    5.338332, 5.35337, 5.358143, 5.352868, 5.338513, 5.316582, 5.288897, 
    5.257421, 5.224789, 5.197577, 5.167107, 5.139554, 5.116156, 5.097363, 
    5.084681, 5.076171, 5.071518, 5.069331, 5.069472, 5.071693, 5.076145, 
    5.082903, 5.093283, 5.107612, 5.127469, 5.151559, 5.179631, 5.210985, 
    5.244498, 5.27869, 5.311812, 5.34193, 5.367047, 5.385226, 5.394764, 
    5.394402, 5.383549, 5.362504, 5.332596, 5.296147, 5.256245, 5.216292, 
    5.179459,
  // momentumX(10,3, 0-49)
    5.123564, 5.156494, 5.193518, 5.232036, 5.268888, 5.30088, 5.325299, 
    5.340286, 5.344973, 5.33944, 5.324524, 5.3016, 5.27236, 5.238668, 
    5.202416, 5.166353, 5.138496, 5.1065, 5.078358, 5.055256, 5.03751, 
    5.026891, 5.020802, 5.018765, 5.018983, 5.021102, 5.024645, 5.029631, 
    5.036055, 5.045497, 5.058444, 5.077137, 5.100204, 5.127726, 5.159303, 
    5.194069, 5.230758, 5.267785, 5.303344, 5.335496, 5.362273, 5.381793, 
    5.39242, 5.392964, 5.382909, 5.362636, 5.33356, 5.298093, 5.259374, 
    5.220767,
  // momentumX(10,4, 0-49)
    5.148277, 5.183551, 5.220681, 5.256588, 5.288019, 5.312116, 5.326862, 
    5.331258, 5.325281, 5.309696, 5.285806, 5.25523, 5.219736, 5.181118, 
    5.141133, 5.102629, 5.075132, 5.042326, 5.01433, 4.99224, 4.976225, 
    4.968293, 4.965206, 4.966337, 4.969534, 4.974173, 4.979482, 4.985287, 
    4.991461, 4.999736, 5.010735, 5.027388, 5.048301, 5.073945, 5.104287, 
    5.138782, 5.176426, 5.215847, 5.255407, 5.293285, 5.327562, 5.356293, 
    5.377622, 5.389924, 5.392003, 5.383332, 5.364291, 5.336296, 5.301751, 
    5.263733,
  // momentumX(10,5, 0-49)
    5.17261, 5.208737, 5.244016, 5.275208, 5.299335, 5.314187, 5.318586, 
    5.31239, 5.29629, 5.271561, 5.239791, 5.202709, 5.162052, 5.119503, 
    5.076645, 5.036462, 5.010109, 4.97695, 4.949606, 4.929027, 4.91522, 
    4.910427, 4.91076, 4.915475, 4.92213, 4.929779, 4.937321, 4.944317, 
    4.950469, 4.957533, 4.96622, 4.980175, 4.998003, 5.020619, 5.048433, 
    5.081285, 5.118479, 5.158883, 5.201038, 5.243255, 5.283694, 5.320426, 
    5.351492, 5.375001, 5.389269, 5.393025, 5.385661, 5.367476, 5.339813, 
    5.305001,
  // momentumX(10,6, 0-49)
    5.194726, 5.230039, 5.261647, 5.286497, 5.302191, 5.307335, 5.301603, 
    5.285583, 5.260492, 5.227921, 5.189589, 5.147222, 5.102467, 5.056863, 
    5.011828, 4.97053, 4.945855, 4.912601, 4.886216, 4.867458, 4.85615, 
    4.854763, 4.858765, 4.867326, 4.877797, 4.888885, 4.899129, 4.907778, 
    4.914294, 4.920318, 4.926564, 4.9374, 4.951415, 4.97002, 4.994144, 
    5.024087, 5.059518, 5.099563, 5.142944, 5.188095, 5.233257, 5.276544, 
    5.315973, 5.349518, 5.375189, 5.391176, 5.396054, 5.389062, 5.370367, 
    5.341236,
  // momentumX(10,7, 0-49)
    5.213053, 5.245964, 5.27248, 5.290026, 5.296961, 5.292734, 5.27777, 
    5.253204, 5.220595, 5.181672, 5.138168, 5.091727, 5.04387, 4.995987, 
    4.949328, 4.907313, 4.88458, 4.851351, 4.826089, 4.809305, 4.800615, 
    4.802724, 4.810457, 4.822952, 4.837451, 4.852314, 4.865723, 4.876563, 
    4.88401, 4.889411, 4.893355, 4.900923, 4.910622, 4.924387, 4.94375, 
    4.969565, 5.001939, 5.040301, 5.083554, 5.130239, 5.178657, 5.226962, 
    5.27318, 5.315236, 5.350972, 5.378225, 5.394969, 5.399563, 5.391072, 
    5.369621,
  // momentumX(10,8, 0-49)
    5.226548, 5.255755, 5.276319, 5.286304, 5.284873, 5.272231, 5.249386, 
    5.217844, 5.179329, 5.135591, 5.088283, 5.038926, 4.98889, 4.939411, 
    4.891582, 4.849094, 4.828224, 4.795094, 4.771032, 4.756248, 4.750131, 
    4.755633, 4.766952, 4.783258, 4.801815, 4.820665, 4.837659, 4.851306, 
    4.860435, 4.865911, 4.868018, 4.872491, 4.877636, 4.885912, 4.899523, 
    4.919997, 4.947987, 4.983297, 5.02504, 5.071846, 5.122056, 5.173835, 
    5.225216, 5.274106, 5.318265, 5.355324, 5.38286, 5.39859, 5.40069, 
    5.388237,
  // momentumX(10,9, 0-49)
    5.234836, 5.259479, 5.273821, 5.276622, 5.26777, 5.248077, 5.218955, 
    5.182111, 5.139313, 5.09224, 5.042422, 4.991228, 4.93987, 4.889423, 
    4.840813, 4.797938, 4.778379, 4.745469, 4.722646, 4.709779, 4.706027, 
    4.714598, 4.729111, 4.748862, 4.77128, 4.794157, 4.815078, 4.832183, 
    4.843925, 4.850475, 4.851599, 4.853556, 4.854271, 4.856665, 4.863659, 
    4.877585, 4.899804, 4.930608, 4.969382, 5.014863, 5.0654, 5.119133, 
    5.17407, 5.228092, 5.27892, 5.324071, 5.360898, 5.386709, 5.399065, 
    5.396215,
  // momentumX(10,10, 0-49)
    5.238247, 5.257951, 5.266341, 5.262815, 5.247848, 5.222678, 5.188955, 
    5.148462, 5.102916, 5.053882, 5.002743, 4.950707, 4.898828, 4.848012, 
    4.798991, 4.755602, 4.736162, 4.703743, 4.682203, 4.671069, 4.66929, 
    4.68035, 4.697388, 4.71993, 4.745744, 4.772466, 4.797513, 4.818703, 
    4.834116, 4.843032, 4.844454, 4.844961, 4.841871, 4.838394, 4.838163, 
    4.844429, 4.859446, 4.88419, 4.918439, 4.961081, 5.01046, 5.064648, 
    5.121579, 5.17908, 5.234825, 5.286284, 5.330706, 5.365195, 5.38696, 
    5.393692,
  // momentumX(10,11, 0-49)
    5.237722, 5.252574, 5.255694, 5.247005, 5.227397, 5.198365, 5.161659, 
    5.119038, 5.072123, 5.022343, 4.970935, 4.918961, 4.86732, 4.81674, 
    4.767717, 4.723385, 4.702055, 4.670654, 4.650481, 4.64079, 4.640394, 
    4.653071, 4.671667, 4.696053, 4.724506, 4.754633, 4.783804, 4.809594, 
    4.829752, 4.842523, 4.845928, 4.846569, 4.840914, 4.832191, 4.824595, 
    4.822354, 4.828823, 4.845907, 4.873978, 4.912177, 4.958867, 5.012014, 
    5.069425, 5.128822, 5.187816, 5.243847, 5.294146, 5.335773, 5.365799, 
    5.381611,
  // momentumX(10,12, 0-49)
    5.234626, 5.245103, 5.243909, 5.231354, 5.20858, 5.177192, 5.138937, 
    5.095491, 5.048359, 4.998839, 4.948044, 4.896914, 4.84622, 4.796515, 
    4.748018, 4.701878, 4.675796, 4.646248, 4.627597, 4.618956, 4.619151, 
    4.632289, 4.651206, 4.676237, 4.706321, 4.739155, 4.772195, 4.802876, 
    4.828703, 4.846828, 4.854155, 4.856939, 4.85062, 4.838054, 4.82369, 
    4.812641, 4.809513, 4.817426, 4.837632, 4.869717, 4.912129, 4.962729, 
    5.019142, 5.078934, 5.139617, 5.198605, 5.253157, 5.300396, 5.33741, 
    5.361478,
  // momentumX(10,13, 0-49)
    5.230535, 5.237388, 5.232965, 5.21782, 5.193212, 5.160748, 5.122097, 
    5.078829, 5.032333, 4.983805, 4.934273, 4.884608, 4.835494, 4.787343, 
    4.740097, 4.690714, 4.656355, 4.629813, 4.612917, 4.604844, 4.60468, 
    4.616896, 4.634736, 4.65907, 4.689609, 4.724247, 4.760649, 4.796208, 
    4.828288, 4.853024, 4.866192, 4.873289, 4.868722, 4.854521, 4.834921, 
    4.81561, 4.802438, 4.8, 4.810771, 4.835072, 4.871596, 4.918133, 4.972108, 
    5.030878, 5.091822, 5.152305, 5.209641, 5.261067, 5.303789, 5.335109,
  // momentumX(10,14, 0-49)
    5.22699, 5.231134, 5.224566, 5.207964, 5.182598, 5.150006, 5.111754, 
    5.069297, 5.023933, 4.976803, 4.928903, 4.881094, 4.834053, 4.788131, 
    4.743088, 4.688396, 4.642111, 4.619964, 4.605116, 4.597078, 4.595531, 
    4.605345, 4.620689, 4.643006, 4.672795, 4.708239, 4.747289, 4.787376, 
    4.82584, 4.857959, 4.878545, 4.891905, 4.89165, 4.878604, 4.856218, 
    4.830238, 4.807499, 4.794166, 4.79429, 4.80929, 4.838372, 4.879369, 
    4.929523, 4.985952, 5.04586, 5.106551, 5.16538, 5.219721, 5.266939, 
    5.304432,
  // momentumX(10,15, 0-49)
    5.225293, 5.227697, 5.219958, 5.202792, 5.177416, 5.145269, 5.107808, 
    5.066401, 5.02229, 4.976607, 4.930377, 4.88452, 4.839792, 4.79663, 
    4.75483, 4.69235, 4.631154, 4.614925, 4.602443, 4.593904, 4.58998, 
    4.595966, 4.607544, 4.62669, 4.65465, 4.689934, 4.730808, 4.7748, 
    4.819294, 4.85896, 4.887938, 4.908922, 4.915213, 4.906217, 4.884106, 
    4.854033, 4.823288, 4.799448, 4.788349, 4.792909, 4.813193, 4.847295, 
    4.892347, 4.94524, 5.002972, 5.062758, 5.12198, 5.17813, 5.228736, 
    5.271329,
  // momentumX(10,16, 0-49)
    5.226336, 5.227925, 5.219817, 5.202703, 5.177724, 5.146221, 5.109568, 
    5.06908, 5.025991, 4.981462, 4.936589, 4.892404, 4.84983, 4.809532, 
    4.771629, 4.699264, 4.621652, 4.61295, 4.603134, 4.593575, 4.586397, 
    4.587306, 4.594104, 4.609207, 4.634496, 4.668808, 4.710706, 4.757823, 
    4.807619, 4.854417, 4.892068, 4.921228, 4.935552, 4.933044, 4.914313, 
    4.883314, 4.847099, 4.81419, 4.792173, 4.785765, 4.796284, 4.822381, 
    4.861237, 4.909564, 4.964163, 5.022121, 5.08082, 5.137845, 5.190862, 
    5.237532,
  // momentumX(10,17, 0-49)
    5.230514, 5.23212, 5.224253, 5.207549, 5.183083, 5.152126, 5.116007, 
    5.076031, 5.033445, 4.989463, 4.945265, 4.902009, 4.860803, 4.822589, 
    4.787977, 4.705591, 4.612271, 4.612747, 4.605839, 4.594719, 4.583512, 
    4.578328, 4.579618, 4.590136, 4.612224, 4.645008, 4.687278, 4.736743, 
    4.790919, 4.844021, 4.890014, 4.927098, 4.949994, 4.955523, 4.94271, 
    4.913936, 4.875333, 4.835699, 4.804019, 4.7869, 4.787251, 4.804621, 
    4.836472, 4.879438, 4.930146, 4.985555, 5.04301, 5.100143, 5.154733, 
    5.204546,
  // momentumX(10,18, 0-49)
    5.237718, 5.240082, 5.232924, 5.216834, 5.19283, 5.162156, 5.126127, 
    5.086053, 5.043212, 4.998859, 4.954231, 4.910549, 4.86899, 4.830619, 
    4.796376, 4.707914, 4.602833, 4.613844, 4.60993, 4.59652, 4.580455, 
    4.568354, 4.563672, 4.569397, 4.588124, 4.619167, 4.66143, 4.712628, 
    4.770273, 4.82866, 4.882247, 4.92637, 4.957467, 4.971514, 4.966166, 
    4.942143, 4.904187, 4.860658, 4.821369, 4.794617, 4.785073, 4.793501, 
    4.817908, 4.85501, 4.901318, 4.953671, 5.009349, 5.066003, 5.121474, 
    5.173612,
  // momentumX(10,19, 0-49)
    5.247415, 5.251267, 5.245289, 5.230013, 5.20642, 5.175728, 5.139245, 
    5.098292, 5.054173, 5.008155, 4.961453, 4.915181, 4.870294, 4.827582, 
    4.788054, 4.702839, 4.595904, 4.617163, 4.615731, 4.598713, 4.576507, 
    4.556717, 4.545831, 4.546948, 4.562612, 4.592149, 4.634409, 4.687026, 
    4.747424, 4.810097, 4.870316, 4.920206, 4.958426, 4.980475, 4.982996, 
    4.965231, 4.930353, 4.885727, 4.841322, 4.806689, 4.788195, 4.788025, 
    4.80498, 4.836047, 4.87772, 4.926739, 4.980312, 5.036072, 5.091892, 
    5.14567,
  // momentumX(10,20, 0-49)
    5.253863, 5.255918, 5.248505, 5.232355, 5.208736, 5.179231, 5.145556, 
    5.109469, 5.072702, 5.036943, 5.003791, 4.974656, 4.950539, 4.931577, 
    4.916345, 0, 4.529047, 4.533604, 4.533447, 4.529254, 4.524078, 4.517531, 
    4.516744, 4.524277, 4.543463, 4.574782, 4.617994, 4.671397, 4.732827, 
    4.797443, 4.86176, 4.91475, 4.957507, 4.985386, 4.994432, 4.982762, 
    4.952068, 4.908407, 4.861261, 4.820816, 4.794822, 4.786893, 4.796811, 
    4.82201, 4.859082, 4.904712, 4.956047, 5.010677, 5.066474, 5.121367,
  // momentumX(10,21, 0-49)
    5.263675, 5.267076, 5.260616, 5.245088, 5.221847, 5.192562, 5.159019, 
    5.122997, 5.086214, 5.050299, 5.016766, 4.986938, 4.961788, 4.941614, 
    4.925509, 0, 4.57267, 4.567389, 4.555607, 4.539651, 4.524162, 4.505689, 
    4.496675, 4.498558, 4.514233, 4.543977, 4.587254, 4.642064, 4.705884, 
    4.773979, 4.843802, 4.901035, 4.949372, 4.984136, 5.000959, 4.997036, 
    4.972662, 4.932421, 4.884916, 4.840544, 4.808241, 4.793121, 4.796153, 
    4.815408, 4.847692, 4.889668, 4.938398, 4.991401, 5.046501, 5.101614,
  // momentumX(10,22, 0-49)
    5.271476, 5.27575, 5.269802, 5.254496, 5.231293, 5.201962, 5.168361, 
    5.132299, 5.095483, 5.059496, 5.025783, 4.995612, 4.969961, 4.949296, 
    4.933185, 0, 4.606127, 4.593786, 4.574115, 4.550414, 4.528358, 4.500781, 
    4.48548, 4.482813, 4.495416, 4.523509, 4.566337, 4.621633, 4.686522, 
    4.756358, 4.829571, 4.888551, 4.939791, 4.978797, 5.001094, 5.003343, 
    4.984809, 4.94875, 4.902673, 4.85667, 4.820312, 4.799883, 4.797452, 
    4.8118, 4.840026, 4.878856, 4.925291, 4.976785, 5.031116, 5.086174,
  // momentumX(10,23, 0-49)
    5.276399, 5.281113, 5.275375, 5.260115, 5.236866, 5.207469, 5.173829, 
    5.13778, 5.101011, 5.065071, 5.031356, 5.001098, 4.975291, 4.954518, 
    4.93868, 0, 4.630615, 4.613832, 4.58922, 4.560673, 4.534565, 4.500163, 
    4.480029, 4.473634, 4.483511, 4.509951, 4.552076, 4.607405, 4.672744, 
    4.743471, 4.818842, 4.878325, 4.930957, 4.972464, 4.998406, 5.005173, 
    4.991349, 4.959182, 4.915194, 4.868976, 4.830346, 4.80637, 4.800004, 
    4.810667, 4.83577, 4.87212, 4.916699, 4.966904, 5.020463, 5.075243,
  // momentumX(10,24, 0-49)
    5.277895, 5.282643, 5.276915, 5.261662, 5.238444, 5.20912, 5.175599, 
    5.139707, 5.103124, 5.067368, 5.033813, 5.003671, 4.977938, 4.957258, 
    4.941692, 0, 4.644578, 4.625749, 4.598795, 4.567974, 4.540061, 4.501756, 
    4.478832, 4.470163, 4.478271, 4.503554, 4.545105, 4.600323, 4.665806, 
    4.736924, 4.813501, 4.87292, 4.926011, 4.96866, 4.996484, 5.005741, 
    4.994654, 4.964887, 4.922336, 4.876217, 4.836404, 4.810391, 4.801668, 
    4.810068, 4.83323, 4.868037, 4.911464, 4.96088, 5.013984, 5.068623,
  // momentumX(10,25, 0-49)
    5.275751, 5.280137, 5.274252, 5.259029, 5.235986, 5.20693, 5.173734, 
    5.138188, 5.10195, 5.066529, 5.033287, 5.003433, 4.977952, 4.957484, 
    4.942075, 0, 4.646362, 4.627713, 4.600918, 4.57033, 4.542782, 4.504051, 
    4.480865, 4.47187, 4.479598, 4.504527, 4.545787, 4.600784, 4.666057, 
    4.736995, 4.813643, 4.872583, 4.925354, 4.967914, 4.995914, 5.005612, 
    4.995152, 4.966033, 4.923948, 4.877962, 4.837917, 4.81139, 4.802017, 
    4.809758, 4.832334, 4.866657, 4.909718, 4.958877, 5.011829, 5.066416,
  // momentumX(10,26, 0-49)
    5.270087, 5.273705, 5.267471, 5.252261, 5.229498, 5.200881, 5.168194, 
    5.133167, 5.097431, 5.062489, 5.029718, 5.00033, 4.975293, 4.955161, 
    4.939804, 0, 4.636261, 4.619933, 4.595723, 4.567776, 4.542617, 4.506954, 
    4.486037, 4.478699, 4.487489, 4.512912, 4.554196, 4.60886, 4.67358, 
    4.743774, 4.819333, 4.877504, 4.92928, 4.970582, 4.997083, 5.005145, 
    4.993102, 4.962729, 4.919972, 4.874004, 4.834575, 4.809024, 4.800726, 
    4.809459, 4.832855, 4.867812, 4.911335, 4.960805, 5.013942, 5.0686,
  // momentumX(10,27, 0-49)
    5.261351, 5.26376, 5.256897, 5.241565, 5.219057, 5.190928, 5.158837, 
    5.124437, 5.089321, 5.054998, 5.022872, 4.994169, 4.969829, 4.950259, 
    4.934984, 0, 4.616155, 4.604306, 4.585077, 4.56209, 4.541208, 4.511642, 
    4.495096, 4.490992, 4.501941, 4.528447, 4.569895, 4.624023, 4.687788, 
    4.756649, 4.829976, 4.887001, 4.937045, 4.975907, 4.999275, 5.003732, 
    4.988097, 4.954829, 4.910524, 4.864675, 4.826832, 4.803771, 4.798227, 
    4.809523, 4.835066, 4.871701, 4.916456, 4.966763, 5.020384, 5.0752,
  // momentumX(10,28, 0-49)
    5.250287, 5.251001, 5.243098, 5.227319, 5.204828, 5.177031, 5.145455, 
    5.111665, 5.077218, 5.043633, 5.012346, 4.984618, 4.961354, 4.942771, 
    4.927911, 0, 4.589266, 4.58401, 4.572131, 4.556344, 4.541521, 4.520256, 
    4.509414, 4.509357, 4.5229, 4.55061, 4.592104, 4.645408, 4.707838, 
    4.774844, 4.844988, 4.900376, 4.947849, 4.983022, 5.001625, 5.000618, 
    4.979618, 4.942165, 4.895842, 4.850533, 4.815399, 4.796301, 4.795027, 
    4.81025, 4.839077, 4.87829, 4.924963, 4.976596, 5.031007, 5.086114,
  // momentumX(10,29, 0-49)
    5.237892, 5.236384, 5.226872, 5.210082, 5.187092, 5.159198, 5.127821, 
    5.094449, 5.060609, 5.027836, 4.997607, 4.971239, 4.949625, 4.9328, 
    4.919292, 0, 4.557674, 4.560971, 4.558987, 4.552932, 4.546215, 4.534846, 
    4.530406, 4.534475, 4.550333, 4.578779, 4.61976, 4.671615, 4.73202, 
    4.796323, 4.862085, 4.914719, 4.958258, 4.988181, 5.000409, 4.992544, 
    4.965331, 4.923674, 4.876193, 4.832937, 4.80229, 4.788859, 4.793301, 
    4.813599, 4.846585, 4.889009, 4.938014, 4.991178, 5.046374, 5.101542,
  // momentumX(10,30, 0-49)
    5.229731, 5.229138, 5.220243, 5.203627, 5.180113, 5.150661, 5.116294, 
    5.078084, 5.037141, 4.994608, 4.951617, 4.909244, 4.868432, 4.829989, 
    4.794954, 4.714292, 4.616234, 4.637926, 4.637839, 4.622587, 4.602194, 
    4.580849, 4.568728, 4.568097, 4.581463, 4.608438, 4.648096, 4.698241, 
    4.756376, 4.817419, 4.877771, 4.926244, 4.964109, 4.986963, 4.99125, 
    4.975613, 4.942276, 4.897612, 4.851018, 4.812195, 4.788252, 4.782269, 
    4.793753, 4.820078, 4.857902, 4.904008, 4.955632, 5.010437, 5.066337, 
    5.121289,
  // momentumX(10,31, 0-49)
    5.219232, 5.216277, 5.205369, 5.187213, 5.162733, 5.132943, 5.098883, 
    5.061612, 5.022202, 4.98176, 4.94143, 4.902367, 4.865702, 4.832438, 
    4.803414, 4.719196, 4.623185, 4.63613, 4.634095, 4.622359, 4.607735, 
    4.594142, 4.588014, 4.591664, 4.607731, 4.635858, 4.675278, 4.723969, 
    4.779628, 4.836938, 4.891286, 4.934981, 4.966794, 4.982536, 4.979336, 
    4.957036, 4.91935, 4.873874, 4.830328, 4.797622, 4.781393, 4.783288, 
    4.801867, 4.834084, 4.87652, 4.926019, 4.979887, 5.035825, 5.091748, 
    5.145588,
  // momentumX(10,32, 0-49)
    5.212204, 5.207666, 5.195166, 5.175536, 5.149817, 5.119109, 5.084501, 
    5.047058, 5.007833, 4.967883, 4.928288, 4.890134, 4.854459, 4.822115, 
    4.793561, 4.715725, 4.631017, 4.635134, 4.631091, 4.622012, 4.61214, 
    4.605616, 4.605232, 4.613331, 4.632458, 4.662114, 4.70151, 4.748676, 
    4.801376, 4.854101, 4.901446, 4.939006, 4.963384, 4.970959, 4.959958, 
    4.931739, 4.891537, 4.847791, 4.809901, 4.785426, 4.77831, 4.788849, 
    4.814866, 4.853093, 4.900144, 4.952962, 5.008929, 5.065755, 5.121329, 
    5.173527,
  // momentumX(10,33, 0-49)
    5.20914, 5.203825, 5.190194, 5.169207, 5.142048, 5.109946, 5.074082, 
    5.035568, 4.995455, 4.954757, 4.914469, 4.875549, 4.838848, 4.804925, 
    4.77372, 4.706617, 4.637273, 4.633828, 4.628059, 4.621222, 4.615577, 
    4.615524, 4.620589, 4.633079, 4.655277, 4.686444, 4.725629, 4.770813, 
    4.819751, 4.866857, 4.906264, 4.936515, 4.952563, 4.951732, 4.933675, 
    4.901386, 4.861358, 4.822259, 4.792506, 4.777924, 4.780762, 4.800201, 
    4.83359, 4.877619, 4.929025, 4.984875, 5.042601, 5.0999, 5.154591, 
    5.204463,
  // momentumX(10,34, 0-49)
    5.210141, 5.204962, 5.190825, 5.168797, 5.140215, 5.106468, 5.068875, 
    5.028635, 4.986836, 4.944474, 4.902484, 4.861712, 4.82285, 4.786231, 
    4.751455, 4.695054, 4.642087, 4.632432, 4.625143, 4.620174, 4.618269, 
    4.623944, 4.634017, 4.650625, 4.67562, 4.707963, 4.746448, 4.788954, 
    4.833173, 4.873645, 4.904438, 4.926645, 4.934232, 4.925783, 4.902545, 
    4.868981, 4.83229, 4.800661, 4.780991, 4.77725, 4.790213, 4.818267, 
    4.858552, 4.907861, 4.963102, 5.021472, 5.080428, 5.137609, 5.190722, 
    5.237449,
  // momentumX(10,35, 0-49)
    5.214813, 5.2108, 5.196992, 5.174516, 5.144845, 5.109542, 5.070085, 
    5.0278, 4.983854, 4.939272, 4.894969, 4.851746, 4.810218, 4.770653, 
    4.732632, 4.684653, 4.646751, 4.632051, 4.62333, 4.619743, 4.620919, 
    4.631336, 4.64574, 4.665937, 4.693183, 4.726111, 4.763205, 4.802227, 
    4.84081, 4.873873, 4.895854, 4.909962, 4.909899, 4.895682, 4.870054, 
    4.838493, 4.808202, 4.78625, 4.777755, 4.784982, 4.807583, 4.843489, 
    4.889846, 4.943633, 5.00196, 5.062129, 5.121593, 5.177893, 5.228593, 
    5.271242,
  // momentumX(10,36, 0-49)
    5.222264, 5.220515, 5.208066, 5.186024, 5.155957, 5.119577, 5.078528, 
    5.03429, 4.988141, 4.941181, 4.894366, 4.848512, 4.804265, 4.76197, 
    4.721433, 4.679046, 4.653185, 4.63448, 4.62433, 4.621491, 4.624862, 
    4.638769, 4.656545, 4.67952, 4.708213, 4.740936, 4.775853, 4.810642, 
    4.842913, 4.868268, 4.881892, 4.888682, 4.882713, 4.865387, 4.840581, 
    4.814148, 4.792623, 4.781571, 4.784374, 4.801928, 4.833148, 4.875787, 
    4.927128, 4.984381, 5.044846, 5.105902, 5.164972, 5.219464, 5.266778, 
    5.30433,
  // momentumX(10,37, 0-49)
    5.231169, 5.232775, 5.222847, 5.202373, 5.172933, 5.13634, 5.094387, 
    5.048704, 5.000711, 4.951622, 4.902481, 4.854186, 4.807487, 4.762895, 
    4.720541, 4.681284, 4.663596, 4.641848, 4.63024, 4.627433, 4.631958, 
    4.647927, 4.667863, 4.692542, 4.721674, 4.753293, 4.785275, 4.815282, 
    4.840997, 4.858955, 4.865395, 4.866431, 4.85696, 4.839487, 4.818485, 
    4.799541, 4.78807, 4.788061, 4.801427, 4.82809, 4.86656, 4.914594, 
    4.969669, 5.029223, 5.090712, 5.15157, 5.209159, 5.260755, 5.303586, 
    5.334973,
  // momentumX(10,38, 0-49)
    5.239892, 5.24584, 5.239644, 5.222045, 5.194521, 5.158906, 5.117092, 
    5.070849, 5.021742, 4.971128, 4.920183, 4.869933, 4.821266, 4.774899, 
    4.73128, 4.693408, 4.680095, 4.656179, 4.643091, 4.639637, 4.644267, 
    4.660845, 4.6816, 4.706756, 4.735232, 4.764845, 4.793278, 4.818267, 
    4.837685, 4.849177, 4.850168, 4.847516, 4.837119, 4.822165, 4.80716, 
    4.796963, 4.795705, 4.805967, 4.828554, 4.862772, 4.906951, 4.958941, 
    5.016412, 5.076992, 5.138256, 5.197663, 5.252513, 5.29996, 5.337116, 
    5.361272,
  // momentumX(10,39, 0-49)
    5.246655, 5.257724, 5.256416, 5.243073, 5.218928, 5.18572, 5.145367, 
    5.099737, 5.050538, 4.999286, 4.947315, 4.895807, 4.845814, 4.798248, 
    4.753822, 4.71631, 4.704317, 4.678978, 4.664438, 4.659803, 4.663629, 
    4.679513, 4.699796, 4.724214, 4.750978, 4.777809, 4.802306, 4.822383, 
    4.83622, 4.842612, 4.840141, 4.835948, 4.826879, 4.816355, 4.808491, 
    4.8072, 4.815392, 4.83454, 4.864683, 4.904767, 4.953069, 5.007549, 
    5.066037, 5.126289, 5.185953, 5.242501, 5.293189, 5.335102, 5.365329, 
    5.381271,
  // momentumX(10,40, 0-49)
    5.249744, 5.266394, 5.270947, 5.263197, 5.243958, 5.214726, 5.177338, 
    5.133704, 5.085651, 5.034855, 4.982824, 4.930913, 4.880349, 4.832219, 
    4.787439, 4.749863, 4.737173, 4.711016, 4.69513, 4.68898, 4.691325, 
    4.705497, 4.724216, 4.746839, 4.771021, 4.794501, 4.81493, 4.830498, 
    4.839759, 4.842586, 4.838536, 4.834641, 4.828501, 4.823401, 4.822832, 
    4.829747, 4.846045, 4.872379, 4.908298, 4.952549, 5.003408, 5.058919, 
    5.117007, 5.175501, 5.232083, 5.284229, 5.329195, 5.364105, 5.386174, 
    5.393111,
  // momentumX(10,41, 0-49)
    5.247719, 5.269979, 5.281053, 5.280043, 5.267168, 5.243511, 5.210688, 
    5.170568, 5.125053, 5.075967, 5.024994, 4.973671, 4.923398, 4.875422, 
    4.830817, 4.79321, 4.778804, 4.752316, 4.735268, 4.727466, 4.727908, 
    4.739669, 4.756018, 4.776052, 4.797035, 4.816849, 4.833313, 4.844961, 
    4.85074, 4.851439, 4.847338, 4.845059, 4.842711, 4.843216, 4.849365, 
    4.863264, 4.886032, 4.917758, 4.95768, 5.004436, 5.056305, 5.111372, 
    5.167601, 5.222831, 5.274746, 5.320846, 5.358463, 5.384906, 5.397736, 
    5.395216,
  // momentumX(10,42, 0-49)
    5.239619, 5.267014, 5.284798, 5.291317, 5.286037, 5.269451, 5.242799, 
    5.207787, 5.166325, 5.120343, 5.071693, 5.02209, 4.973096, 4.926105, 
    4.88232, 4.845045, 4.828703, 4.802299, 4.784326, 4.774885, 4.773208, 
    4.78215, 4.795608, 4.812541, 4.829976, 4.846041, 4.858818, 4.867209, 
    4.870528, 4.870278, 4.867199, 4.867313, 4.869003, 4.87472, 4.886584, 
    4.906005, 4.933528, 4.968866, 5.01106, 5.058681, 5.109999, 5.1631, 
    5.215928, 5.266298, 5.311891, 5.350265, 5.378949, 5.395628, 5.398466, 
    5.386536,
  // momentumX(10,43, 0-49)
    5.225125, 5.256631, 5.280723, 5.295022, 5.298166, 5.289894, 5.270908, 
    5.242608, 5.206801, 5.165462, 5.120562, 5.073971, 5.027399, 4.982369, 
    4.940185, 4.903838, 4.885886, 4.85994, 4.841307, 4.830328, 4.826455, 
    4.832383, 4.842665, 4.856229, 4.869998, 4.882415, 4.891881, 4.897665, 
    4.899386, 4.899063, 4.897659, 4.900507, 4.90607, 4.916288, 4.932685, 
    4.956121, 4.986723, 5.023946, 5.066707, 5.113532, 5.16267, 5.212178, 
    5.259955, 5.303786, 5.34137, 5.370416, 5.388793, 5.394788, 5.38742, 
    5.366787,
  // momentumX(10,44, 0-49)
    5.204635, 5.238729, 5.268057, 5.289697, 5.30149, 5.302343, 5.292276, 
    5.272214, 5.243718, 5.20869, 5.169145, 5.127045, 5.08421, 5.042264, 
    5.0026, 4.967926, 4.949046, 4.92391, 4.904885, 4.892501, 4.88643, 
    4.88929, 4.896282, 4.906398, 4.916552, 4.925547, 4.932125, 4.93589, 
    4.936687, 4.936886, 4.937493, 4.94312, 4.952159, 4.966044, 4.985777, 
    5.011779, 5.043863, 5.081303, 5.122929, 5.167236, 5.212452, 5.256604, 
    5.297564, 5.333117, 5.361072, 5.379413, 5.386541, 5.381553, 5.364513, 
    5.336632,
  // momentumX(10,45, 0-49)
    5.179212, 5.214012, 5.246877, 5.274645, 5.294554, 5.304733, 5.304421, 
    5.293918, 5.274354, 5.247395, 5.214958, 5.179004, 5.14139, 5.103791, 
    5.067675, 5.035524, 5.016601, 4.992625, 4.973468, 4.959824, 4.951601, 
    4.951439, 4.955157, 4.961893, 4.9686, 4.974474, 4.978585, 4.980832, 
    4.981196, 4.982283, 4.985005, 4.993274, 5.005284, 5.021986, 5.043922, 
    5.071142, 5.103206, 5.139245, 5.178025, 5.218019, 5.257449, 5.294353, 
    5.326642, 5.352213, 5.369123, 5.375821, 5.371424, 5.355994, 5.330694, 
    5.29772,
  // momentumX(10,46, 0-49)
    5.15041, 5.183906, 5.218145, 5.250115, 5.276795, 5.295731, 5.305416, 
    5.305406, 5.296213, 5.27905, 5.255547, 5.227502, 5.196701, 5.164815, 
    5.133346, 5.104626, 5.08668, 5.064239, 5.04522, 5.03049, 5.020214, 
    5.017181, 5.017759, 5.021304, 5.024827, 5.027922, 5.029962, 5.031085, 
    5.031336, 5.033477, 5.038228, 5.048871, 5.063292, 5.081979, 5.10506, 
    5.132253, 5.162891, 5.19597, 5.230196, 5.264036, 5.295753, 5.323472, 
    5.345274, 5.359347, 5.364205, 5.358969, 5.343636, 5.319263, 5.287948, 
    5.25254,
  // momentumX(10,47, 0-49)
    5.119985, 5.150326, 5.183611, 5.217366, 5.248749, 5.275069, 5.294239, 
    5.305062, 5.307268, 5.30139, 5.288529, 5.270121, 5.247734, 5.222944, 
    5.197252, 5.1729, 5.157071, 5.136595, 5.11804, 5.102479, 5.090351, 
    5.084734, 5.082446, 5.08311, 5.083791, 5.084471, 5.08479, 5.085076, 
    5.085362, 5.088531, 5.095047, 5.107666, 5.123862, 5.143695, 5.166904, 
    5.192897, 5.220782, 5.249414, 5.27744, 5.303342, 5.32549, 5.342224, 
    5.351979, 5.353467, 5.345912, 5.329299, 5.304561, 5.273603, 5.239101, 
    5.204047,
  // momentumX(10,48, 0-49)
    5.089595, 5.115337, 5.145545, 5.178566, 5.212147, 5.243782, 5.271115, 
    5.29231, 5.306252, 5.312603, 5.311698, 5.304386, 5.291848, 5.275453, 
    5.25664, 5.23762, 5.225192, 5.207209, 5.189566, 5.173572, 5.159956, 
    5.152224, 5.147508, 5.145734, 5.143994, 5.142636, 5.141529, 5.141139, 
    5.141435, 5.145405, 5.153227, 5.167259, 5.184483, 5.204558, 5.226863, 
    5.250508, 5.274375, 5.297177, 5.317502, 5.333895, 5.344922, 5.349295, 
    5.346019, 5.33458, 5.315123, 5.288604, 5.256801, 5.222151, 5.187412, 
    5.155191,
  // momentumX(10,49, 0-49)
    5.053679, 5.072524, 5.096591, 5.125384, 5.157755, 5.191944, 5.225796, 
    5.257071, 5.283777, 5.304451, 5.318295, 5.325191, 5.325613, 5.320494, 
    5.311103, 5.300251, 5.299141, 5.285053, 5.268355, 5.251288, 5.235315, 
    5.227765, 5.223431, 5.222784, 5.22031, 5.217353, 5.213843, 5.210539, 
    5.206765, 5.208167, 5.214479, 5.229855, 5.247833, 5.267559, 5.287977, 
    5.307836, 5.32576, 5.340317, 5.350102, 5.353841, 5.350516, 5.339516, 
    5.320797, 5.295008, 5.263525, 5.228363, 5.191968, 5.156848, 5.125219, 
    5.098701,
  // momentumX(11,0, 0-49)
    5.173462, 5.206308, 5.240257, 5.272574, 5.300474, 5.321579, 5.334246, 
    5.337715, 5.33208, 5.318138, 5.297173, 5.270765, 5.240604, 5.208375, 
    5.175654, 5.144077, 5.116427, 5.090436, 5.068562, 5.051296, 5.038685, 
    5.030923, 5.027062, 5.026567, 5.028524, 5.032345, 5.037494, 5.043713, 
    5.050945, 5.059712, 5.070448, 5.084126, 5.100892, 5.121141, 5.144976, 
    5.172139, 5.202004, 5.233603, 5.265666, 5.296687, 5.325003, 5.348888, 
    5.366683, 5.376942, 5.378628, 5.371307, 5.355311, 5.331816, 5.302765, 
    5.270608,
  // momentumX(11,1, 0-49)
    5.194742, 5.228152, 5.26071, 5.289646, 5.312393, 5.32699, 5.332311, 
    5.328114, 5.314935, 5.29389, 5.266475, 5.234376, 5.199319, 5.162972, 
    5.126867, 5.092795, 5.064954, 5.037652, 5.015035, 4.997619, 4.985379, 
    4.97889, 4.976613, 4.977965, 4.981647, 4.987005, 4.993341, 5.000309, 
    5.007703, 5.0163, 5.026547, 5.039942, 5.056371, 5.076459, 5.100532, 
    5.128533, 5.160006, 5.194112, 5.229676, 5.265248, 5.299183, 5.329723, 
    5.355093, 5.373639, 5.383974, 5.385177, 5.376961, 5.359829, 5.335091, 
    5.304753,
  // momentumX(11,2, 0-49)
    5.215133, 5.247335, 5.276393, 5.299809, 5.315543, 5.322279, 5.319528, 
    5.307566, 5.287278, 5.259983, 5.227242, 5.190721, 5.152076, 5.112883, 
    5.074576, 5.039062, 5.011899, 4.983998, 4.961249, 4.944171, 4.93268, 
    4.927715, 4.927212, 4.93057, 4.936181, 4.943317, 4.951117, 4.959096, 
    4.966879, 4.975387, 4.985026, 4.997762, 5.013227, 5.032263, 5.055445, 
    5.082962, 5.114574, 5.149624, 5.187086, 5.225627, 5.263697, 5.299596, 
    5.33156, 5.357855, 5.376884, 5.387331, 5.388323, 5.37959, 5.3616, 5.335593,
  // momentumX(11,3, 0-49)
    5.23278, 5.262092, 5.285949, 5.302372, 5.310034, 5.308362, 5.297498, 
    5.278173, 5.251532, 5.218977, 5.182038, 5.142278, 5.101216, 5.060287, 
    5.020789, 4.984736, 4.959036, 4.931108, 4.908727, 4.892389, 4.881948, 
    4.878703, 4.880101, 4.885571, 4.893275, 4.902404, 4.911927, 4.921201, 
    4.929637, 4.9382, 4.947193, 4.959, 4.972971, 4.990158, 5.011407, 
    5.037199, 5.067567, 5.102092, 5.139944, 5.17996, 5.220726, 5.260663, 
    5.298082, 5.331253, 5.358465, 5.378115, 5.388823, 5.389595, 5.380008, 
    5.360395,
  // momentumX(11,4, 0-49)
    5.246124, 5.271151, 5.28868, 5.297393, 5.296728, 5.286824, 5.26838, 
    5.242476, 5.21042, 5.173625, 5.133534, 5.091561, 5.049062, 5.007304, 
    4.967432, 4.931567, 4.908005, 4.880484, 4.858866, 4.843581, 4.83441, 
    4.833011, 4.836378, 4.843999, 4.853899, 4.86519, 4.876671, 4.887522, 
    4.896918, 4.905757, 4.914163, 4.924904, 4.936983, 4.951648, 4.970031, 
    4.992957, 5.020799, 5.053441, 5.090303, 5.130426, 5.172563, 5.215267, 
    5.256948, 5.295912, 5.330392, 5.358579, 5.378705, 5.389174, 5.388783, 
    5.376987,
  // momentumX(11,5, 0-49)
    5.254175, 5.273928, 5.284616, 5.285609, 5.277045, 5.259663, 5.234583, 
    5.203132, 5.1667, 5.126667, 5.08436, 5.041042, 4.997897, 4.956021, 
    4.916396, 4.881262, 4.860361, 4.83355, 4.812981, 4.798963, 4.791189, 
    4.79168, 4.796989, 4.80671, 4.818825, 4.832373, 4.846004, 4.858711, 
    4.86942, 4.878846, 4.88686, 4.896566, 4.906542, 4.918179, 4.932914, 
    4.951959, 4.976102, 5.005606, 5.040208, 5.079185, 5.121468, 5.165733, 
    5.210474, 5.254028, 5.294588, 5.330204, 5.358836, 5.378459, 5.387281, 
    5.384035,
  // momentumX(11,6, 0-49)
    5.256631, 5.270588, 5.274484, 5.268309, 5.25277, 5.229043, 5.198534, 
    5.162709, 5.122982, 5.080671, 5.036992, 4.993062, 4.949906, 4.90846, 
    4.869534, 4.835497, 4.817565, 4.791654, 4.772311, 4.759662, 4.753291, 
    4.755591, 4.762683, 4.77432, 4.788547, 4.804348, 4.820257, 4.835084, 
    4.847507, 4.857955, 4.865939, 4.874877, 4.882786, 4.891138, 4.901649, 
    4.915957, 4.935346, 4.960551, 4.991693, 5.028335, 5.069591, 5.114242, 
    5.160832, 5.2077, 5.252995, 5.294673, 5.33052, 5.358258, 5.375719, 
    5.381134,
  // momentumX(11,7, 0-49)
    5.253899, 5.261981, 5.259573, 5.247164, 5.225865, 5.197128, 5.162515, 
    5.123538, 5.081592, 5.037923, 4.993641, 4.949739, 4.907105, 4.866518, 
    4.828615, 4.795863, 4.780922, 4.756021, 4.737971, 4.726662, 4.721548, 
    4.72541, 4.733949, 4.747142, 4.763211, 4.781125, 4.799346, 4.816528, 
    4.831117, 4.843144, 4.851673, 4.860385, 4.866592, 4.871735, 4.877743, 
    4.88669, 4.900416, 4.920234, 4.94675, 4.979874, 5.018923, 5.062773, 
    5.109976, 5.158839, 5.207454, 5.253706, 5.295303, 5.329849, 5.355006, 
    5.36871,
  // momentumX(11,8, 0-49)
    5.246972, 5.249469, 5.241543, 5.224041, 5.198316, 5.165953, 5.128552, 
    5.087615, 5.044479, 5.000314, 4.956141, 4.912849, 4.871207, 4.831842, 
    4.795206, 4.763745, 4.751428, 4.727627, 4.710842, 4.700696, 4.696517, 
    4.701485, 4.710924, 4.725105, 4.742551, 4.762268, 4.782706, 4.802408, 
    4.81963, 4.83391, 4.843769, 4.853097, 4.858361, 4.860801, 4.86244, 
    4.865728, 4.873104, 4.886553, 4.907292, 4.935679, 4.971288, 5.01309, 
    5.059626, 5.109141, 5.159651, 5.208991, 5.254846, 5.29482, 5.326542, 
    5.347835,
  // momentumX(11,9, 0-49)
    5.237248, 5.234728, 5.222235, 5.200835, 5.17199, 5.1373, 5.09833, 
    5.056515, 5.013119, 4.96924, 4.925823, 4.883679, 4.843467, 4.805668, 
    4.770514, 4.740153, 4.729591, 4.707032, 4.691422, 4.682123, 4.678374, 
    4.683771, 4.693341, 4.707723, 4.725875, 4.746894, 4.769297, 4.791569, 
    4.811847, 4.829095, 4.841227, 4.852277, 4.857747, 4.858494, 4.856425, 
    4.854231, 4.854913, 4.861206, 4.875076, 4.897473, 4.92833, 4.966763, 
    5.011302, 5.060114, 5.111127, 5.162135, 5.210836, 5.254894, 5.292007, 
    5.319999,
  // momentumX(11,10, 0-49)
    5.226325, 5.219534, 5.203464, 5.179299, 5.148501, 5.112608, 5.073096, 
    5.031306, 4.988426, 4.94549, 4.903389, 4.862872, 4.824508, 4.788627, 
    4.755206, 4.725522, 4.715262, 4.694233, 4.679683, 4.670805, 4.666822, 
    4.671776, 4.680524, 4.694141, 4.712152, 4.733792, 4.757727, 4.782455, 
    4.806074, 4.826941, 4.84233, 4.856339, 4.863483, 4.86403, 4.859515, 
    4.852623, 4.846785, 4.845483, 4.851567, 4.866756, 4.891508, 4.925184, 
    4.966353, 5.013109, 5.063296, 5.114656, 5.164914, 5.211822, 5.253187, 
    5.286903,
  // momentumX(11,11, 0-49)
    5.215777, 5.205538, 5.186835, 5.160881, 5.129076, 5.092853, 5.05357, 
    5.01247, 4.970669, 4.929159, 4.888799, 4.850304, 4.814176, 4.780593, 
    4.749253, 4.719546, 4.70758, 4.688578, 4.67502, 4.666077, 4.661113, 
    4.664628, 4.671499, 4.683293, 4.700191, 4.72163, 4.746493, 4.773363, 
    4.800385, 4.825321, 4.844834, 4.86298, 4.873383, 4.875564, 4.870417, 
    4.860304, 4.848796, 4.840018, 4.837758, 4.844696, 4.862033, 4.889554, 
    4.925972, 4.969349, 5.01745, 5.067966, 5.118637, 5.167293, 5.211854, 
    5.250307,
  // momentumX(11,12, 0-49)
    5.206971, 5.194101, 5.173579, 5.146593, 5.114454, 5.078471, 5.039887, 
    4.99986, 4.959449, 4.919629, 4.88126, 4.845059, 4.811492, 4.78062, 
    4.751868, 4.72114, 4.705098, 4.688858, 4.676319, 4.666856, 4.660173, 
    4.661228, 4.665177, 4.674097, 4.688881, 4.709216, 4.734272, 4.762765, 
    4.792983, 4.822137, 4.846368, 4.869545, 4.884646, 4.890373, 4.886761, 
    4.875495, 4.859918, 4.844513, 4.833935, 4.83196, 4.84078, 4.860842, 
    4.891177, 4.929914, 4.974764, 5.023362, 5.073436, 5.12287, 5.169671, 
    5.211904,
  // momentumX(11,13, 0-49)
    5.200899, 5.186135, 5.164429, 5.136922, 5.104827, 5.069341, 5.031617, 
    4.992749, 4.953773, 4.915673, 4.879345, 4.845548, 4.814764, 4.787011, 
    4.761545, 4.728561, 4.7061, 4.693552, 4.682205, 4.671872, 4.662838, 
    4.660499, 4.66059, 4.665687, 4.677411, 4.695735, 4.72017, 4.749611, 
    4.782543, 4.815727, 4.844905, 4.873561, 4.8944, 4.905334, 4.90543, 
    4.895422, 4.878002, 4.857599, 4.839486, 4.828537, 4.828136, 4.839681, 
    4.862757, 4.895705, 4.936254, 4.981984, 5.030586, 5.079952, 5.128131, 
    5.173246,
  // momentumX(11,14, 0-49)
    5.198095, 5.182048, 5.159592, 5.13182, 5.099866, 5.064854, 5.027873, 
    4.989992, 4.952253, 4.915678, 4.881233, 4.849756, 4.82182, 4.797526, 
    4.776157, 4.739671, 4.70902, 4.701211, 4.69137, 4.679989, 4.668147, 
    4.661624, 4.657088, 4.65757, 4.665394, 4.680862, 4.703853, 4.733477, 
    4.768441, 4.805169, 4.839162, 4.873245, 4.9003, 4.917571, 4.923186, 
    4.916782, 4.900061, 4.876922, 4.852844, 4.83361, 4.823883, 4.826264, 
    4.841175, 4.867381, 4.902731, 4.944778, 4.991159, 5.039723, 5.088521, 
    5.135692,
  // momentumX(11,15, 0-49)
    5.198611, 5.181742, 5.158781, 5.130789, 5.098861, 5.064082, 5.027527, 
    4.990268, 4.953382, 4.917949, 4.885024, 4.855564, 4.83031, 4.809587, 
    4.793001, 4.752295, 4.712822, 4.710817, 4.702914, 4.690477, 4.67556, 
    4.664219, 4.654443, 4.649671, 4.652883, 4.664748, 4.685534, 4.714571, 
    4.750784, 4.790377, 4.82878, 4.867803, 4.900972, 4.92504, 4.93734, 
    4.936428, 4.922827, 4.899501, 4.871641, 4.845568, 4.827119, 4.820251, 
    4.826494, 4.845283, 4.874737, 4.912448, 4.955987, 5.003134, 5.051886, 
    5.100367,
  // momentumX(11,16, 0-49)
    5.202085, 5.184723, 5.161361, 5.133057, 5.10091, 5.066013, 5.029459, 
    4.99235, 4.955808, 4.920977, 4.889006, 4.860992, 4.837896, 4.820388, 
    4.808672, 4.76449, 4.717262, 4.722044, 4.716553, 4.703173, 4.685042, 
    4.668344, 4.652804, 4.642239, 4.640246, 4.647893, 4.665833, 4.693597, 
    4.730288, 4.771996, 4.814262, 4.857442, 4.896148, 4.926826, 4.946223, 
    4.951967, 4.943392, 4.922285, 4.893093, 4.862197, 4.836313, 4.820743, 
    4.818316, 4.829373, 4.852494, 4.885402, 4.925627, 4.970856, 5.019004, 
    5.068143,
  // momentumX(11,17, 0-49)
    5.207882, 5.190274, 5.166554, 5.137811, 5.105181, 5.069798, 5.032796, 
    4.995312, 4.95851, 4.923584, 4.891758, 4.864257, 4.842258, 4.826826, 
    4.818871, 4.77463, 4.723094, 4.735348, 4.732672, 4.718445, 4.696949, 
    4.674356, 4.652512, 4.635655, 4.627968, 4.630945, 4.645575, 4.671546, 
    4.708066, 4.751193, 4.796754, 4.843171, 4.886521, 4.923114, 4.949328, 
    4.962093, 4.959697, 4.942693, 4.914481, 4.881027, 4.849508, 4.826371, 
    4.815795, 4.819218, 4.835872, 4.863728, 4.900331, 4.943276, 4.990375, 
    5.039623,
  // momentumX(11,18, 0-49)
    5.215275, 5.197681, 5.173691, 5.144443, 5.111129, 5.074939, 5.037043, 
    4.998607, 4.960812, 4.924872, 4.892043, 4.863613, 4.840909, 4.825321, 
    4.818491, 4.781203, 4.73237, 4.751977, 4.752251, 4.737044, 4.711777, 
    4.682581, 4.653769, 4.630121, 4.616386, 4.614459, 4.625572, 4.649482, 
    4.685395, 4.729392, 4.777759, 4.826488, 4.873441, 4.914927, 4.947153, 
    4.966595, 4.970727, 4.958978, 4.933579, 4.899727, 4.8646, 4.835458, 
    4.817726, 4.814026, 4.824396, 4.847192, 4.880045, 4.920485, 4.966215, 
    5.015142,
  // momentumX(11,19, 0-49)
    5.223647, 5.206471, 5.182448, 5.152765, 5.118663, 5.081373, 5.042089, 
    5.001988, 4.962242, 4.924037, 4.888577, 4.857102, 4.830956, 4.811839, 
    4.802468, 4.782428, 4.748799, 4.774101, 4.776849, 4.759989, 4.72988, 
    4.692934, 4.656215, 4.62528, 4.605374, 4.598666, 4.606437, 4.628368, 
    4.663541, 4.708077, 4.758886, 4.809097, 4.858589, 4.903782, 4.940869, 
    4.966106, 4.976411, 4.9703, 4.948884, 4.916395, 4.87963, 4.846251, 
    4.822695, 4.812732, 4.817303, 4.835267, 4.864427, 4.902291, 4.94647, 
    4.994776,
  // momentumX(11,20, 0-49)
    5.228605, 5.209377, 5.183713, 5.153066, 5.118945, 5.08285, 5.046243, 
    5.010551, 4.977164, 4.947405, 4.922451, 4.903156, 4.889757, 4.881487, 
    4.876232, 0, 4.74619, 4.746288, 4.737542, 4.720608, 4.697607, 4.668127, 
    4.638677, 4.612827, 4.595506, 4.58938, 4.596458, 4.617135, 4.651025, 
    4.694868, 4.746641, 4.79661, 4.846766, 4.893705, 4.933717, 4.963015, 
    4.978206, 4.977147, 4.959987, 4.929938, 4.893122, 4.857208, 4.829299, 
    4.814166, 4.813659, 4.827224, 4.852918, 4.888282, 4.930861, 4.978384,
  // momentumX(11,21, 0-49)
    5.2353, 5.216488, 5.190962, 5.160259, 5.125952, 5.089577, 5.052596, 
    5.016393, 4.982272, 4.951435, 4.92492, 4.903454, 4.887238, 4.875626, 
    4.866798, 0, 4.797721, 4.792305, 4.77688, 4.75208, 4.720561, 4.678942, 
    4.639472, 4.605354, 4.581752, 4.571404, 4.576097, 4.595869, 4.629888, 
    4.674782, 4.72919, 4.780305, 4.832267, 4.881819, 4.925358, 4.959108, 
    4.979494, 4.983882, 4.97161, 4.944922, 4.909168, 4.871809, 4.840419, 
    4.820678, 4.815356, 4.824558, 4.846657, 4.879263, 4.919861, 4.966089,
  // momentumX(11,22, 0-49)
    5.239971, 5.221348, 5.19583, 5.165015, 5.130526, 5.093925, 5.056665, 
    5.020096, 4.985459, 4.95387, 4.926275, 4.903344, 4.885296, 4.871654, 
    4.860947, 0, 4.835303, 4.825794, 4.806291, 4.777096, 4.740961, 4.690882, 
    4.644479, 4.604306, 4.575753, 4.561767, 4.564087, 4.582548, 4.615982, 
    4.660958, 4.716836, 4.767711, 4.819979, 4.870557, 4.915993, 4.952604, 
    4.976768, 4.985557, 4.977713, 4.954643, 4.920895, 4.883494, 4.850173, 
    4.82724, 4.818252, 4.823944, 4.84304, 4.873272, 4.912107, 4.957114,
  // momentumX(11,23, 0-49)
    5.242476, 5.223934, 5.198411, 5.167542, 5.132972, 5.096276, 5.058898, 
    5.022161, 4.987256, 4.95525, 4.927035, 4.903254, 4.884159, 4.869406, 
    4.857812, 0, 4.860757, 4.848539, 4.826694, 4.795172, 4.756673, 4.700799, 
    4.649669, 4.605175, 4.572934, 4.556139, 4.556563, 4.573909, 4.606749, 
    4.651597, 4.708432, 4.75862, 4.810601, 4.861441, 4.90783, 4.9462, 
    4.97295, 4.984998, 4.980686, 4.960799, 4.929197, 4.892447, 4.858245, 
    4.833289, 4.82172, 4.824795, 4.841565, 4.869889, 4.907241, 4.951149,
  // momentumX(11,24, 0-49)
    5.242755, 5.224256, 5.198783, 5.167976, 5.133484, 5.096869, 5.059566, 
    5.022881, 4.987978, 4.955898, 4.927505, 4.903431, 4.883943, 4.868771, 
    4.856884, 0, 4.873823, 4.860311, 4.837456, 4.80504, 4.765738, 4.706779, 
    4.653216, 4.606438, 4.572193, 4.55386, 4.553253, 4.570012, 4.602548, 
    4.647337, 4.704798, 4.75439, 4.805976, 4.856723, 4.903411, 4.942552, 
    4.970578, 4.984347, 4.981996, 4.963964, 4.933707, 4.897477, 4.862895, 
    4.836847, 4.823806, 4.825346, 4.840734, 4.867923, 4.904401, 4.947665,
  // momentumX(11,25, 0-49)
    5.240794, 5.22232, 5.196975, 5.166369, 5.132127, 5.095788, 5.058773, 
    5.022375, 4.987755, 4.955944, 4.927806, 4.903964, 4.884675, 4.869664, 
    4.8579, 0, 4.873703, 4.860322, 4.837665, 4.805562, 4.766716, 4.707583, 
    4.654046, 4.607269, 4.572984, 4.554605, 4.553962, 4.570693, 4.603181, 
    4.647916, 4.705504, 4.754699, 4.80592, 4.856369, 4.902862, 4.941946, 
    4.970081, 4.984127, 4.982181, 4.964595, 4.934705, 4.898656, 4.864019, 
    4.837709, 4.824278, 4.825392, 4.84038, 4.86723, 4.903439, 4.946502,
  // momentumX(11,26, 0-49)
    5.236609, 5.218122, 5.192966, 5.162689, 5.128861, 5.092988, 5.056469, 
    5.020595, 4.98654, 4.955349, 4.927902, 4.904818, 4.886321, 4.872047, 
    4.860817, 0, 4.860604, 4.848742, 4.827468, 4.796851, 4.759639, 4.703284, 
    4.652233, 4.607754, 4.575406, 4.558476, 4.558778, 4.576014, 4.608685, 
    4.653347, 4.710508, 4.75958, 4.810529, 4.860532, 4.90638, 4.944607, 
    4.971689, 4.984544, 4.981393, 4.962756, 4.932151, 4.895843, 4.8614, 
    4.835618, 4.82288, 4.824695, 4.8403, 4.867644, 4.904226, 4.947563,
  // momentumX(11,27, 0-49)
    5.230247, 5.211652, 5.186687, 5.156816, 5.12353, 5.088286, 5.052456, 
    5.017334, 4.984122, 4.953905, 4.927598, 4.90583, 4.888774, 4.875917, 
    4.8658, 0, 4.835612, 4.826562, 4.807929, 4.780112, 4.745865, 4.695104, 
    4.648843, 4.608716, 4.580005, 4.565769, 4.567803, 4.585944, 4.618935, 
    4.663445, 4.719617, 4.768734, 4.819421, 4.868762, 4.913473, 4.950031, 
    4.97492, 4.985185, 4.979329, 4.958301, 4.926076, 4.889226, 4.855335, 
    4.83092, 4.819949, 4.823555, 4.84074, 4.869361, 4.906916, 4.950954,
  // momentumX(11,28, 0-49)
    5.221816, 5.202913, 5.178044, 5.148566, 5.115879, 5.081367, 5.046379, 
    5.012208, 4.980105, 4.951216, 4.926524, 4.906692, 4.891847, 4.881296, 
    4.873246, 0, 4.800921, 4.795757, 4.781104, 4.757642, 4.728002, 4.685359, 
    4.64586, 4.611671, 4.58779, 4.577054, 4.5813, 4.600579, 4.633968, 
    4.678254, 4.733004, 4.782204, 4.832494, 4.880813, 4.923745, 4.957682, 
    4.979128, 4.985353, 4.975339, 4.950729, 4.91621, 4.878789, 4.846007, 
    4.823902, 4.815784, 4.822229, 4.841906, 4.872549, 4.91166, 4.956846,
  // momentumX(11,29, 0-49)
    5.211528, 5.191969, 5.166947, 5.13771, 5.105555, 5.071788, 5.037718, 
    5.004653, 4.97389, 4.946674, 4.924098, 4.906909, 4.895241, 4.888247, 
    4.883862, 0, 4.758096, 4.757624, 4.74851, 4.73148, 4.7087, 4.676564, 
    4.645609, 4.618504, 4.600053, 4.593021, 4.59944, 4.61967, 4.653188, 
    4.696864, 4.749561, 4.798358, 4.847646, 4.894192, 4.934445, 4.964732, 
    4.981649, 4.982831, 4.967932, 4.939481, 4.902971, 4.865784, 4.835213, 
    4.816581, 4.812366, 4.8225, 4.845302, 4.8784, 4.919327, 4.965767,
  // momentumX(11,30, 0-49)
    5.203184, 5.185256, 5.161644, 5.13331, 5.101258, 5.066503, 5.030076, 
    4.993026, 4.956442, 4.921446, 4.889181, 4.860801, 4.837526, 4.82086, 
    4.81322, 4.793564, 4.759291, 4.783369, 4.786592, 4.771524, 4.744068, 
    4.707412, 4.671654, 4.641252, 4.621176, 4.613644, 4.620066, 4.640306, 
    4.673593, 4.716428, 4.766704, 4.814546, 4.862028, 4.905797, 4.942236, 
    4.967708, 4.97907, 4.974526, 4.954614, 4.922864, 4.885518, 4.850087, 
    4.823308, 4.809544, 4.810329, 4.82495, 4.851427, 4.887334, 4.930273, 
    4.978027,
  // momentumX(11,31, 0-49)
    5.191897, 5.173043, 5.149139, 5.121112, 5.08991, 5.056485, 5.021814, 
    4.986914, 4.952852, 4.920757, 4.891789, 4.867128, 4.847923, 4.835331, 
    4.830701, 4.793941, 4.74672, 4.765321, 4.765812, 4.751783, 4.728415, 
    4.699248, 4.671027, 4.647578, 4.633379, 4.630328, 4.639804, 4.661777, 
    4.695667, 4.737928, 4.785717, 4.832349, 4.877781, 4.918511, 4.950845, 
    4.971227, 4.976875, 4.966708, 4.942261, 4.908067, 4.87096, 4.838338, 
    4.81617, 4.807773, 4.813767, 4.832868, 4.862859, 4.901292, 4.945847, 
    4.994394,
  // momentumX(11,32, 0-49)
    5.182117, 5.162619, 5.138494, 5.110645, 5.079966, 5.047355, 5.013735, 
    4.980078, 4.947419, 4.916849, 4.889486, 4.866421, 4.848642, 4.836962, 
    4.832007, 4.788759, 4.739945, 4.751895, 4.749567, 4.736239, 4.716129, 
    4.69341, 4.671788, 4.654728, 4.646223, 4.647764, 4.660519, 4.684406, 
    4.718903, 4.760376, 4.805366, 4.850052, 4.892422, 4.928905, 4.955868, 
    4.970041, 4.969263, 4.95342, 4.925176, 4.889977, 4.854934, 4.826926, 
    4.810857, 4.808888, 4.820767, 4.844739, 4.87844, 4.919459, 4.965571, 
    5.014742,
  // momentumX(11,33, 0-49)
    5.174572, 5.154589, 5.13018, 5.102248, 5.071674, 5.039321, 5.00607, 
    4.972849, 4.940649, 4.910503, 4.883449, 4.860447, 4.842265, 4.829318, 
    4.82152, 4.779136, 4.735283, 4.740807, 4.736142, 4.723701, 4.706699, 
    4.689884, 4.674292, 4.663169, 4.660039, 4.665985, 4.681876, 4.707491, 
    4.742249, 4.782453, 4.824167, 4.866026, 4.904251, 4.935326, 4.955851, 
    4.96308, 4.955732, 4.934846, 4.90422, 4.869962, 4.83904, 4.817427, 
    4.808751, 4.814018, 4.832221, 4.861261, 4.898711, 4.942233, 4.989711, 
    5.039204,
  // momentumX(11,34, 0-49)
    5.170084, 5.149796, 5.125022, 5.096713, 5.065773, 5.033074, 4.999493, 
    4.965929, 4.933328, 4.902668, 4.874899, 4.850855, 4.831088, 4.815667, 
    4.803902, 4.766072, 4.730641, 4.730635, 4.724333, 4.713195, 4.699438, 
    4.68818, 4.678235, 4.672667, 4.674529, 4.684519, 4.703167, 4.730061, 
    4.764484, 4.802741, 4.840598, 4.878656, 4.91169, 4.936383, 4.949773, 
    4.949892, 4.936552, 4.912015, 4.881037, 4.849986, 4.825233, 4.811538, 
    4.81119, 4.824152, 4.848831, 4.882911, 4.923972, 4.969772, 5.0183, 
    5.067683,
  // momentumX(11,35, 0-49)
    5.16936, 5.149054, 5.123928, 5.095007, 5.063273, 5.029659, 4.99507, 
    4.960418, 4.926631, 4.894642, 4.865333, 4.839435, 4.817364, 4.798974, 
    4.783234, 4.750862, 4.725138, 4.7207, 4.713482, 4.704073, 4.693744, 
    4.687737, 4.683125, 4.682759, 4.689171, 4.702719, 4.723572, 4.751113, 
    4.784435, 4.819942, 4.853301, 4.886603, 4.913572, 4.931258, 4.937376, 
    4.930943, 4.912982, 4.886868, 4.857957, 4.832395, 4.815557, 4.810833, 
    4.819266, 4.839981, 4.870982, 4.909855, 4.954227, 5.001952, 5.051094, 
    5.099827,
  // momentumX(11,36, 0-49)
    5.172808, 5.152929, 5.127627, 5.098027, 5.065219, 5.030244, 4.994094, 
    4.95773, 4.922098, 4.888113, 4.856624, 4.828312, 4.803537, 4.782102, 
    4.762949, 4.735329, 4.718907, 4.711125, 4.703607, 4.696209, 4.689353, 
    4.688214, 4.688584, 4.693012, 4.703455, 4.719961, 4.742342, 4.769779, 
    4.801148, 4.833087, 4.861357, 4.889116, 4.909484, 4.920085, 4.919499, 
    4.907862, 4.887349, 4.862151, 4.837749, 4.819602, 4.811847, 4.816537, 
    4.833683, 4.861814, 4.898704, 4.941922, 4.989157, 5.038332, 5.08755, 
    5.134997,
  // momentumX(11,37, 0-49)
    5.180398, 5.161556, 5.136457, 5.106329, 5.072402, 5.035862, 4.997823, 
    4.959341, 4.921418, 4.884993, 4.850913, 4.819863, 4.792229, 4.767898, 
    4.746009, 4.72179, 4.713002, 4.702868, 4.695462, 4.6901, 4.686528, 
    4.689706, 4.694558, 4.703251, 4.717091, 4.735848, 4.758998, 4.785535, 
    4.814129, 4.841794, 4.864573, 4.886342, 4.900098, 4.904203, 4.898227, 
    4.883398, 4.862806, 4.841026, 4.823173, 4.813704, 4.815465, 4.829372, 
    4.854675, 4.889541, 4.931647, 4.978592, 5.028115, 5.07816, 5.126826, 
    5.172269,
  // momentumX(11,38, 0-49)
    5.191592, 5.174534, 5.150224, 5.119972, 5.085162, 5.047144, 5.007191, 
    4.966487, 4.926123, 4.887098, 4.850299, 4.816452, 4.786022, 4.759057, 
    4.735008, 4.712789, 4.70924, 4.697576, 4.690451, 4.686867, 4.686113, 
    4.692836, 4.701461, 4.713706, 4.730173, 4.750387, 4.773516, 4.798402, 
    4.82355, 4.846487, 4.86371, 4.879532, 4.88728, 4.886151, 4.876693, 
    4.861042, 4.842818, 4.826513, 4.816519, 4.816159, 4.827136, 4.849496, 
    4.882006, 4.922656, 4.969118, 5.019029, 5.070147, 5.120387, 5.167787, 
    5.210437,
  // momentumX(11,39, 0-49)
    5.205347, 5.190912, 5.168145, 5.138416, 5.103247, 5.064161, 5.022605, 
    4.979915, 4.937297, 4.895839, 4.856494, 4.820059, 4.787104, 4.757856, 
    4.732081, 4.710703, 4.709868, 4.697269, 4.690359, 4.688056, 4.689408, 
    4.698699, 4.710176, 4.72507, 4.743271, 4.764093, 4.786444, 4.809061, 
    4.830353, 4.848471, 4.860497, 4.870972, 4.873897, 4.869296, 4.858545, 
    4.844366, 4.830497, 4.82097, 4.819266, 4.827655, 4.846931, 4.876558, 
    4.915043, 4.960332, 5.010135, 5.06212, 5.114024, 5.163682, 5.209023, 
    5.248034,
  // momentumX(11,40, 0-49)
    5.220186, 5.209238, 5.188896, 5.160541, 5.125803, 5.086365, 5.043848, 
    4.999744, 4.955394, 4.911988, 4.870568, 4.832009, 4.796983, 4.765884, 
    4.73874, 4.717393, 4.717087, 4.703911, 4.69698, 4.695314, 4.697904, 
    4.708665, 4.721914, 4.738419, 4.75739, 4.777978, 4.798889, 4.81882, 
    4.836173, 4.849782, 4.857394, 4.863602, 4.863284, 4.857172, 4.847208, 
    4.836345, 4.828079, 4.825771, 4.831997, 4.848148, 4.874382, 4.90982, 
    4.95287, 5.001508, 5.053501, 5.106535, 5.158285, 5.206468, 5.248866, 
    5.283354,
  // momentumX(11,41, 0-49)
    5.23431, 5.227661, 5.210699, 5.184736, 5.151451, 5.112651, 5.070111, 
    5.025473, 4.980214, 4.935633, 4.892861, 4.852852, 4.816367, 4.783926, 
    4.755749, 4.733974, 4.732622, 4.719017, 4.711739, 4.710033, 4.712957, 
    4.724083, 4.737983, 4.755019, 4.773808, 4.793388, 4.812348, 4.829412, 
    4.84305, 4.852812, 4.85709, 4.860407, 4.858553, 4.852761, 4.845245, 
    4.838876, 4.836684, 4.841298, 4.854504, 4.87704, 4.908657, 4.948308, 
    4.994401, 5.044983, 5.097881, 5.150779, 5.201279, 5.246957, 5.285442, 
    5.314502,
  // momentumX(11,42, 0-49)
    5.245757, 5.244094, 5.231469, 5.209024, 5.178406, 5.141475, 5.100114, 
    5.056091, 5.011003, 4.966255, 4.923054, 4.882427, 4.845201, 4.811985, 
    4.783129, 4.76075, 4.75743, 4.7434, 4.735441, 4.733069, 4.735492, 
    4.745985, 4.759491, 4.776057, 4.793811, 4.811748, 4.828418, 4.84264, 
    4.853035, 4.859815, 4.861965, 4.863824, 4.861996, 4.857988, 4.854019, 
    4.852657, 4.856369, 4.867102, 4.886012, 4.913383, 4.948726, 4.99094, 
    5.038484, 5.089493, 5.141856, 5.193256, 5.241224, 5.283213, 5.316723, 
    5.33947,
  // momentumX(11,43, 0-49)
    5.252583, 5.256382, 5.248981, 5.231237, 5.20464, 5.171007, 5.132254, 
    5.090226, 5.046606, 5.002879, 4.96032, 4.92001, 4.882821, 4.849424, 
    4.820261, 4.797302, 4.791629, 4.777101, 4.768164, 4.764614, 4.765842, 
    4.774894, 4.787142, 4.802403, 4.818435, 4.834261, 4.848473, 4.860041, 
    4.867776, 4.872492, 4.873652, 4.875337, 4.87478, 4.873552, 4.873688, 
    4.877326, 4.886364, 4.902164, 4.925396, 4.95604, 4.993475, 5.036603, 
    5.083958, 5.133768, 5.18399, 5.232327, 5.276277, 5.313229, 5.340635, 
    5.356261,
  // momentumX(11,44, 0-49)
    5.253074, 5.262515, 5.261069, 5.249179, 5.228035, 5.199276, 5.164745, 
    5.12628, 5.085594, 5.044218, 5.003467, 4.964456, 4.928098, 4.895112, 
    4.866016, 4.842618, 4.834599, 4.819472, 4.809327, 4.804217, 4.803734, 
    4.810767, 4.821117, 4.834463, 4.848287, 4.861711, 4.873432, 4.882618, 
    4.888287, 4.891765, 4.892875, 4.89539, 4.896967, 4.89908, 4.90345, 
    4.911751, 4.925344, 4.945101, 4.971322, 5.003768, 5.041742, 5.084168, 
    5.129661, 5.176544, 5.222858, 5.266371, 5.304625, 5.335056, 5.355216, 
    5.363077,
  // momentumX(11,45, 0-49)
    5.245976, 5.260865, 5.26584, 5.260825, 5.246549, 5.224311, 5.19573, 
    5.162527, 5.126361, 5.08875, 5.05102, 5.014307, 4.97956, 4.947553, 
    4.918889, 4.895254, 4.885153, 4.869344, 4.85784, 4.850928, 4.848397, 
    4.853063, 4.861111, 4.872155, 4.883486, 4.894375, 4.903677, 4.910774, 
    4.914892, 4.917789, 4.919525, 4.923557, 4.927764, 4.933413, 4.941857, 
    4.954303, 4.971632, 4.994293, 5.02229, 5.055206, 5.092278, 5.13245, 
    5.174401, 5.216556, 5.257073, 5.293852, 5.324604, 5.34698, 5.358833, 
    5.358551,
  // momentumX(11,46, 0-49)
    5.230698, 5.250425, 5.261923, 5.264531, 5.258378, 5.244246, 5.223355, 
    5.197155, 5.167138, 5.134735, 5.101245, 5.067813, 5.035434, 5.004955, 
    4.977088, 4.953472, 4.941727, 4.925207, 4.912287, 4.903466, 4.898721, 
    4.900876, 4.90643, 4.914997, 4.923724, 4.932077, 4.939089, 4.944373, 
    4.94734, 4.950113, 4.952881, 4.958815, 4.965834, 4.974938, 4.987098, 
    5.003079, 5.023328, 5.047932, 5.076622, 5.108816, 5.143669, 5.180115, 
    5.216885, 5.252507, 5.285301, 5.313405, 5.334856, 5.347742, 5.35046, 
    5.342037,
  // momentumX(11,47, 0-49)
    5.207477, 5.23103, 5.248695, 5.259253, 5.262141, 5.257459, 5.24584, 
    5.228285, 5.205985, 5.18019, 5.152124, 5.122934, 5.093671, 5.065282, 
    5.03861, 5.015327, 5.00253, 4.985361, 4.971079, 4.96038, 4.953408, 
    4.953086, 4.956131, 4.962209, 4.968366, 4.974279, 4.979176, 4.982888, 
    4.984988, 4.987902, 4.991867, 4.999817, 5.009564, 5.021826, 5.037194, 
    5.056029, 5.07839, 5.104032, 5.132427, 5.162814, 5.194239, 5.225595, 
    5.255641, 5.283024, 5.306286, 5.323929, 5.334507, 5.336784, 5.329955, 
    5.313877,
  // momentumX(11,48, 0-49)
    5.177426, 5.203481, 5.226476, 5.244749, 5.257052, 5.262691, 5.261548, 
    5.253999, 5.240782, 5.222868, 5.201346, 5.177341, 5.151967, 5.126286, 
    5.101289, 5.078762, 5.06565, 5.04801, 5.03255, 5.020142, 5.011084, 
    5.008462, 5.009127, 5.012832, 5.016562, 5.020209, 5.023188, 5.025537, 
    5.026949, 5.030105, 5.035226, 5.045074, 5.057245, 5.072175, 5.090107, 
    5.111032, 5.134658, 5.16043, 5.187572, 5.215123, 5.242, 5.267024, 
    5.288981, 5.30666, 5.318905, 5.324718, 5.323361, 5.314494, 5.298303, 
    5.275572,
  // momentumX(11,49, 0-49)
    5.130487, 5.157133, 5.184359, 5.21029, 5.233043, 5.250996, 5.26301, 
    5.268517, 5.267499, 5.260395, 5.247995, 5.231311, 5.211483, 5.189702, 
    5.167173, 5.146682, 5.140685, 5.122538, 5.104847, 5.089356, 5.0769, 
    5.074059, 5.074942, 5.079597, 5.082418, 5.084044, 5.083921, 5.082497, 
    5.079126, 5.079224, 5.082874, 5.095003, 5.110043, 5.128022, 5.148745, 
    5.171737, 5.196276, 5.221437, 5.24613, 5.269165, 5.289305, 5.305318, 
    5.316079, 5.32065, 5.318389, 5.309089, 5.293078, 5.271255, 5.245065, 
    5.216325,
  // momentumX(12,0, 0-49)
    5.283156, 5.303393, 5.315825, 5.319623, 5.31465, 5.301387, 5.280786, 
    5.254111, 5.222781, 5.188264, 5.151982, 5.115261, 5.079288, 5.045088, 
    5.013504, 4.985375, 4.962522, 4.942296, 4.926528, 4.915215, 4.908121, 
    4.905272, 4.90585, 4.909438, 4.915286, 4.922814, 4.93137, 4.940413, 
    4.949502, 4.958674, 4.967987, 4.978175, 4.989471, 5.002637, 5.018452, 
    5.037585, 5.060488, 5.087313, 5.117883, 5.15169, 5.18792, 5.225489, 
    5.263074, 5.299156, 5.332043, 5.359944, 5.381062, 5.393738, 5.396669, 
    5.389134,
  // momentumX(12,1, 0-49)
    5.289672, 5.306209, 5.313846, 5.31217, 5.301459, 5.28255, 5.256652, 
    5.225194, 5.189679, 5.15159, 5.112332, 5.073187, 5.035285, 4.999592, 
    4.966884, 4.938138, 4.916506, 4.896032, 4.880301, 4.86932, 4.862805, 
    4.861174, 4.863127, 4.868292, 4.875661, 4.884639, 4.894459, 4.904496, 
    4.91414, 4.923573, 4.932739, 4.942745, 4.953437, 4.965678, 4.980408, 
    4.998491, 5.020582, 5.047031, 5.077825, 5.112586, 5.150586, 5.19079, 
    5.231888, 5.272332, 5.310356, 5.344034, 5.371366, 5.390417, 5.399523, 
    5.397548,
  // momentumX(12,2, 0-49)
    5.289351, 5.301156, 5.303457, 5.296273, 5.280246, 5.256473, 5.226311, 
    5.191248, 5.152781, 5.112347, 5.071281, 5.030792, 4.991937, 4.955608, 
    4.922512, 4.893762, 4.873818, 4.853418, 4.837952, 4.827422, 4.821506, 
    4.821013, 4.824201, 4.830774, 4.839534, 4.849892, 4.860994, 4.872135, 
    4.882534, 4.892459, 4.901697, 4.911676, 4.921791, 4.932947, 4.946202, 
    4.962606, 4.983036, 5.008065, 5.037891, 5.072294, 5.110664, 5.152039, 
    5.195147, 5.238437, 5.280128, 5.318251, 5.350725, 5.375486, 5.390674, 
    5.394858,
  // momentumX(12,3, 0-49)
    5.282612, 5.289087, 5.285932, 5.273549, 5.252862, 5.225129, 5.191766, 
    5.154241, 5.113979, 5.072326, 5.030522, 4.989674, 4.950751, 4.914566, 
    4.881744, 4.85353, 4.835714, 4.815639, 4.800602, 4.790585, 4.785224, 
    4.785729, 4.789946, 4.797691, 4.807655, 4.819279, 4.831649, 4.843991, 
    4.855368, 4.866057, 4.875648, 4.885847, 4.895519, 4.905539, 4.917031, 
    4.931207, 4.949178, 4.971781, 4.999463, 5.032219, 5.069589, 5.110712, 
    5.154368, 5.199042, 5.24297, 5.2842, 5.320669, 5.350304, 5.37118, 5.381702,
  // momentumX(12,4, 0-49)
    5.270433, 5.271401, 5.263016, 5.245987, 5.221428, 5.190666, 5.15511, 
    5.116154, 5.07512, 5.033241, 4.991632, 4.951296, 4.9131, 4.877757, 
    4.845793, 4.818586, 4.803279, 4.783717, 4.769216, 4.759707, 4.754789, 
    4.756079, 4.761035, 4.769634, 4.780541, 4.793252, 4.806829, 4.820447, 
    4.833023, 4.844786, 4.855074, 4.865842, 4.87534, 4.884321, 4.893908, 
    4.905432, 4.92024, 4.93947, 4.963875, 4.993721, 5.02876, 5.068261, 
    5.111091, 5.155785, 5.200624, 5.243716, 5.283067, 5.316677, 5.342657, 
    5.359342,
  // momentumX(12,5, 0-49)
    5.254186, 5.249829, 5.236703, 5.215734, 5.188132, 5.155237, 5.118395, 
    5.078903, 5.037965, 4.996687, 4.956069, 4.916993, 4.880211, 4.84632, 
    4.815726, 4.789899, 4.777379, 4.758461, 4.744543, 4.735467, 4.730793, 
    4.732566, 4.737878, 4.74691, 4.758401, 4.771935, 4.786589, 4.801508, 
    4.815494, 4.828657, 4.840042, 4.851838, 4.861586, 4.869823, 4.877574, 
    4.886226, 4.897335, 4.912361, 4.932431, 4.958163, 4.989584, 5.026161, 
    5.066878, 5.110339, 5.154894, 5.19872, 5.239929, 5.276628, 5.30701, 
    5.329417,
  // momentumX(12,6, 0-49)
    5.235466, 5.226234, 5.209022, 5.184886, 5.155065, 5.120851, 5.083508, 
    5.044224, 5.004089, 4.964089, 4.925107, 4.88791, 4.853123, 4.821205, 
    4.792401, 4.768209, 4.758565, 4.740386, 4.727033, 4.718237, 4.713521, 
    4.715374, 4.720548, 4.729478, 4.741088, 4.755076, 4.770578, 4.786751, 
    4.802309, 4.817187, 4.830103, 4.84348, 4.854072, 4.862099, 4.868368, 
    4.874223, 4.881364, 4.891574, 4.906406, 4.926915, 4.953505, 4.985915, 
    5.023302, 5.064378, 5.107562, 5.151116, 5.193247, 5.232182, 5.266211, 
    5.293715,
  // momentumX(12,7, 0-49)
    5.215919, 5.202434, 5.181869, 5.155337, 5.124051, 5.089231, 5.052039, 
    5.013558, 4.974773, 4.936571, 4.899731, 4.864904, 4.832586, 4.803066, 
    4.776391, 4.753929, 4.746964, 4.729606, 4.716753, 4.708011, 4.702882, 
    4.704314, 4.708754, 4.716944, 4.728096, 4.742053, 4.758061, 4.775326, 
    4.792534, 4.809388, 4.824256, 4.839813, 4.851985, 4.860579, 4.86606, 
    4.869582, 4.872879, 4.878002, 4.88695, 4.901301, 4.921952, 4.949025, 
    4.981931, 5.019534, 5.060344, 5.102702, 5.144898, 5.185256, 5.222154, 
    5.254018,
  // momentumX(12,8, 0-49)
    5.197084, 5.180053, 5.15687, 5.128651, 5.096552, 5.0617, 5.02516, 
    4.987918, 4.950877, 4.914841, 4.880503, 4.848413, 4.818925, 4.792144, 
    4.76786, 4.747036, 4.742175, 4.725766, 4.713326, 4.70436, 4.698389, 
    4.698829, 4.701871, 4.708604, 4.71863, 4.731961, 4.748012, 4.766073, 
    4.784878, 4.803852, 4.82102, 4.839316, 4.853869, 4.863999, 4.869711, 
    4.871802, 4.871869, 4.872107, 4.874922, 4.882471, 4.896258, 4.916928, 
    4.944264, 4.977354, 5.014838, 5.055129, 5.096582, 5.137584, 5.17657, 
    5.212003,
  // momentumX(12,9, 0-49)
    5.180264, 5.160401, 5.13527, 5.105958, 5.07355, 5.03908, 5.003524, 
    4.967793, 4.932725, 4.899067, 4.86745, 4.838332, 4.811933, 4.788154, 
    4.766489, 4.747004, 4.743248, 4.728023, 4.715933, 4.706465, 4.699218, 
    4.698076, 4.699035, 4.70357, 4.711748, 4.723778, 4.739289, 4.757714, 
    4.777895, 4.798965, 4.818629, 4.840088, 4.857762, 4.870472, 4.877666, 
    4.879622, 4.877593, 4.873718, 4.870685, 4.871213, 4.877508, 4.890886, 
    4.911653, 4.939244, 4.972483, 5.00987, 5.049802, 5.090693, 5.131, 5.169196,
  // momentumX(12,10, 0-49)
    5.166411, 5.144372, 5.117849, 5.087887, 5.0555, 5.021643, 4.987225, 
    4.9531, 4.920068, 4.888845, 4.86002, 4.833982, 4.810833, 4.790262, 
    4.771456, 4.752806, 4.748785, 4.735146, 4.723433, 4.713244, 4.704352, 
    4.701074, 4.699321, 4.700947, 4.706553, 4.716559, 4.730864, 4.749084, 
    4.770245, 4.79319, 4.815342, 4.840149, 4.861498, 4.877731, 4.887707, 
    4.891069, 4.888515, 4.881875, 4.873897, 4.867746, 4.866354, 4.871841, 
    4.885215, 4.906405, 4.934523, 4.968196, 5.005853, 5.045899, 5.086775, 
    5.126939,
  // momentumX(12,11, 0-49)
    5.156057, 5.132392, 5.104886, 5.074547, 5.042329, 5.009131, 4.975822, 
    4.943227, 4.912133, 4.883249, 4.85715, 4.83418, 4.814344, 4.797164, 
    4.781535, 4.763055, 4.757185, 4.745727, 4.734569, 4.723561, 4.712773, 
    4.706907, 4.701915, 4.700012, 4.70236, 4.709619, 4.721997, 4.739341, 
    4.760933, 4.785336, 4.809756, 4.837816, 4.863089, 4.883525, 4.89742, 
    4.90373, 4.902445, 4.894832, 4.883407, 4.871558, 4.862848, 4.860272, 
    4.865705, 4.879758, 4.901966, 4.931159, 4.965813, 5.004309, 5.045033, 
    5.086396,
  // momentumX(12,12, 0-49)
    5.149285, 5.12441, 5.096178, 5.065566, 5.033495, 5.000843, 4.968459, 
    4.937173, 4.907782, 4.881011, 4.857444, 4.837414, 4.820879, 4.807252, 
    4.795251, 4.776213, 4.766981, 4.758471, 4.748212, 4.73646, 4.723689, 
    4.714914, 4.706287, 4.700346, 4.698822, 4.702633, 4.712355, 4.728104, 
    4.74946, 4.774756, 4.801041, 4.831972, 4.861088, 4.886032, 4.904624, 
    4.915174, 4.916892, 4.910286, 4.897347, 4.881368, 4.866335, 4.856068, 
    4.853416, 4.859857, 4.875521, 4.899554, 4.930533, 4.966812, 5.006703, 
    5.048541,
  // momentumX(12,13, 0-49)
    5.145769, 5.119963, 5.09112, 5.060205, 5.028135, 4.995795, 4.964047, 
    4.933748, 4.905724, 4.880737, 4.859405, 4.842088, 4.828754, 4.818828, 
    4.811018, 4.790828, 4.777141, 4.772433, 4.763588, 4.751352, 4.736684, 
    4.724803, 4.712266, 4.701881, 4.695943, 4.695662, 4.70202, 4.715442, 
    4.735847, 4.761384, 4.789021, 4.822229, 4.854795, 4.884152, 4.90777, 
    4.923401, 4.929517, 4.925776, 4.913407, 4.895278, 4.875484, 4.858485, 
    4.848105, 4.846823, 4.855548, 4.87389, 4.900612, 4.934071, 4.9725, 5.01414,
  // momentumX(12,14, 0-49)
    5.144871, 5.118295, 5.088853, 5.057521, 5.02524, 4.992924, 4.961475, 
    4.931789, 4.904742, 4.881144, 4.861664, 4.846729, 4.836396, 4.830227, 
    4.827164, 4.805708, 4.787249, 4.787188, 4.780379, 4.768078, 4.751752, 
    4.736667, 4.720029, 4.704872, 4.694035, 4.689069, 4.691406, 4.701812, 
    4.720558, 4.745669, 4.774117, 4.808887, 4.844282, 4.877623, 4.906136, 
    4.927167, 4.938556, 4.939137, 4.929252, 4.911079, 4.888462, 4.866208, 
    4.848984, 4.840306, 4.842016, 4.854346, 4.876366, 4.906497, 4.942909, 
    4.983748,
  // momentumX(12,15, 0-49)
    5.145796, 5.118527, 5.088447, 5.056561, 5.023852, 4.991281, 4.959796, 
    4.930346, 4.903856, 4.881192, 4.863095, 4.850088, 4.842387, 4.839818, 
    4.841783, 4.819959, 4.797536, 4.802824, 4.798692, 4.786848, 4.769209, 
    4.750873, 4.72998, 4.709755, 4.693579, 4.683396, 4.681126, 4.687901, 
    4.70434, 4.728413, 4.75718, 4.792764, 4.83025, 4.866904, 4.899821, 
    4.926082, 4.943048, 4.948842, 4.942933, 4.92663, 4.903234, 4.877543, 
    4.854808, 4.839509, 4.834488, 4.840753, 4.857808, 4.884229, 4.918171, 
    4.957691,
  // momentumX(12,16, 0-49)
    5.14775, 5.119838, 5.089086, 5.056542, 5.023234, 4.99017, 4.958349, 
    4.928762, 4.902383, 4.88013, 4.862822, 4.851107, 4.845402, 4.84588, 
    4.852536, 4.832886, 4.808788, 4.819836, 4.818934, 4.808081, 4.789505, 
    4.767872, 4.742556, 4.716972, 4.695046, 4.67918, 4.671813, 4.674458, 
    4.688052, 4.710579, 4.739286, 4.774993, 4.813807, 4.852983, 4.889573, 
    4.920512, 4.942851, 4.954165, 4.953143, 4.940207, 4.917892, 4.890668, 
    4.864047, 4.843275, 4.83217, 4.832603, 4.844646, 4.867138, 4.898277, 
    4.936063,
  // momentumX(12,17, 0-49)
    5.150093, 5.121617, 5.090219, 5.056981, 5.022968, 4.989228, 4.956792, 
    4.926682, 4.899899, 4.877413, 4.860113, 4.84878, 4.844049, 4.846456, 
    4.856596, 4.843801, 4.822259, 4.838977, 4.841652, 4.832212, 4.813004, 
    4.787975, 4.758004, 4.726743, 4.698685, 4.676764, 4.663949, 4.662121, 
    4.672501, 4.693131, 4.72155, 4.756793, 4.796225, 4.837117, 4.876529, 
    4.911358, 4.938486, 4.955118, 4.959318, 4.950685, 4.930918, 4.903908, 
    4.875101, 4.850234, 4.833983, 4.829096, 4.836311, 4.854834, 4.882985, 
    4.918743,
  // momentumX(12,18, 0-49)
    5.152446, 5.123583, 5.091654, 5.057766, 5.023003, 4.988423, 4.955067, 
    4.923962, 4.896122, 4.872548, 4.854192, 4.841951, 4.836679, 4.839291, 
    4.851016, 4.851833, 4.839601, 4.861182, 4.867465, 4.859635, 4.839867, 
    4.81117, 4.776155, 4.738822, 4.704293, 4.676091, 4.657684, 4.651282, 
    4.65831, 4.676892, 4.704975, 4.739322, 4.778765, 4.820615, 4.861983, 
    4.8998, 4.930897, 4.952261, 4.961515, 4.957573, 4.941316, 4.915917, 
    4.886491, 4.85898, 4.838706, 4.829237, 4.832021, 4.846715, 4.871841, 
    4.905409,
  // momentumX(12,19, 0-49)
    5.154763, 5.125841, 5.093623, 5.059199, 5.023643, 4.987998, 4.95329, 
    4.920535, 4.890742, 4.864912, 4.844035, 4.829114, 4.82127, 4.821993, 
    4.833523, 4.855882, 4.862566, 4.887558, 4.897141, 4.890828, 4.870145, 
    4.837114, 4.796288, 4.752288, 4.710979, 4.67649, 4.652683, 4.64197, 
    4.645842, 4.66249, 4.690382, 4.723572, 4.762553, 4.804698, 4.847201, 
    4.887078, 4.921197, 4.946469, 4.960234, 4.960886, 4.948586, 4.925761, 
    4.897009, 4.868209, 4.845094, 4.831927, 4.83085, 4.842024, 4.864239, 
    4.895589,
  // momentumX(12,20, 0-49)
    5.154693, 5.1242, 5.09093, 5.056166, 5.021146, 4.987069, 4.955105, 
    4.926386, 4.901967, 4.88274, 4.869288, 4.861674, 4.859224, 4.860402, 
    4.862944, 0, 4.887241, 4.889175, 4.884861, 4.87331, 4.854144, 4.824542, 
    4.78899, 4.749675, 4.711314, 4.677715, 4.653001, 4.640221, 4.641569, 
    4.655976, 4.682993, 4.71405, 4.751464, 4.792706, 4.835068, 4.875674, 
    4.911485, 4.939419, 4.956679, 4.961297, 4.952844, 4.933036, 4.905849, 
    4.876883, 4.852042, 4.836103, 4.831837, 4.839926, 4.859478, 4.888717,
  // momentumX(12,21, 0-49)
    5.155864, 5.125593, 5.092457, 5.057732, 5.02263, 4.988307, 4.955864, 
    4.926349, 4.90071, 4.879722, 4.863865, 4.853156, 4.846985, 4.843976, 
    4.841977, 0, 4.928431, 4.928067, 4.921334, 4.906662, 4.883474, 4.84574, 
    4.802858, 4.756638, 4.712227, 4.67375, 4.64543, 4.630235, 4.630127, 
    4.64397, 4.671875, 4.702372, 4.7396, 4.78107, 4.82414, 4.866025, 
    4.903787, 4.934397, 4.954999, 4.963388, 4.958678, 4.941965, 4.916625, 
    4.887901, 4.861739, 4.843331, 4.83602, 4.841007, 4.857741, 4.884601,
  // momentumX(12,22, 0-49)
    5.156168, 5.126009, 5.092949, 5.05825, 5.023098, 4.988604, 4.955816, 
    4.925714, 4.899168, 4.876884, 4.859283, 4.846379, 4.837635, 4.831826, 
    4.826962, 0, 4.95737, 4.955109, 4.947015, 4.931, 4.906226, 4.863213, 
    4.81588, 4.765259, 4.716686, 4.674536, 4.643195, 4.62569, 4.623909, 
    4.63674, 4.664946, 4.694184, 4.7305, 4.771442, 4.814431, 4.856776, 
    4.895633, 4.928053, 4.951179, 4.962662, 4.96128, 4.947614, 4.924472, 
    4.896675, 4.870069, 4.850082, 4.840516, 4.843034, 4.857418, 4.882221,
  // momentumX(12,23, 0-49)
    5.155862, 5.125789, 5.092804, 5.058161, 5.023019, 4.988459, 4.955489, 
    4.925042, 4.897942, 4.874845, 4.856148, 4.84187, 4.831531, 4.824033, 
    4.817537, 0, 4.976377, 4.972693, 4.963794, 4.947212, 4.921901, 4.875348, 
    4.825215, 4.771749, 4.720391, 4.675718, 4.642266, 4.623123, 4.620123, 
    4.632184, 4.660638, 4.688662, 4.724012, 4.764284, 4.806946, 4.849384, 
    4.888843, 4.92245, 4.947373, 4.961187, 4.962439, 4.951327, 4.930201, 
    4.903494, 4.876895, 4.855958, 4.8448, 4.845447, 4.857971, 4.881085,
  // momentumX(12,24, 0-49)
    5.155117, 5.125144, 5.092268, 5.057733, 5.022682, 4.988179, 4.955212, 
    4.924688, 4.897405, 4.873996, 4.85484, 4.839958, 4.828905, 4.820646, 
    4.81344, 0, 4.985891, 4.981441, 4.972165, 4.95543, 4.930089, 4.881607, 
    4.830071, 4.775189, 4.722447, 4.676545, 4.642097, 4.622215, 4.618693, 
    4.630451, 4.65923, 4.686486, 4.721179, 4.760937, 4.803261, 4.84558, 
    4.885197, 4.919293, 4.945075, 4.960088, 4.962771, 4.953119, 4.93321, 
    4.907235, 4.880754, 4.85936, 4.84734, 4.846935, 4.858387, 4.880515,
  // momentumX(12,25, 0-49)
    5.154003, 5.124162, 5.091442, 5.057076, 5.022206, 4.987893, 4.955125, 
    4.924804, 4.897723, 4.874507, 4.855525, 4.840787, 4.829843, 4.821658, 
    4.814504, 0, 4.985445, 4.981015, 4.971813, 4.955236, 4.930161, 4.881445, 
    4.829905, 4.775073, 4.722418, 4.676649, 4.642362, 4.622644, 4.61925, 
    4.63111, 4.66012, 4.687131, 4.721565, 4.761066, 4.803155, 4.84528, 
    4.884767, 4.918823, 4.94467, 4.959867, 4.962834, 4.953512, 4.933909, 
    4.908139, 4.88171, 4.860214, 4.847972, 4.847279, 4.858426, 4.880264,
  // momentumX(12,26, 0-49)
    5.152479, 5.122794, 5.090271, 5.056139, 5.021544, 4.98756, 4.955191, 
    4.925356, 4.898864, 4.876347, 4.858164, 4.84431, 4.834285, 4.826993, 
    4.820641, 0, 4.975043, 4.971416, 4.962752, 4.946657, 4.92212, 4.874942, 
    4.824836, 4.771557, 4.72049, 4.676219, 4.64323, 4.624537, 4.621883, 
    4.634203, 4.663285, 4.690606, 4.725205, 4.764738, 4.80672, 4.848597, 
    4.887678, 4.921165, 4.946287, 4.960632, 4.962692, 4.952519, 4.932245, 
    4.906088, 4.879598, 4.858325, 4.846496, 4.846295, 4.857932, 4.880213,
  // momentumX(12,27, 0-49)
    5.150397, 5.120863, 5.088561, 5.054716, 5.020484, 4.986965, 4.955193, 
    4.926123, 4.900596, 4.879271, 4.862515, 4.85029, 4.842027, 4.836516, 
    4.831839, 0, 4.955084, 4.952917, 4.945256, 4.930057, 4.906505, 4.862667, 
    4.815493, 4.76527, 4.717227, 4.67572, 4.645051, 4.628139, 4.626747, 
    4.639816, 4.668792, 4.696878, 4.731983, 4.77176, 4.813708, 4.855239, 
    4.893616, 4.925999, 4.949613, 4.96211, 4.962144, 4.950032, 4.928223, 
    4.901196, 4.874612, 4.853933, 4.843158, 4.844211, 4.857095, 4.880501,
  // momentumX(12,28, 0-49)
    5.147523, 5.118073, 5.085974, 5.052443, 5.018648, 4.985715, 4.954721, 
    4.926675, 4.902474, 4.882824, 4.868122, 4.858309, 4.85273, 4.850033, 
    4.848179, 0, 4.926608, 4.926298, 4.920071, 4.906347, 4.884541, 4.845834, 
    4.803155, 4.757463, 4.713751, 4.676086, 4.648576, 4.634062, 4.63437, 
    4.648452, 4.677229, 4.706404, 4.742229, 4.782332, 4.82418, 4.865112, 
    4.902321, 4.932904, 4.95409, 4.963649, 4.960521, 4.945456, 4.921401, 
    4.893226, 4.866715, 4.847156, 4.838172, 4.84128, 4.85618, 4.881395,
  // momentumX(12,29, 0-49)
    5.143562, 5.11403, 5.082041, 5.048799, 5.015478, 4.983227, 4.953168, 
    4.926374, 4.903827, 4.886317, 4.874309, 4.867758, 4.86593, 4.867328, 
    4.869853, 0, 4.889934, 4.891613, 4.88732, 4.875996, 4.857266, 4.825638, 
    4.789297, 4.749714, 4.711526, 4.678509, 4.654641, 4.642774, 4.644877, 
    4.659924, 4.688231, 4.718379, 4.754757, 4.794957, 4.836395, 4.876332, 
    4.911868, 4.940042, 4.958111, 4.964036, 4.957141, 4.938742, 4.912372, 
    4.883308, 4.857393, 4.839608, 4.833077, 4.838827, 4.856208, 4.883573,
  // momentumX(12,30, 0-49)
    5.140514, 5.112536, 5.081708, 5.049011, 5.015432, 4.981946, 4.949521, 
    4.919111, 4.891653, 4.868042, 4.849143, 4.835805, 4.82899, 4.830027, 
    4.841019, 4.861464, 4.864655, 4.888956, 4.899061, 4.894265, 4.875897, 
    4.843383, 4.804152, 4.761779, 4.721758, 4.68805, 4.664435, 4.653369, 
    4.656442, 4.672151, 4.699848, 4.730855, 4.767568, 4.807538, 4.848127, 
    4.886528, 4.91977, 4.944874, 4.959198, 4.960996, 4.950107, 4.928501, 
    4.900321, 4.871173, 4.846792, 4.831698, 4.828403, 4.837403, 4.857709, 
    4.887527,
  // momentumX(12,31, 0-49)
    5.134956, 5.106979, 5.076535, 5.044599, 5.012144, 4.980138, 4.949538, 
    4.921287, 4.896299, 4.875444, 4.859525, 4.84926, 4.845331, 4.848502, 
    4.859925, 4.859009, 4.845135, 4.865917, 4.872577, 4.866015, 4.848228, 
    4.820029, 4.786397, 4.750472, 4.717049, 4.68944, 4.671017, 4.664021, 
    4.67, 4.687367, 4.714871, 4.746837, 4.783939, 4.823677, 4.863338, 
    4.900009, 4.93064, 4.952261, 4.962398, 4.959703, 4.944641, 4.919906, 
    4.890231, 4.861438, 4.83902, 4.826921, 4.826994, 4.839206, 4.862264, 
    4.894248,
  // momentumX(12,32, 0-49)
    5.129212, 5.101433, 5.071481, 5.040294, 5.008811, 4.97796, 4.948673, 
    4.921868, 4.898431, 4.87919, 4.864866, 4.856045, 4.853179, 4.856658, 
    4.867016, 4.852871, 4.831022, 4.847097, 4.850173, 4.841893, 4.824452, 
    4.79999, 4.771226, 4.741108, 4.713883, 4.692271, 4.679163, 4.676469, 
    4.685562, 4.704714, 4.732142, 4.764843, 4.801892, 4.840762, 4.878683, 
    4.912685, 4.939712, 4.956912, 4.96214, 4.954616, 4.93555, 4.908378, 
    4.878297, 4.851113, 4.831837, 4.823677, 4.827783, 4.84363, 4.869668, 
    4.90391,
  // momentumX(12,33, 0-49)
    5.12343, 5.095872, 5.066374, 5.035829, 5.005118, 4.975122, 4.946723, 
    4.920801, 4.898202, 4.879708, 4.865957, 4.8574, 4.854257, 4.856545, 
    4.864198, 4.843874, 4.820434, 4.831309, 4.831038, 4.821383, 4.804472, 
    4.783561, 4.75934, 4.73466, 4.713286, 4.697415, 4.689446, 4.690929, 
    4.70299, 4.723768, 4.751048, 4.784074, 4.82048, 4.857722, 4.89301, 
    4.92337, 4.945841, 4.957834, 4.957703, 4.945395, 4.922944, 4.894461, 
    4.865391, 4.841245, 4.82632, 4.822978, 4.831672, 4.851446, 4.880571, 
    4.91704,
  // momentumX(12,34, 0-49)
    5.118104, 5.090694, 5.0615, 5.031375, 5.001149, 4.971647, 4.943697, 
    4.918133, 4.895763, 4.877318, 4.863366, 4.854235, 4.849931, 4.850104, 
    4.854072, 4.83257, 4.811661, 4.817543, 4.81448, 4.804032, 4.788081, 
    4.770701, 4.75087, 4.731368, 4.715502, 4.705021, 4.701844, 4.707161, 
    4.721816, 4.74386, 4.770767, 4.803555, 4.838606, 4.873378, 4.905098, 
    4.930877, 4.947974, 4.954234, 4.948682, 4.932118, 4.907397, 4.87913, 
    4.852721, 4.83309, 4.823634, 4.825835, 4.8395, 4.863335, 4.895511, 
    4.934046,
  // momentumX(12,35, 0-49)
    5.113986, 5.086621, 5.057515, 5.027502, 4.997377, 4.967923, 4.939924, 
    4.914174, 4.891447, 4.872436, 4.85766, 4.847354, 4.841359, 4.839027, 
    4.839162, 4.81933, 4.803371, 4.80494, 4.799863, 4.789345, 4.774886, 
    4.761084, 4.745565, 4.731028, 4.720322, 4.714813, 4.715966, 4.724633, 
    4.74135, 4.764152, 4.790324, 4.822191, 4.855091, 4.886513, 4.913769, 
    4.934159, 4.945316, 4.945704, 4.935174, 4.915422, 4.890007, 4.863766, 
    4.841733, 4.827977, 4.824899, 4.833127, 4.851935, 4.879796, 4.914845, 
    4.955168,
  // momentumX(12,36, 0-49)
    5.111942, 5.084561, 5.055326, 5.025081, 4.994619, 4.964703, 4.936105, 
    4.909595, 4.885931, 4.865786, 4.849653, 4.83772, 4.829732, 4.824864, 
    4.821609, 4.804615, 4.794687, 4.792881, 4.786672, 4.776821, 4.764374, 
    4.754197, 4.742932, 4.733154, 4.727239, 4.726232, 4.731174, 4.742603, 
    4.760743, 4.7837, 4.808667, 4.838854, 4.868789, 4.896034, 4.918074, 
    4.932533, 4.937595, 4.932491, 4.91799, 4.896621, 4.872406, 4.850078, 
    4.833977, 4.827167, 4.831044, 4.845499, 4.8694, 4.901079, 4.938695, 
    4.980416,
  // momentumX(12,37, 0-49)
    5.112801, 5.08544, 5.055923, 5.025138, 4.993912, 4.963036, 4.933292, 
    4.905466, 4.880316, 4.858521, 4.840577, 4.826664, 4.81651, 4.809246, 
    4.803285, 4.789212, 4.785302, 4.781154, 4.774646, 4.766088, 4.756061, 
    4.7495, 4.742392, 4.737138, 4.735608, 4.738574, 4.746701, 4.76024, 
    4.779102, 4.801551, 4.82479, 4.852537, 4.878767, 4.901183, 4.917546, 
    4.92596, 4.9253, 4.915676, 4.898742, 4.877671, 4.856634, 4.839904, 
    4.830922, 4.831695, 4.84272, 4.863298, 4.892019, 4.927155, 4.966915, 
    5.009552,
  // momentumX(12,38, 0-49)
    5.117163, 5.089993, 5.060169, 5.028653, 4.996345, 4.964101, 4.932761, 
    4.903154, 4.876072, 4.852218, 4.83211, 4.815961, 4.803544, 4.794055, 
    4.786015, 4.774364, 4.77559, 4.770068, 4.763923, 4.757067, 4.749672, 
    4.746599, 4.743455, 4.742412, 4.744793, 4.75115, 4.761802, 4.776754, 
    4.795622, 4.81691, 4.837911, 4.862556, 4.884535, 4.90178, 4.912446, 
    4.915242, 4.909836, 4.897208, 4.879747, 4.860974, 4.844863, 4.834976, 
    4.833762, 4.842255, 4.86022, 4.886531, 4.919603, 4.957696, 4.999078, 
    5.042069,
  // momentumX(12,39, 0-49)
    5.125264, 5.098615, 5.068628, 5.036368, 5.002841, 4.969013, 4.935816, 
    4.904154, 4.874874, 4.84872, 4.826249, 4.807725, 4.793006, 4.781432, 
    4.771742, 4.761746, 4.766644, 4.760505, 4.755105, 4.750071, 4.74527, 
    4.745384, 4.745862, 4.74859, 4.754327, 4.763429, 4.775914, 4.791576, 
    4.809772, 4.829317, 4.847673, 4.868758, 4.88626, 4.898421, 4.903902, 
    4.902092, 4.893451, 4.879701, 4.863706, 4.849003, 4.839085, 4.836678, 
    4.843287, 4.859147, 4.883482, 4.914883, 4.951668, 4.992102, 5.034494, 
    5.077206,
  // momentumX(12,40, 0-49)
    5.136877, 5.111238, 5.081432, 5.048639, 5.014005, 4.978633, 4.943581, 
    4.909848, 4.878351, 4.849883, 4.825041, 4.804149, 4.787166, 4.773599, 
    4.76246, 4.753274, 4.760116, 4.753808, 4.749212, 4.745819, 4.743309, 
    4.746111, 4.749687, 4.755607, 4.764044, 4.775191, 4.788807, 4.804513, 
    4.821455, 4.83882, 4.854307, 4.871682, 4.884876, 4.892533, 4.893868, 
    4.888951, 4.878927, 4.866021, 4.853262, 4.843918, 4.840827, 4.845891, 
    4.859829, 4.882285, 4.912125, 4.94777, 4.987484, 5.029533, 5.072239, 
    5.113965,
  // momentumX(12,41, 0-49)
    5.151308, 5.127309, 5.098226, 5.065358, 5.030005, 4.993429, 4.956825, 
    4.921301, 4.887843, 4.857288, 4.830274, 4.807172, 4.78804, 4.772555, 
    4.759991, 4.750806, 4.757907, 4.751545, 4.747518, 4.745323, 4.744565, 
    4.749381, 4.755365, 4.763759, 4.774164, 4.786629, 4.800695, 4.81586, 
    4.83112, 4.846073, 4.858711, 4.872571, 4.882043, 4.886209, 4.884839, 
    4.878588, 4.869079, 4.858769, 4.850559, 4.847245, 4.850982, 4.862956, 
    4.883301, 4.911276, 4.945533, 4.98441, 5.026139, 5.068966, 5.111191, 
    5.151146,
  // momentumX(12,42, 0-49)
    5.167433, 5.145825, 5.118198, 5.085958, 5.05056, 5.013422, 4.975871, 
    4.939118, 4.904213, 4.872023, 4.84321, 4.818187, 4.797098, 4.779766, 
    4.765706, 4.755823, 4.761775, 4.755195, 4.751298, 4.749695, 4.749995, 
    4.756035, 4.763631, 4.773695, 4.7853, 4.798368, 4.81227, 4.826428, 
    4.839757, 4.852291, 4.862344, 4.873213, 4.879873, 4.881848, 4.879389, 
    4.873567, 4.866244, 4.859843, 4.856923, 4.859726, 4.86978, 4.887712, 
    4.91327, 4.945491, 4.982934, 5.023899, 5.066599, 5.109246, 5.150087, 
    5.187401,
  // momentumX(12,43, 0-49)
    5.183809, 5.165433, 5.140165, 5.109489, 5.074985, 5.038198, 5.000572, 
    4.963393, 4.927755, 4.894545, 4.864434, 4.837869, 4.815063, 4.795979, 
    4.780333, 4.769211, 4.773004, 4.765872, 4.76158, 4.759906, 4.760523, 
    4.766987, 4.77537, 4.786294, 4.798351, 4.811367, 4.824594, 4.837421, 
    4.848752, 4.859057, 4.866989, 4.875616, 4.880549, 4.881706, 4.879692, 
    4.875801, 4.871909, 4.870196, 4.872773, 4.881325, 4.896852, 4.919589, 
    4.94904, 4.984147, 5.023449, 5.065253, 5.107759, 5.149135, 5.187568, 
    5.22127,
  // momentumX(12,44, 0-49)
    5.198803, 5.184547, 5.162685, 5.134711, 5.102264, 5.066974, 5.03035, 
    4.993721, 4.9582, 4.924677, 4.893834, 4.866149, 4.841905, 4.821187, 
    4.803893, 4.791168, 4.792223, 4.784158, 4.778965, 4.776611, 4.77686, 
    4.783025, 4.79144, 4.802482, 4.814332, 4.826746, 4.838907, 4.85022, 
    4.859634, 4.868042, 4.874416, 4.881635, 4.88592, 4.887495, 4.887174, 
    4.886299, 4.886583, 4.889843, 4.897708, 4.911355, 4.931366, 4.957692, 
    4.989709, 5.026331, 5.066129, 5.10744, 5.148468, 5.187353, 5.222224, 
    5.251262,
  // momentumX(12,45, 0-49)
    5.210752, 5.201502, 5.184183, 5.160196, 5.131147, 5.098663, 5.064255, 
    5.029252, 4.994759, 4.961669, 4.930681, 4.902313, 4.876929, 4.854733, 
    4.835791, 4.821271, 4.819385, 4.810057, 4.803559, 4.800041, 4.799366, 
    4.804659, 4.81249, 4.82304, 4.834153, 4.845552, 4.856387, 4.866125, 
    4.873801, 4.880695, 4.886077, 4.892675, 4.897229, 4.900172, 4.9024, 
    4.905163, 4.909904, 4.918032, 4.9307, 4.948648, 4.972125, 5.000875, 
    5.034193, 5.071006, 5.109934, 5.149368, 5.187541, 5.222595, 5.252655, 
    5.275915,
  // momentumX(12,46, 0-49)
    5.218122, 5.214686, 5.20306, 5.184418, 5.160201, 5.131918, 5.101005, 
    5.068739, 5.036206, 5.004301, 4.973755, 4.945153, 4.91895, 4.895483, 
    4.874975, 4.858628, 4.853901, 4.843082, 4.835012, 4.830008, 4.828019, 
    4.832044, 4.838839, 4.848449, 4.858446, 4.868553, 4.87793, 4.886125, 
    4.892288, 4.898044, 4.902914, 4.909524, 4.915015, 4.919935, 4.925162, 
    4.93177, 4.940877, 4.953484, 4.970314, 4.991725, 5.017685, 5.047775, 
    5.081226, 5.116975, 5.153697, 5.189855, 5.223742, 5.253561, 5.277506, 
    5.293887,
  // momentumX(12,47, 0-49)
    5.21968, 5.222688, 5.21781, 5.205827, 5.18786, 5.16517, 5.139026, 
    5.110605, 5.080956, 5.050987, 5.021486, 4.993125, 4.966475, 4.942011, 
    4.920112, 4.902047, 4.89479, 4.88238, 4.87262, 4.865965, 4.86244, 
    4.86497, 4.870446, 4.87882, 4.88747, 4.896142, 4.904027, 4.910778, 
    4.91566, 4.9206, 4.925312, 4.932374, 4.939193, 4.946368, 4.954691, 
    4.965012, 4.978126, 4.994638, 5.014892, 5.038917, 5.066428, 5.09685, 
    5.129348, 5.162853, 5.19609, 5.227598, 5.255783, 5.278975, 5.295548, 
    5.304067,
  // momentumX(12,48, 0-49)
    5.214645, 5.224436, 5.227116, 5.222918, 5.212476, 5.196669, 5.176497, 
    5.152991, 5.127141, 5.099882, 5.07207, 5.044486, 5.017835, 4.992734, 
    4.969724, 4.950169, 4.940837, 4.926858, 4.91543, 4.907111, 4.90198, 
    4.902931, 4.906935, 4.913908, 4.921101, 4.9283, 4.934745, 4.940191, 
    4.944019, 4.94839, 4.953168, 4.960919, 4.969209, 4.978634, 4.989865, 
    5.003521, 5.020082, 5.039804, 5.062685, 5.088459, 5.11661, 5.146403, 
    5.176918, 5.207063, 5.235599, 5.261165, 5.28232, 5.297623, 5.305756, 
    5.305692,
  // momentumX(12,49, 0-49)
    5.192284, 5.210041, 5.222421, 5.228807, 5.229014, 5.22324, 5.211989, 
    5.195982, 5.176065, 5.153151, 5.128168, 5.102034, 5.075628, 5.049784, 
    5.025281, 5.004552, 5.000236, 4.983833, 4.969202, 4.957649, 4.949624, 
    4.951151, 4.956371, 4.96534, 4.972784, 4.978915, 4.982822, 4.984548, 
    4.983208, 4.98358, 4.985592, 4.994268, 5.004465, 5.016714, 5.031483, 
    5.049073, 5.069549, 5.092734, 5.118204, 5.145324, 5.173291, 5.201159, 
    5.227886, 5.252362, 5.273417, 5.289875, 5.300619, 5.304664, 5.301308, 
    5.290269,
  // momentumX(13,0, 0-49)
    5.302906, 5.297866, 5.283644, 5.261401, 5.232627, 5.198957, 5.162014, 
    5.123312, 5.084203, 5.045848, 5.009209, 4.975058, 4.943973, 4.916348, 
    4.892391, 4.872317, 4.857236, 4.844203, 4.834624, 4.828238, 4.824745, 
    4.82422, 4.826094, 4.830255, 4.836333, 4.844073, 4.853085, 4.862946, 
    4.873157, 4.88348, 4.893552, 4.903595, 4.913329, 4.923114, 4.933573, 
    4.945522, 4.959881, 4.977537, 4.999209, 5.025342, 5.056015, 5.090916, 
    5.129323, 5.170135, 5.211916, 5.252959, 5.291361, 5.325141, 5.352355, 
    5.371239,
  // momentumX(13,1, 0-49)
    5.28951, 5.280722, 5.263025, 5.237669, 5.206186, 5.170209, 5.131349, 
    5.091095, 5.05077, 5.011506, 4.974237, 4.939699, 4.908432, 4.880779, 
    4.856899, 4.837128, 4.823848, 4.810921, 4.801519, 4.795393, 4.792206, 
    4.792432, 4.795098, 4.800194, 4.807179, 4.81584, 4.825731, 4.836394, 
    4.847203, 4.858047, 4.868423, 4.878859, 4.888578, 4.897897, 4.907441, 
    4.918092, 4.930884, 4.946864, 4.966928, 4.991677, 5.021327, 5.055649, 
    5.093979, 5.135242, 5.178015, 5.220617, 5.26118, 5.297764, 5.328457, 
    5.351484,
  // momentumX(13,2, 0-49)
    5.270072, 5.257787, 5.237234, 5.209664, 5.176543, 5.139416, 5.099804, 
    5.059119, 5.018622, 4.979402, 4.942351, 4.90817, 4.877359, 4.850216, 
    4.826835, 4.807679, 4.796417, 4.78367, 4.774438, 4.768469, 4.765407, 
    4.766132, 4.769279, 4.774964, 4.782534, 4.791835, 4.802403, 4.813765, 
    4.825194, 4.836684, 4.847581, 4.858711, 4.868759, 4.877928, 4.886779, 
    4.896184, 4.907245, 4.921134, 4.938916, 4.961381, 4.988906, 5.021394, 
    5.058273, 5.098534, 5.14082, 5.18352, 5.224868, 5.263035, 5.29622, 
    5.322726,
  // momentumX(13,3, 0-49)
    5.246368, 5.230927, 5.208125, 5.179145, 5.145323, 5.108055, 5.068716, 
    5.028602, 4.988883, 4.950584, 4.914549, 4.881436, 4.851695, 4.825564, 
    4.803069, 4.78479, 4.775711, 4.763161, 4.754032, 4.748058, 4.744871, 
    4.745768, 4.749006, 4.754856, 4.762612, 4.77221, 4.783199, 4.795122, 
    4.807179, 4.819442, 4.831099, 4.843277, 4.85408, 4.863536, 4.872057, 
    4.880424, 4.889727, 4.901223, 4.916138, 4.935462, 4.959786, 4.989203, 
    5.023292, 5.061168, 5.10159, 5.143067, 5.183972, 5.222636, 5.257412, 
    5.286727,
  // momentumX(13,4, 0-49)
    5.220337, 5.202127, 5.177616, 5.147886, 5.114111, 5.077507, 5.039276, 
    5.000571, 4.962453, 4.925858, 4.89157, 4.860184, 4.83209, 4.80745, 
    4.786195, 4.768989, 4.762178, 4.749801, 4.740659, 4.734465, 4.730842, 
    4.731516, 4.734381, 4.73989, 4.747362, 4.756843, 4.767935, 4.780223, 
    4.792881, 4.806018, 4.818665, 4.832267, 4.844315, 4.854602, 4.863307, 
    4.871026, 4.878742, 4.887725, 4.899331, 4.91477, 4.934896, 4.960064, 
    4.990092, 5.024294, 5.061602, 5.100693, 5.140108, 5.178351, 5.21394, 
    5.245433,
  // momentumX(13,5, 0-49)
    5.193888, 5.173308, 5.147536, 5.117548, 5.084359, 5.048999, 5.012493, 
    4.975842, 4.939978, 4.905743, 4.873834, 4.84477, 4.818851, 4.796136, 
    4.776439, 4.760425, 4.755842, 4.743599, 4.734304, 4.72764, 4.723233, 
    4.723243, 4.725216, 4.729818, 4.736472, 4.745353, 4.756155, 4.768545, 
    4.781706, 4.795761, 4.809578, 4.824949, 4.838744, 4.850475, 4.860016, 
    4.867673, 4.874217, 4.880829, 4.88893, 4.899941, 4.915029, 4.9349, 
    4.959711, 4.989072, 5.022166, 5.057874, 5.094924, 5.131988, 5.167728, 
    5.200819,
  // momentumX(13,6, 0-49)
    5.168723, 5.146162, 5.119484, 5.089571, 5.057295, 5.023526, 4.989129, 
    4.954954, 4.92181, 4.890425, 4.861399, 4.835148, 4.811861, 4.791458, 
    4.773588, 4.758794, 4.756223, 4.744107, 4.734529, 4.727149, 4.721606, 
    4.720503, 4.721052, 4.724154, 4.729415, 4.737158, 4.74721, 4.759347, 
    4.772826, 4.78774, 4.802809, 4.820201, 4.836185, 4.849976, 4.861088, 
    4.869447, 4.875493, 4.880192, 4.884932, 4.891296, 4.900784, 4.914537, 
    4.933163, 4.956684, 4.984612, 5.016095, 5.050054, 5.085308, 5.12063, 
    5.154777,
  // momentumX(13,7, 0-49)
    5.146191, 5.122014, 5.094694, 5.065038, 5.033816, 5.001769, 4.969636, 
    4.938137, 4.907962, 4.879731, 4.853929, 4.830854, 4.810551, 4.792776, 
    4.776973, 4.763321, 4.762328, 4.750426, 4.740496, 4.732202, 4.72523, 
    4.722604, 4.721231, 4.72226, 4.725554, 4.73159, 4.740366, 4.751813, 
    4.765307, 4.780891, 4.797148, 4.816651, 4.835127, 4.851506, 4.864916, 
    4.874842, 4.881288, 4.884869, 4.886801, 4.888733, 4.892467, 4.899627, 
    4.911375, 4.928267, 4.950256, 4.976807, 5.007057, 5.039953, 5.074344, 
    5.109021,
  // momentumX(13,8, 0-49)
    5.12719, 5.101721, 5.073936, 5.044599, 5.01441, 4.984032, 4.95411, 
    4.92527, 4.898105, 4.873127, 4.850711, 4.831019, 4.81394, 4.799034, 
    4.785518, 4.77283, 4.772757, 4.761313, 4.751078, 4.74178, 4.733187, 
    4.728723, 4.725017, 4.723469, 4.724253, 4.728013, 4.734952, 4.745189, 
    4.758284, 4.7742, 4.791411, 4.812908, 4.833974, 4.853284, 4.869596, 
    4.881938, 4.889804, 4.893339, 4.893427, 4.891637, 4.889973, 4.890526, 
    4.895082, 4.90484, 4.920309, 4.941354, 4.96736, 4.997399, 5.030363, 
    5.06504,
  // momentumX(13,9, 0-49)
    5.112118, 5.085622, 5.057474, 5.028415, 4.999117, 4.970207, 4.94228, 
    4.915903, 4.891597, 4.869787, 4.850737, 4.834479, 4.820738, 4.808884, 
    4.7979, 4.785911, 4.785915, 4.775369, 4.765037, 4.754792, 4.744537, 
    4.73805, 4.731728, 4.727205, 4.725008, 4.725948, 4.730473, 4.738923, 
    4.7511, 4.766879, 4.784646, 4.8078, 4.831308, 4.853636, 4.873232, 
    4.888683, 4.898961, 4.903659, 4.903191, 4.898856, 4.892699, 4.88718, 
    4.884699, 4.887177, 4.895783, 4.910887, 4.932183, 4.958889, 4.989927, 
    5.024058,
  // momentumX(13,10, 0-49)
    5.100892, 5.073568, 5.045088, 5.016195, 4.987566, 4.959826, 4.933566, 
    4.909325, 4.887583, 4.868696, 4.852839, 4.839923, 4.829534, 4.820874, 
    4.812728, 4.801129, 4.800285, 4.791276, 4.781237, 4.770275, 4.758482, 
    4.749933, 4.740851, 4.733079, 4.727515, 4.725141, 4.726683, 4.732738, 
    4.743409, 4.758473, 4.776271, 4.800553, 4.826117, 4.851284, 4.874251, 
    4.893243, 4.906741, 4.913769, 4.914171, 4.908805, 4.899549, 4.88904, 
    4.880201, 4.875673, 4.877369, 4.886271, 4.902476, 4.925397, 4.954008, 
    4.987036,
  // momentumX(13,11, 0-49)
    5.093023, 5.064999, 5.036164, 5.007285, 4.979065, 4.952162, 4.927186, 
    4.904684, 4.885119, 4.868808, 4.855855, 4.846086, 4.838981, 4.833637, 
    4.828726, 4.817231, 4.814683, 4.807994, 4.798809, 4.787527, 4.774482, 
    4.76396, 4.75211, 4.74093, 4.731703, 4.725581, 4.723604, 4.726661, 
    4.7352, 4.748919, 4.766147, 4.790886, 4.817931, 4.845511, 4.87165, 
    4.894293, 4.911518, 4.921821, 4.924446, 4.919686, 4.909037, 4.895079, 
    4.881061, 4.870255, 4.86534, 4.868004, 4.878853, 4.897589, 4.923282, 
    4.954648,
  // momentumX(13,12, 0-49)
    5.087749, 5.05909, 5.029847, 5.00082, 4.972756, 4.946362, 4.92229, 
    4.901118, 4.883312, 4.869174, 4.858771, 4.851879, 4.847934, 4.846014, 
    4.844818, 4.833281, 4.828422, 4.824882, 4.817225, 4.80616, 4.792282, 
    4.779981, 4.765455, 4.75081, 4.737704, 4.727466, 4.721484, 4.720968, 
    4.72675, 4.738482, 4.754528, 4.778989, 4.806825, 4.836215, 4.865081, 
    4.891179, 4.912287, 4.926467, 4.932404, 4.92977, 4.919513, 4.903913, 
    4.886283, 4.870348, 4.859491, 4.856153, 4.861555, 4.875796, 4.898129, 
    4.927302,
  // momentumX(13,13, 0-49)
    5.084192, 5.054919, 5.025204, 4.995886, 4.967764, 4.941601, 4.918097, 
    4.897873, 4.881418, 4.86904, 4.860798, 4.856464, 4.8555, 4.857069, 
    4.860056, 4.848661, 4.84133, 4.84169, 4.836272, 4.826051, 4.811856, 
    4.798031, 4.780994, 4.762904, 4.745772, 4.731121, 4.720706, 4.716094, 
    4.718533, 4.727675, 4.741975, 4.765423, 4.793318, 4.823824, 4.854806, 
    4.883918, 4.908742, 4.927023, 4.936974, 4.937667, 4.929421, 4.914011, 
    4.894545, 4.874947, 4.859157, 4.850342, 4.850424, 4.860008, 4.878631, 
    4.905142,
  // momentumX(13,14, 0-49)
    5.081517, 5.05163, 5.021392, 4.991681, 4.963344, 4.937195, 4.913986, 
    4.89438, 4.878895, 4.867865, 4.861372, 4.85923, 4.860987, 4.865987, 
    4.87346, 4.863003, 4.853669, 4.858477, 4.855946, 4.847213, 4.833271, 
    4.818205, 4.798866, 4.777408, 4.756172, 4.736881, 4.721683, 4.712525, 
    4.7111, 4.717124, 4.729209, 4.750969, 4.778223, 4.809133, 4.841548, 
    4.873077, 4.901201, 4.923458, 4.937708, 4.942506, 4.937534, 4.923936, 
    4.904391, 4.882751, 4.863289, 4.849806, 4.844934, 4.849881, 4.864576, 
    4.888054,
  // momentumX(13,15, 0-49)
    5.079049, 5.048556, 5.017774, 4.987615, 4.958967, 4.932677, 4.909543, 
    4.890262, 4.875388, 4.865291, 4.8601, 4.859703, 4.863788, 4.871943, 
    4.883821, 4.876032, 4.865983, 4.875477, 4.876322, 4.869667, 4.856545, 
    4.840522, 4.819111, 4.794412, 4.769051, 4.744977, 4.724737, 4.710681, 
    4.704965, 4.707441, 4.716984, 4.73648, 4.762472, 4.793127, 4.826293, 
    4.859575, 4.890423, 4.916268, 4.934734, 4.94397, 4.943079, 4.932546, 
    4.914461, 4.892363, 4.870615, 4.853478, 4.844249, 4.844784, 4.855497, 
    4.875701,
  // momentumX(13,16, 0-49)
    5.076357, 5.04529, 5.013985, 4.983371, 4.954356, 4.927814, 4.90456, 
    4.885322, 4.870687, 4.861065, 4.85665, 4.857431, 4.863256, 4.873969, 
    4.889624, 4.887436, 4.878976, 4.892997, 4.897475, 4.893355, 4.881554, 
    4.864819, 4.841561, 4.813771, 4.784333, 4.755423, 4.729992, 4.710805, 
    4.700493, 4.699131, 4.705956, 4.722753, 4.746984, 4.776818, 4.810111, 
    4.844488, 4.877415, 4.906292, 4.928608, 4.942223, 4.945766, 4.939097, 
    4.923651, 4.902481, 4.879802, 4.860133, 4.84732, 4.843862, 4.850718, 
    4.867552,
  // momentumX(13,17, 0-49)
    5.073276, 5.041718, 5.00995, 4.978906, 4.949494, 4.922585, 4.899002, 
    4.879483, 4.864644, 4.854941, 4.850645, 4.851858, 4.858593, 4.870928, 
    4.889231, 4.896774, 4.893412, 4.911368, 4.919476, 4.918165, 4.908042, 
    4.890761, 4.865815, 4.835064, 4.801618, 4.767901, 4.737255, 4.712861, 
    4.697815, 4.692492, 4.696613, 4.710435, 4.732548, 4.761121, 4.794013, 
    4.828882, 4.86324, 4.894509, 4.920127, 4.937771, 4.94571, 4.943258, 
    4.931211, 4.912036, 4.889621, 4.86853, 4.853006, 4.846128, 4.849413, 
    4.862942,
  // momentumX(13,18, 0-49)
    5.069894, 5.037993, 5.005871, 4.974439, 4.94458, 4.917144, 4.89294, 
    4.872707, 4.857082, 4.846572, 4.841537, 4.842215, 4.848804, 4.861626, 
    4.881323, 4.903514, 4.910012, 4.930978, 4.94249, 4.944072, 4.935783, 
    4.917948, 4.891298, 4.857579, 4.820136, 4.781682, 4.745924, 4.716439, 
    4.696753, 4.687572, 4.689219, 4.699979, 4.719781, 4.746784, 4.778859, 
    4.813701, 4.848888, 4.881894, 4.910168, 4.931293, 4.943286, 4.945026, 
    4.936729, 4.920257, 4.899048, 4.877536, 4.860189, 4.850558, 4.850698, 
    4.861127,
  // momentumX(13,19, 0-49)
    5.066533, 5.034526, 5.002198, 4.970406, 4.939985, 4.911748, 4.886477, 
    4.864903, 4.847689, 4.835394, 4.828495, 4.827422, 4.832679, 4.845, 
    4.865422, 4.907155, 4.92915, 4.952248, 4.966908, 4.971374, 4.964861, 
    4.946195, 4.917465, 4.88041, 4.838736, 4.795547, 4.754904, 4.720706, 
    4.696789, 4.684154, 4.683802, 4.691631, 4.709097, 4.734366, 4.765323, 
    4.799715, 4.83519, 4.869302, 4.899551, 4.923498, 4.939002, 4.944619, 
    4.940077, 4.926665, 4.907319, 4.886206, 4.86786, 4.856178, 4.853689, 
    4.861349,
  // momentumX(13,20, 0-49)
    5.062326, 5.029428, 4.996673, 4.965066, 4.935573, 4.909109, 4.88653, 
    4.868585, 4.85582, 4.848474, 4.846332, 4.848631, 4.854045, 4.860835, 
    4.867209, 0, 4.960554, 4.96489, 4.966611, 4.9642, 4.956264, 4.938369, 
    4.913416, 4.881072, 4.843659, 4.803276, 4.763498, 4.72832, 4.70213, 
    4.68676, 4.684481, 4.689006, 4.70359, 4.72649, 4.755638, 4.788839, 
    4.823808, 4.858182, 4.88953, 4.915427, 4.93366, 4.942553, 4.941444, 
    4.931111, 4.913975, 4.893856, 4.875212, 4.86215, 4.857589, 4.862891,
  // momentumX(13,21, 0-49)
    5.05939, 5.026729, 4.99416, 4.962648, 4.9331, 4.906367, 4.883225, 
    4.864333, 4.850152, 4.840854, 4.836205, 4.83551, 4.837572, 4.840788, 
    4.843318, 0, 4.988412, 4.991874, 4.992982, 4.989769, 4.980573, 4.958037, 
    4.92908, 4.892868, 4.851937, 4.808477, 4.766072, 4.728681, 4.700647, 
    4.683903, 4.681386, 4.684261, 4.697501, 4.719358, 4.747776, 4.780595, 
    4.815596, 4.850495, 4.882943, 4.910565, 4.93112, 4.942796, 4.944633, 
    4.936992, 4.921839, 4.902638, 4.883723, 4.869337, 4.862715, 4.865593,
  // momentumX(13,22, 0-49)
    5.056715, 5.024198, 4.991746, 4.960288, 4.930684, 4.903732, 4.880151, 
    4.860536, 4.845291, 4.834549, 4.828082, 4.825235, 4.824912, 4.825584, 
    4.825378, 0, 5.007531, 5.01016, 5.010991, 5.007695, 4.998391, 4.972798, 
    4.941637, 4.903322, 4.860387, 4.814988, 4.770687, 4.731456, 4.701693, 
    4.683507, 4.680566, 4.681566, 4.693231, 4.713815, 4.741263, 4.773442, 
    4.808179, 4.843255, 4.876388, 4.905256, 4.92762, 4.941576, 4.94595, 
    4.940767, 4.927596, 4.90955, 4.890788, 4.875599, 4.867455, 4.868394,
  // momentumX(13,23, 0-49)
    5.054629, 5.022224, 4.989868, 4.958463, 4.928839, 4.901758, 4.877898, 
    4.857814, 4.841877, 4.830197, 4.822548, 4.818313, 4.816451, 4.815497, 
    4.813565, 0, 5.020011, 5.021922, 5.022535, 5.019291, 5.010156, 4.982364, 
    4.949795, 4.910171, 4.86599, 4.819386, 4.773896, 4.733502, 4.702621, 
    4.683495, 4.680393, 4.679896, 4.690282, 4.709814, 4.73644, 4.768047, 
    4.802501, 4.837631, 4.871211, 4.900962, 4.924655, 4.940331, 4.946666, 
    4.94344, 4.931912, 4.914906, 4.89641, 4.880715, 4.871446, 4.870869,
  // momentumX(13,24, 0-49)
    5.053342, 5.021052, 4.988799, 4.957475, 4.927895, 4.900801, 4.876853, 
    4.856582, 4.840339, 4.828224, 4.820012, 4.8151, 4.812484, 4.810732, 
    4.807968, 0, 5.026357, 5.027834, 5.028316, 5.025136, 5.016194, 4.987086, 
    4.953739, 4.913423, 4.868618, 4.821458, 4.775474, 4.734633, 4.703346, 
    4.683897, 4.680958, 4.67964, 4.689296, 4.708194, 4.734291, 4.765488, 
    4.799673, 4.834713, 4.868412, 4.898533, 4.92286, 4.939422, 4.946823, 
    4.944707, 4.934157, 4.91782, 4.899562, 4.883654, 4.873792, 4.872372,
  // momentumX(13,25, 0-49)
    5.052937, 5.020776, 4.988652, 4.957452, 4.927993, 4.901019, 4.877185, 
    4.857019, 4.840869, 4.828824, 4.820656, 4.815761, 4.813137, 4.811367, 
    4.80859, 0, 5.026131, 5.027595, 5.028104, 5.025001, 5.016189, 4.986772, 
    4.953303, 4.912925, 4.868127, 4.821061, 4.775249, 4.73463, 4.703572, 
    4.684343, 4.681725, 4.680303, 4.68982, 4.708557, 4.734481, 4.76551, 
    4.799545, 4.834464, 4.868091, 4.898201, 4.922594, 4.939297, 4.946908, 
    4.945036, 4.934718, 4.918549, 4.900354, 4.884392, 4.874371, 4.872713,
  // momentumX(13,26, 0-49)
    5.053365, 5.021352, 4.989378, 4.958348, 4.92909, 4.902367, 4.878851, 
    4.859085, 4.843421, 4.831948, 4.824425, 4.82023, 4.81834, 4.817324, 
    4.815344, 0, 5.019228, 5.021117, 5.02184, 5.018843, 5.010098, 4.981457, 
    4.948575, 4.908823, 4.864714, 4.818419, 4.773448, 4.7337, 4.703471, 
    4.684952, 4.682744, 4.681938, 4.691911, 4.710961, 4.737072, 4.768174, 
    4.802174, 4.836944, 4.870301, 4.900016, 4.923895, 4.939982, 4.946925, 
    4.944401, 4.933534, 4.917, 4.89867, 4.8828, 4.873055, 4.871789,
  // momentumX(13,27, 0-49)
    5.054453, 5.022583, 4.990769, 4.959939, 4.930949, 4.904599, 4.881593, 
    4.862506, 4.847711, 4.837303, 4.831028, 4.82823, 4.827834, 4.828379, 
    4.828067, 0, 5.005809, 5.008458, 5.00954, 5.006703, 4.998044, 4.971261, 
    4.939735, 4.901355, 4.858659, 4.813832, 4.770372, 4.732119, 4.703287, 
    4.685929, 4.684206, 4.684655, 4.695604, 4.715379, 4.741986, 4.773363, 
    4.807406, 4.841971, 4.874848, 4.903781, 4.926571, 4.941309, 4.946741, 
    4.942723, 4.93059, 4.913219, 4.894607, 4.879008, 4.86998, 4.869713,
  // momentumX(13,28, 0-49)
    5.055897, 5.024127, 4.992451, 4.961824, 4.933147, 4.907266, 4.884938, 
    4.866787, 4.853227, 4.844376, 4.839968, 4.839299, 4.841219, 4.844214, 
    4.846556, 0, 4.986444, 4.989986, 4.991482, 4.988878, 4.980467, 4.956567, 
    4.927253, 4.891089, 4.850602, 4.80798, 4.766706, 4.730566, 4.703684, 
    4.687934, 4.686851, 4.689076, 4.701419, 4.722225, 4.749526, 4.781257, 
    4.815298, 4.849463, 4.8815, 4.909118, 4.930127, 4.942695, 4.945752, 
    4.939439, 4.925432, 4.906913, 4.88804, 4.873039, 4.865275, 4.866679,
  // momentumX(13,29, 0-49)
    5.057277, 5.025501, 4.993886, 4.963425, 4.935068, 4.909718, 4.888201, 
    4.871215, 4.859243, 4.852449, 4.850572, 4.852848, 4.858019, 4.864477, 
    4.870577, 0, 4.960837, 4.965211, 4.967146, 4.96498, 4.957272, 4.937307, 
    4.911318, 4.878489, 4.841214, 4.801627, 4.763185, 4.72964, 4.705064, 
    4.691149, 4.690714, 4.694875, 4.708726, 4.730634, 4.758652, 4.790708, 
    4.824646, 4.858231, 4.889145, 4.915062, 4.933808, 4.943669, 4.943821, 
    4.934777, 4.918635, 4.898928, 4.87997, 4.865904, 4.859822, 4.863319,
  // momentumX(13,30, 0-49)
    5.059418, 5.028654, 4.997622, 4.96715, 4.938057, 4.911136, 4.887138, 
    4.866747, 4.850553, 4.839038, 4.832601, 4.831628, 4.836618, 4.848354, 
    4.867994, 4.90837, 4.928143, 4.951606, 4.967244, 4.973113, 4.968354, 
    4.949694, 4.92203, 4.886323, 4.846043, 4.804104, 4.764419, 4.730797, 
    4.707057, 4.694342, 4.694369, 4.700532, 4.715995, 4.739077, 4.76782, 
    4.800131, 4.833815, 4.866575, 4.896039, 4.919852, 4.935893, 4.942627, 
    4.93956, 4.927652, 4.909478, 4.888913, 4.870369, 4.857808, 4.853965, 
    4.860042,
  // momentumX(13,31, 0-49)
    5.060282, 5.029759, 4.999126, 4.96925, 4.940992, 4.915175, 4.892564, 
    4.873836, 4.859542, 4.850095, 4.845772, 4.846765, 4.85328, 4.865714, 
    4.884841, 4.905748, 4.911053, 4.932447, 4.945031, 4.948086, 4.941575, 
    4.923994, 4.898461, 4.866093, 4.830063, 4.792876, 4.758057, 4.729052, 
    4.709362, 4.699802, 4.701348, 4.710032, 4.727447, 4.751931, 4.781534, 
    4.814127, 4.847456, 4.879147, 4.906764, 4.927947, 4.940672, 4.94366, 
    4.936833, 4.921684, 4.90129, 4.879853, 4.861801, 4.850834, 4.849262, 
    4.857854,
  // momentumX(13,32, 0-49)
    5.060558, 5.030423, 5.000259, 4.970952, 4.943376, 4.918372, 4.896713, 
    4.879066, 4.865955, 4.857725, 4.854555, 4.856493, 4.863556, 4.875896, 
    4.894008, 4.900531, 4.896977, 4.915523, 4.924882, 4.9252, 4.916963, 
    4.900275, 4.876549, 4.847143, 4.815058, 4.782508, 4.752657, 4.728541, 
    4.713242, 4.707185, 4.710644, 4.721965, 4.741295, 4.766997, 4.797129, 
    4.829546, 4.861939, 4.891879, 4.916902, 4.9347, 4.943443, 4.94221, 
    4.931443, 4.913217, 4.891095, 4.869491, 4.85271, 4.844056, 4.845331, 
    4.856855,
  // momentumX(13,33, 0-49)
    5.059862, 5.03015, 5.000467, 4.971692, 4.944696, 4.920317, 4.899325, 
    4.882373, 4.869952, 4.862354, 4.859664, 4.861796, 4.868586, 4.879933, 
    4.896007, 4.893321, 4.885574, 4.900522, 4.906545, 4.904282, 4.894521, 
    4.878765, 4.856861, 4.8304, 4.802221, 4.774295, 4.749418, 4.730218, 
    4.719326, 4.716811, 4.722351, 4.736221, 4.757266, 4.783872, 4.814105, 
    4.845798, 4.876605, 4.904065, 4.925737, 4.939448, 4.943662, 4.93793, 
    4.923305, 4.902457, 4.879358, 4.858486, 4.843853, 4.838239, 4.842885, 
    4.857669,
  // momentumX(13,34, 0-49)
    5.058055, 5.028715, 4.999457, 4.971143, 4.944623, 4.920722, 4.900189, 
    4.883659, 4.871587, 4.864218, 4.861553, 4.863379, 4.869329, 4.879015, 
    4.892175, 4.88469, 4.876192, 4.887134, 4.889908, 4.885369, 4.874451, 
    4.859777, 4.839851, 4.816452, 4.79222, 4.768898, 4.748909, 4.734482, 
    4.727811, 4.728682, 4.736307, 4.752478, 4.774912, 4.802001, 4.831811, 
    4.862161, 4.890678, 4.914915, 4.93252, 4.941554, 4.94089, 4.930667, 
    4.912594, 4.889904, 4.866834, 4.847734, 4.836153, 4.834247, 4.842685, 
    4.860934,
  // momentumX(13,35, 0-49)
    5.055274, 5.02619, 4.997241, 4.969266, 4.943089, 4.919506, 4.899241, 
    4.882901, 4.870915, 4.863482, 4.860535, 4.861737, 4.866537, 4.874239, 
    4.884109, 4.875016, 4.868087, 4.875023, 4.874868, 4.868522, 4.85693, 
    4.843543, 4.825792, 4.805592, 4.785332, 4.766533, 4.751252, 4.741336, 
    4.738557, 4.742521, 4.752098, 4.770198, 4.793586, 4.820644, 4.849438, 
    4.87777, 4.90328, 4.923584, 4.936518, 4.940488, 4.934902, 4.920564, 
    4.899837, 4.876399, 4.854555, 4.838321, 4.830633, 4.832978, 4.845473, 
    4.86724,
  // momentumX(13,36, 0-49)
    5.051935, 5.022963, 4.994163, 4.966357, 4.940342, 4.916883, 4.896673, 
    4.880292, 4.868145, 4.860397, 4.856926, 4.857306, 4.860819, 4.866513, 
    4.873233, 4.864482, 4.860516, 4.863798, 4.861239, 4.853672, 4.841947, 
    4.830064, 4.814686, 4.797793, 4.781472, 4.767046, 4.756203, 4.750443, 
    4.751133, 4.757798, 4.76908, 4.788637, 4.812456, 4.838905, 4.86604, 
    4.891673, 4.9135, 4.929286, 4.937158, 4.935996, 4.925839, 4.908185, 
    4.885969, 4.863123, 4.843789, 4.831448, 4.828336, 4.835277, 4.851907, 
    4.87708,
  // momentumX(13,37, 0-49)
    5.048712, 5.019714, 4.990895, 4.963061, 4.936992, 4.91342, 4.893018, 
    4.876333, 4.863755, 4.855429, 4.851202, 4.850588, 4.852764, 4.856591, 
    4.860627, 4.853176, 4.852786, 4.853034, 4.848742, 4.840593, 4.829271, 
    4.819106, 4.806266, 4.79274, 4.780269, 4.769989, 4.763242, 4.761208, 
    4.764874, 4.773776, 4.78642, 4.806883, 4.830554, 4.855775, 4.880613, 
    4.902925, 4.920528, 4.931437, 4.934191, 4.928248, 4.914334, 4.894584, 
    4.87234, 4.851547, 4.83594, 4.828331, 4.830231, 4.841869, 4.862504, 
    4.890805,
  // momentumX(13,38, 0-49)
    5.046463, 5.017363, 4.988382, 4.960333, 4.933984, 4.910048, 4.889175, 
    4.871894, 4.858581, 4.849375, 4.84412, 4.842312, 4.843084, 4.84521, 
    4.847122, 4.841239, 4.84439, 4.842373, 4.837064, 4.828948, 4.818515, 
    4.810253, 4.800081, 4.789934, 4.781161, 4.774736, 4.771679, 4.772884, 
    4.778982, 4.789603, 4.803183, 4.82395, 4.846866, 4.87026, 4.892232, 
    4.910744, 4.923823, 4.92984, 4.927855, 4.917969, 4.901567, 4.881282, 
    4.860622, 4.843279, 4.832405, 4.830073, 4.83712, 4.853296, 4.877594, 
    4.908586,
  // momentumX(13,39, 0-49)
    5.046107, 5.016935, 4.987735, 4.959342, 4.932527, 4.907993, 4.886375, 
    4.86819, 4.853814, 4.843393, 4.836789, 4.833525, 4.832754, 4.833261, 
    4.833495, 4.82901, 4.835154, 4.83167, 4.826, 4.818432, 4.809279, 
    4.803062, 4.795628, 4.788808, 4.783522, 4.780604, 4.780778, 4.78469, 
    4.79264, 4.804419, 4.818454, 4.838909, 4.860484, 4.881526, 4.900217, 
    4.914691, 4.92329, 4.924838, 4.918981, 4.90646, 4.889201, 4.870115, 
    4.852602, 4.839882, 4.834409, 4.837548, 4.849568, 4.869874, 4.897309, 
    4.930414,
  // momentumX(13,40, 0-49)
    5.048494, 5.019421, 4.990073, 4.961317, 4.933938, 4.90864, 4.886052, 
    4.866689, 4.850931, 4.838945, 4.830641, 4.8256, 4.823055, 4.82189, 
    4.82068, 4.817156, 4.825377, 4.821116, 4.815586, 4.808927, 4.801313, 
    4.797197, 4.792489, 4.788867, 4.786796, 4.786984, 4.789888, 4.795939, 
    4.805148, 4.817516, 4.831503, 4.85106, 4.870792, 4.889106, 4.904329, 
    4.914861, 4.919432, 4.917396, 4.908987, 4.895493, 4.879183, 4.862983, 
    4.84994, 4.842655, 4.842869, 4.851325, 4.86787, 4.891695, 4.921583, 
    4.956109,
  // momentumX(13,41, 0-49)
    5.05427, 5.025635, 4.996369, 4.967378, 4.939467, 4.913352, 4.889659, 
    4.868913, 4.851506, 4.837645, 4.827295, 4.820136, 4.815523, 4.812502, 
    4.809849, 4.806692, 4.81588, 4.811314, 4.806209, 4.800623, 4.794641, 
    4.79257, 4.790468, 4.789821, 4.790624, 4.793467, 4.798572, 4.806185, 
    4.816072, 4.828482, 4.841944, 4.860108, 4.877642, 4.893072, 4.90494, 
    4.911988, 4.913404, 4.909066, 4.899735, 4.887073, 4.87345, 4.861562, 
    4.85393, 4.852476, 4.858293, 4.871628, 4.892047, 4.918634, 4.950186, 
    4.985343,
  // momentumX(13,42, 0-49)
    5.063781, 5.036088, 5.007306, 4.978371, 4.950112, 4.923259, 4.898448, 
    4.876221, 4.856994, 4.841022, 4.828345, 4.818758, 4.811777, 4.806639, 
    4.802362, 4.798909, 4.80793, 4.803259, 4.798624, 4.794068, 4.789628, 
    4.789413, 4.789672, 4.791672, 4.794939, 4.799946, 4.806708, 4.815324, 
    4.825358, 4.837329, 4.84987, 4.866296, 4.881484, 4.894133, 4.903078, 
    4.907446, 4.906895, 4.90178, 4.893241, 4.883102, 4.873612, 4.867048, 
    4.865321, 4.869707, 4.880752, 4.898339, 4.921859, 4.950371, 4.982732, 
    5.017666,
  // momentumX(13,43, 0-49)
    5.077024, 5.050926, 5.02318, 4.994742, 4.966463, 4.939089, 4.913278, 
    4.889596, 4.868496, 4.850291, 4.835114, 4.822883, 4.813281, 4.80576, 
    4.799586, 4.79519, 4.80303, 4.798201, 4.793865, 4.790109, 4.786953, 
    4.788271, 4.790523, 4.794739, 4.799999, 4.80666, 4.814556, 4.823662, 
    4.8334, 4.84456, 4.855913, 4.87045, 4.883365, 4.893603, 4.900323, 
    4.903059, 4.901888, 4.897532, 4.891333, 4.885078, 4.880715, 4.880008, 
    4.884263, 4.894188, 4.909894, 4.931011, 4.956826, 4.986413, 5.018707, 
    5.052526,
  // momentumX(13,44, 0-49)
    5.09363, 5.069897, 5.04386, 5.016483, 4.988629, 4.96107, 4.934496, 
    4.909508, 4.886611, 4.866188, 4.848468, 4.833498, 4.82113, 4.811025, 
    4.802682, 4.796786, 4.802666, 4.797429, 4.793074, 4.789756, 4.787496, 
    4.789924, 4.7937, 4.79963, 4.806377, 4.814182, 4.822727, 4.831895, 
    4.841009, 4.85113, 4.861181, 4.873878, 4.884815, 4.893214, 4.898576, 
    4.900804, 4.900312, 4.898042, 4.895368, 4.893885, 4.895139, 4.900371, 
    4.910341, 4.925292, 4.945001, 4.968908, 4.996238, 5.026088, 5.057459, 
    5.089253,
  // momentumX(13,45, 0-49)
    5.112896, 5.092362, 5.068785, 5.043111, 5.016217, 4.988903, 4.961903, 
    4.935873, 4.911382, 4.88889, 4.868727, 4.851068, 4.835922, 4.823139, 
    4.812431, 4.804618, 4.808037, 4.802051, 4.79729, 4.793986, 4.792167, 
    4.79523, 4.800014, 4.807119, 4.814841, 4.823317, 4.832101, 4.841004, 
    4.8493, 4.858297, 4.867085, 4.878168, 4.887572, 4.894811, 4.899705, 
    4.902462, 4.903721, 4.904501, 4.906074, 4.909746, 4.916643, 4.927522, 
    4.942692, 4.962025, 4.985044, 5.011038, 5.039169, 5.068532, 5.098169, 
    5.127051,
  // momentumX(13,46, 0-49)
    5.133814, 5.117327, 5.096988, 5.073705, 5.048361, 5.021798, 4.994802, 
    4.968101, 4.942336, 4.918055, 4.895684, 4.87552, 4.857718, 4.842292, 
    4.829139, 4.81916, 4.819887, 4.812812, 4.807271, 4.803571, 4.801742, 
    4.80497, 4.81025, 4.818002, 4.826226, 4.834962, 4.843659, 4.852087, 
    4.859497, 4.867418, 4.875102, 4.884908, 4.893291, 4.900041, 4.905254, 
    4.909355, 4.913095, 4.917461, 4.923537, 4.932306, 4.944498, 4.960462, 
    4.980148, 5.003146, 5.028774, 5.056185, 5.084462, 5.112659, 5.139817, 
    5.164942,
  // momentumX(13,47, 0-49)
    5.155118, 5.143477, 5.127144, 5.10696, 5.083807, 5.058568, 5.032099, 
    5.005201, 4.978597, 4.952922, 4.928703, 4.906341, 4.886123, 4.868207, 
    4.85265, 4.840416, 4.838448, 4.830011, 4.823393, 4.818952, 4.816723, 
    4.819705, 4.825018, 4.832941, 4.841257, 4.849924, 4.85831, 4.866159, 
    4.872729, 4.879717, 4.886525, 4.895436, 4.903288, 4.910117, 4.91623, 
    4.922192, 4.928778, 4.936869, 4.947312, 4.960783, 4.977658, 4.997964, 
    5.021375, 5.047264, 5.074781, 5.102951, 5.130748, 5.157147, 5.181139, 
    5.201734,
  // momentumX(13,48, 0-49)
    5.17534, 5.169244, 5.157641, 5.141272, 5.120998, 5.09774, 5.072417, 
    5.045903, 5.019007, 4.992444, 4.966833, 4.942678, 4.920383, 4.900235, 
    4.882427, 4.867987, 4.863477, 4.85351, 4.845624, 4.840209, 4.837288, 
    4.839696, 4.844657, 4.852349, 4.860429, 4.868786, 4.876736, 4.884, 
    4.889857, 4.896114, 4.9023, 4.910675, 4.918396, 4.925701, 4.933056, 
    4.941097, 4.950563, 4.962187, 4.976577, 4.994122, 5.014909, 5.038708, 
    5.064978, 5.092928, 5.121566, 5.149796, 5.176466, 5.200438, 5.22062, 5.236,
  // momentumX(13,49, 0-49)
    5.18919, 5.190837, 5.186273, 5.175988, 5.160712, 5.141308, 5.11869, 
    5.09377, 5.067405, 5.04039, 5.013444, 4.987204, 4.962228, 4.938995, 
    4.917903, 4.901022, 4.900822, 4.888001, 4.877112, 4.869137, 4.864331, 
    4.86836, 4.875689, 4.886596, 4.896372, 4.905116, 4.911828, 4.916348, 
    4.917615, 4.919777, 4.922395, 4.930235, 4.938002, 4.946137, 4.955254, 
    4.966011, 4.979034, 4.994824, 5.013668, 5.035591, 5.060346, 5.087408, 
    5.116018, 5.145223, 5.173903, 5.200845, 5.22479, 5.244488, 5.258783, 
    5.266685,
  // momentumX(14,0, 0-49)
    5.229131, 5.206501, 5.178502, 5.14638, 5.111412, 5.074858, 5.037918, 
    5.001689, 4.967128, 4.935019, 4.905952, 4.880305, 4.858244, 4.839743, 
    4.824595, 4.812624, 4.804584, 4.797328, 4.792109, 4.788625, 4.78663, 
    4.786323, 4.787329, 4.789779, 4.793612, 4.798909, 4.805624, 4.813658, 
    4.822749, 4.832749, 4.84324, 4.854219, 4.865003, 4.875406, 4.885445, 
    4.89538, 4.905724, 4.917185, 4.930576, 4.94668, 4.966119, 4.989237, 
    5.016041, 5.046188, 5.079033, 5.113686, 5.149096, 5.184103, 5.21749, 
    5.247988,
  // momentumX(14,1, 0-49)
    5.207026, 5.182279, 5.152763, 5.119683, 5.084245, 5.047626, 5.010942, 
    4.975212, 4.941328, 4.910021, 4.881835, 4.857101, 4.835941, 4.818269, 
    4.80382, 4.79253, 4.786399, 4.779195, 4.773937, 4.770339, 4.768142, 
    4.767947, 4.769014, 4.771609, 4.775563, 4.781028, 4.787959, 4.796264, 
    4.805616, 4.816019, 4.826934, 4.838686, 4.850087, 4.860837, 4.870841, 
    4.880264, 4.889561, 4.899436, 4.910755, 4.924414, 4.941188, 4.961601, 
    4.985838, 5.013726, 5.044766, 5.078192, 5.113054, 5.148269, 5.182673, 
    5.215027,
  // momentumX(14,2, 0-49)
    5.183304, 5.15703, 5.12666, 5.093325, 5.058139, 5.022183, 4.986475, 
    4.951942, 4.919401, 4.889516, 4.862769, 4.839439, 4.819584, 4.803053, 
    4.789515, 4.779003, 4.774808, 4.767579, 4.762142, 4.758224, 4.755566, 
    4.755175, 4.755948, 4.758294, 4.761974, 4.767229, 4.774033, 4.782334, 
    4.791769, 4.802477, 4.813826, 4.826488, 4.838775, 4.850249, 4.860665, 
    4.870028, 4.878657, 4.887173, 4.896429, 4.907394, 4.921, 4.937978, 
    4.958755, 4.983394, 5.011603, 5.042788, 5.076122, 5.110613, 5.14515, 
    5.178529,
  // momentumX(14,3, 0-49)
    5.159269, 5.132011, 5.101366, 5.068372, 5.034046, 4.999361, 4.965226, 
    4.932481, 4.901851, 4.873924, 4.849108, 4.82761, 4.809415, 4.794293, 
    4.781828, 4.772121, 4.769814, 4.762452, 4.756672, 4.752212, 4.748813, 
    4.747893, 4.747982, 4.749643, 4.752614, 4.757233, 4.763523, 4.771494, 
    4.780782, 4.791656, 4.803401, 4.817072, 4.830497, 4.84309, 4.854418, 
    4.864275, 4.872768, 4.880341, 4.887757, 4.896002, 4.906137, 4.919126, 
    4.935688, 4.956191, 4.980619, 5.008601, 5.039472, 5.072342, 5.106161, 
    5.139763,
  // momentumX(14,4, 0-49)
    5.136073, 5.108289, 5.077836, 5.045656, 5.012658, 4.979708, 4.947617, 
    4.91712, 4.888855, 4.863318, 4.840836, 4.821526, 4.805284, 4.791785, 
    4.780509, 4.771574, 4.771007, 4.763416, 4.75714, 4.751925, 4.747519, 
    4.745743, 4.744758, 4.745288, 4.747094, 4.75062, 4.755964, 4.763226, 
    4.772083, 4.782914, 4.794947, 4.809652, 4.824399, 4.838461, 4.851204, 
    4.862165, 4.871171, 4.878408, 4.884452, 4.890225, 4.896865, 4.905565, 
    4.917366, 4.933001, 4.952807, 4.976699, 5.004219, 5.034612, 5.066907, 
    5.099984,
  // momentumX(14,5, 0-49)
    5.114647, 5.08669, 5.056768, 5.025724, 4.994371, 4.96347, 4.933736, 
    4.905807, 4.880225, 4.857395, 4.837543, 4.82069, 4.806624, 4.794909, 
    4.784913, 4.776653, 4.77757, 4.769712, 4.76284, 4.756712, 4.751087, 
    4.748175, 4.745767, 4.744746, 4.744943, 4.746911, 4.750852, 4.756979, 
    4.765056, 4.775557, 4.787667, 4.803314, 4.819453, 4.835233, 4.849818, 
    4.862471, 4.872696, 4.88035, 4.885726, 4.889578, 4.893041, 4.89748, 
    4.90426, 4.914527, 4.929033, 4.948059, 4.97142, 4.998543, 5.028562, 
    5.060421,
  // momentumX(14,6, 0-49)
    5.095639, 5.06775, 5.038558, 5.008825, 4.979269, 4.950567, 4.923344, 
    4.898149, 4.875429, 4.855488, 4.838451, 4.824225, 4.812485, 4.802677, 
    4.79404, 4.786319, 4.788359, 4.780312, 4.772842, 4.76574, 4.758781, 
    4.754543, 4.750437, 4.747506, 4.745694, 4.74566, 4.747729, 4.752261, 
    4.759154, 4.768952, 4.780826, 4.797183, 4.814626, 4.832209, 4.848913, 
    4.86374, 4.875854, 4.884737, 4.890322, 4.893084, 4.894041, 4.894635, 
    4.896505, 4.901212, 4.909982, 4.923539, 4.942053, 4.9652, 4.992265, 
    5.022275,
  // momentumX(14,7, 0-49)
    5.079382, 5.051685, 5.023293, 4.994893, 4.967136, 4.940629, 4.915915, 
    4.893468, 4.873641, 4.856643, 4.842487, 4.830967, 4.821641, 4.813837, 
    4.806674, 4.799337, 4.802044, 4.794051, 4.786124, 4.778114, 4.769837, 
    4.764191, 4.758224, 4.753119, 4.748968, 4.746531, 4.746279, 4.748741, 
    4.754, 4.762649, 4.773867, 4.790557, 4.809045, 4.82832, 4.847221, 
    4.864514, 4.879047, 4.889917, 4.896648, 4.899345, 4.898779, 4.896335, 
    4.893821, 4.893167, 4.896089, 4.903821, 4.916978, 4.935566, 4.959084, 
    4.986681,
  // momentumX(14,8, 0-49)
    5.065872, 5.038401, 5.01076, 4.983597, 4.95751, 4.933054, 4.910717, 
    4.890898, 4.87387, 4.859747, 4.848433, 4.839616, 4.832747, 4.827052, 
    4.821545, 4.814451, 4.817304, 4.809798, 4.801712, 4.793008, 4.783563, 
    4.776557, 4.76869, 4.761254, 4.754529, 4.749352, 4.746367, 4.746292, 
    4.749443, 4.756443, 4.766504, 4.783024, 4.80213, 4.822789, 4.843732, 
    4.863547, 4.880808, 4.894256, 4.903001, 4.906718, 4.905815, 4.901471, 
    4.895508, 4.890118, 4.887469, 4.889338, 4.896865, 4.91048, 4.92997, 
    4.954655,
  // momentumX(14,9, 0-49)
    5.054821, 5.027532, 5.000518, 4.974404, 4.949765, 4.927123, 4.906926, 
    4.889516, 4.875094, 4.863682, 4.855093, 4.848915, 4.84452, 4.841063, 
    4.837492, 4.83054, 4.83301, 4.826586, 4.818791, 4.809748, 4.799422, 
    4.791223, 4.781535, 4.77173, 4.762289, 4.754117, 4.748044, 4.744996, 
    4.74556, 4.750387, 4.75874, 4.774489, 4.79366, 4.815218, 4.837843, 
    4.859991, 4.880027, 4.896397, 4.907828, 4.913559, 4.913555, 4.908646, 
    4.9005, 4.891405, 4.883876, 4.880214, 4.88213, 4.890561, 4.905677, 
    4.927028,
  // momentumX(14,10, 0-49)
    5.04573, 5.018534, 4.991975, 4.96668, 4.943219, 4.922101, 4.903752, 
    4.888469, 4.876389, 4.867462, 4.861423, 4.857787, 4.855875, 4.854819, 
    4.85357, 4.846726, 4.848333, 4.843694, 4.836761, 4.827849, 4.817042, 
    4.807907, 4.796583, 4.784479, 4.772281, 4.760951, 4.751504, 4.745098, 
    4.742626, 4.744754, 4.750842, 4.765165, 4.783755, 4.805612, 4.829389, 
    4.853467, 4.876074, 4.895433, 4.909956, 4.918473, 4.920488, 4.916383, 
    4.907503, 4.896041, 4.8847, 4.876213, 4.872857, 4.876142, 4.886695, 
    4.904379,
  // momentumX(14,11, 0-49)
    5.038, 5.010782, 4.984499, 4.959789, 4.937232, 4.917344, 4.900531, 
    4.887064, 4.877037, 4.870335, 4.866637, 4.86542, 4.865989, 4.867517, 
    4.869044, 4.862404, 4.862796, 4.860651, 4.855209, 4.846973, 4.836166, 
    4.826419, 4.813724, 4.799486, 4.784587, 4.770025, 4.757013, 4.746933, 
    4.741017, 4.73996, 4.74325, 4.755486, 4.772819, 4.794303, 4.818602, 
    4.844064, 4.868836, 4.890996, 4.908724, 4.92051, 4.925418, 4.923341, 
    4.915177, 4.902844, 4.889031, 4.87675, 4.86878, 4.867208, 4.873197, 
    4.886992,
  // momentumX(14,12, 0-49)
    5.031034, 5.003688, 4.977518, 4.953181, 4.931284, 4.912348, 4.896778, 
    4.884824, 4.876548, 4.871799, 4.870219, 4.871272, 4.8743, 4.878574, 
    4.883319, 4.877185, 4.876233, 4.87719, 4.873849, 4.866863, 4.856576, 
    4.846573, 4.832829, 4.816703, 4.799254, 4.781491, 4.764815, 4.750834, 
    4.741136, 4.736468, 4.736497, 4.746009, 4.761425, 4.781863, 4.806017, 
    4.832239, 4.858638, 4.883218, 4.904005, 4.919235, 4.927595, 4.928498, 
    4.922335, 4.910599, 4.895769, 4.880947, 4.869279, 4.863392, 4.865007, 
    4.874826,
  // momentumX(14,13, 0-49)
    5.024333, 4.99677, 4.970584, 4.946457, 4.925018, 4.906796, 4.892203, 
    4.881479, 4.874665, 4.87159, 4.871881, 4.875025, 4.880433, 4.887527, 
    4.895803, 4.890821, 4.888721, 4.893181, 4.89245, 4.887251, 4.878012, 
    4.868104, 4.853672, 4.835969, 4.816206, 4.795377, 4.775051, 4.757049, 
    4.743318, 4.734697, 4.731096, 4.73732, 4.750211, 4.768974, 4.792344, 
    4.818688, 4.846123, 4.872623, 4.896131, 4.91471, 4.926751, 4.931248, 
    4.928075, 4.918214, 4.903775, 4.887743, 4.873465, 4.864006, 4.861628, 
    4.867535,
  // momentumX(14,14, 0-49)
    5.017553, 4.989715, 4.963422, 4.939384, 4.918242, 4.90054, 4.88669, 
    4.876932, 4.871295, 4.869604, 4.871495, 4.876493, 4.884107, 4.893934, 
    4.905785, 4.903114, 4.900491, 4.908577, 4.910793, 4.907833, 4.900127, 
    4.890634, 4.875879, 4.856959, 4.835193, 4.811535, 4.787686, 4.765656, 
    4.747746, 4.734937, 4.727468, 4.729933, 4.739788, 4.756329, 4.778342, 
    4.804221, 4.832108, 4.85998, 4.88575, 4.90738, 4.923053, 4.931413, 
    4.931864, 4.92485, 4.912005, 4.896032, 4.880286, 4.868128, 4.8623, 
    4.864512,
  // momentumX(14,15, 0-49)
    5.010522, 4.982379, 4.955929, 4.931895, 4.910927, 4.893575, 4.880256, 
    4.871205, 4.866455, 4.865833, 4.869004, 4.875539, 4.885052, 4.897312, 
    4.912402, 4.913854, 4.911866, 4.923392, 4.928685, 4.928277, 4.922505, 
    4.913686, 4.898948, 4.879184, 4.855774, 4.829604, 4.802463, 4.776515, 
    4.754398, 4.737293, 4.725864, 4.724226, 4.730651, 4.744537, 4.764725, 
    4.789639, 4.817448, 4.846156, 4.873679, 4.897934, 4.916968, 4.929162, 
    4.933515, 4.929967, 4.919626, 4.90479, 4.888655, 4.874717, 4.866093, 
    4.864969,
  // momentumX(14,16, 0-49)
    5.003232, 4.974789, 4.948159, 4.924067, 4.903166, 4.886005, 4.872997, 
    4.864381, 4.860195, 4.860283, 4.864339, 4.872, 4.882958, 4.897115, 
    4.91473, 4.922801, 4.923217, 4.937708, 4.946001, 4.948301, 4.94475, 
    4.936777, 4.92233, 4.902053, 4.877351, 4.849022, 4.818892, 4.789238, 
    4.76301, 4.74164, 4.726334, 4.720396, 4.723143, 4.734078, 4.752094, 
    4.775647, 4.802935, 4.831992, 4.860762, 4.887154, 4.909132, 4.924897, 
    4.93313, 4.933318, 4.926054, 4.91317, 4.897569, 4.882729, 4.872013, 
    4.868022,
  // momentumX(14,17, 0-49)
    4.995819, 4.967114, 4.940305, 4.916105, 4.895159, 4.878008, 4.865059, 
    4.856553, 4.85254, 4.852895, 4.857356, 4.865614, 4.877438, 4.892803, 
    4.912023, 4.929695, 4.934912, 4.951701, 4.962767, 4.967796, 4.966612, 
    4.959546, 4.945543, 4.924974, 4.899243, 4.869065, 4.836262, 4.803187, 
    4.773059, 4.747612, 4.728692, 4.718437, 4.717418, 4.725255, 4.740889, 
    4.762807, 4.789228, 4.818224, 4.84777, 4.875792, 4.900223, 4.919144, 
    4.930996, 4.934896, 4.930968, 4.920557, 4.906198, 4.891222, 4.879112, 
    4.872787,
  // momentumX(14,18, 0-49)
    4.988537, 4.959641, 4.932666, 4.9083, 4.887167, 4.869789, 4.856569, 
    4.847752, 4.843416, 4.843479, 4.847744, 4.855983, 4.868048, 4.88397, 
    4.904027, 4.934335, 4.947203, 4.965634, 4.979208, 4.98692, 4.988139, 
    4.981914, 4.968329, 4.947478, 4.920774, 4.888891, 4.85365, 4.81746, 
    4.783762, 4.754593, 4.73253, 4.71814, 4.713455, 4.718208, 4.731387, 
    4.75151, 4.776821, 4.805424, 4.835332, 4.864502, 4.890868, 4.912439, 
    4.927494, 4.934857, 4.934252, 4.926565, 4.913923, 4.899424, 4.88655, 
    4.878451,
  // momentumX(14,19, 0-49)
    4.981731, 4.952747, 4.925626, 4.901007, 4.879478, 4.86154, 4.847589, 
    4.837891, 4.832567, 4.831611, 4.834948, 4.842501, 4.854297, 4.870481, 
    4.891221, 4.936656, 4.959976, 4.979749, 4.995747, 5.00617, 5.009804, 
    5.004245, 4.990828, 4.969369, 4.941361, 4.907585, 4.869937, 4.830897, 
    4.794071, 4.761743, 4.73723, 4.719127, 4.711077, 4.712924, 4.723711, 
    4.741991, 4.766041, 4.793996, 4.823914, 4.853789, 4.881576, 4.90526, 
    4.923007, 4.933437, 4.93594, 4.930997, 4.920331, 4.906754, 4.893658, 
    4.88432,
  // momentumX(14,20, 0-49)
    4.975356, 4.946013, 4.918895, 4.894783, 4.874384, 4.858284, 4.846906, 
    4.840438, 4.838765, 4.841401, 4.847481, 4.8558, 4.864954, 4.87357, 
    4.880587, 0, 4.989855, 4.995119, 5.000073, 5.003455, 5.004048, 4.997201, 
    4.985688, 4.96794, 4.944427, 4.914887, 4.880343, 4.842763, 4.805717, 
    4.771926, 4.745841, 4.724278, 4.712812, 4.711535, 4.719627, 4.735713, 
    4.758105, 4.784973, 4.814407, 4.844437, 4.873043, 4.898208, 4.918039, 
    4.931002, 4.936229, 4.933856, 4.92523, 4.912845, 4.899946, 4.889857,
  // momentumX(14,21, 0-49)
    4.970289, 4.941153, 4.914182, 4.890114, 4.869606, 4.853193, 4.841239, 
    4.833877, 4.830952, 4.831978, 4.836136, 4.842323, 4.849247, 4.85558, 
    4.860119, 0, 5.006929, 5.011988, 5.017016, 5.020457, 5.020889, 5.011185, 
    4.997466, 4.977767, 4.952747, 4.922137, 4.886837, 4.848618, 4.81087, 
    4.776311, 4.749987, 4.726534, 4.71325, 4.710298, 4.716912, 4.731764, 
    4.753213, 4.779468, 4.808661, 4.838869, 4.868112, 4.894393, 4.915797, 
    4.930689, 4.938019, 4.937646, 4.930596, 4.919082, 4.906178, 4.895215,
  // momentumX(14,22, 0-49)
    4.96617, 4.937153, 4.910255, 4.886184, 4.865558, 4.848874, 4.83646, 
    4.828418, 4.824572, 4.824438, 4.827231, 4.831902, 4.837212, 4.841824, 
    4.844385, 0, 5.018405, 5.023205, 5.02841, 5.032224, 5.033048, 5.021325, 
    5.00638, 4.985718, 4.960042, 4.928993, 4.893322, 4.85464, 4.816243, 
    4.780902, 4.754295, 4.728978, 4.713942, 4.709406, 4.71464, 4.728346, 
    4.748909, 4.774562, 4.803468, 4.833735, 4.863416, 4.890533, 4.913163, 
    4.929612, 4.938688, 4.940041, 4.934431, 4.923813, 4.911096, 4.899575,
  // momentumX(14,23, 0-49)
    4.96328, 4.934348, 4.907502, 4.883425, 4.862714, 4.845841, 4.833112, 
    4.824607, 4.820145, 4.819244, 4.821142, 4.824821, 4.829068, 4.832527, 
    4.833734, 0, 5.025937, 5.030453, 5.035746, 5.039857, 5.041064, 5.027761, 
    5.011934, 4.990608, 4.964503, 4.9332, 4.897349, 4.85845, 4.819719, 
    4.783957, 4.757343, 4.730652, 4.714336, 4.708647, 4.712873, 4.725742, 
    4.745659, 4.770877, 4.799579, 4.829896, 4.859901, 4.887634, 4.911168, 
    4.928766, 4.939146, 4.941798, 4.937283, 4.927362, 4.914799, 4.902847,
  // momentumX(14,24, 0-49)
    4.961791, 4.932945, 4.906162, 4.882113, 4.861383, 4.844429, 4.831546, 
    4.822805, 4.81802, 4.816717, 4.818145, 4.821302, 4.824994, 4.827858, 
    4.828371, 0, 5.029955, 5.034287, 5.039621, 5.043921, 5.045398, 5.031094, 
    5.014718, 4.992973, 4.966591, 4.935138, 4.899226, 4.8603, 4.821521, 
    4.785698, 4.759323, 4.731932, 4.714949, 4.708636, 4.712295, 4.724666, 
    4.744171, 4.76908, 4.797589, 4.827847, 4.857946, 4.88594, 4.909908, 
    4.928101, 4.939186, 4.942573, 4.93871, 4.929234, 4.916815, 4.904671,
  // momentumX(14,25, 0-49)
    4.961771, 4.933026, 4.906334, 4.882361, 4.86169, 4.844777, 4.831912, 
    4.823165, 4.818351, 4.816997, 4.818359, 4.821449, 4.825079, 4.827899, 
    4.828384, 0, 5.03003, 5.034381, 5.039783, 5.044186, 5.045787, 5.031203, 
    5.014672, 4.992793, 4.966319, 4.934835, 4.89897, 4.860161, 4.821557, 
    4.785944, 4.759897, 4.732482, 4.715449, 4.709057, 4.712609, 4.724858, 
    4.744236, 4.769025, 4.797433, 4.827615, 4.857674, 4.88567, 4.909687, 
    4.927975, 4.939195, 4.942734, 4.939016, 4.929639, 4.917246, 4.905041,
  // momentumX(14,26, 0-49)
    4.963167, 4.93454, 4.907962, 4.884112, 4.863579, 4.846827, 4.834151, 
    4.825628, 4.821076, 4.820027, 4.821736, 4.825215, 4.829287, 4.832619, 
    4.833757, 0, 5.026039, 5.030636, 5.036156, 5.040594, 5.042174, 5.028095, 
    5.011848, 4.990179, 4.963848, 4.932496, 4.896807, 4.858271, 4.820046, 
    4.784883, 4.759194, 4.73243, 4.715955, 4.710011, 4.713904, 4.726387, 
    4.745905, 4.770749, 4.799131, 4.829207, 4.85908, 4.886809, 4.91048, 
    4.928358, 4.939132, 4.942234, 4.938139, 4.928508, 4.91602, 4.903892,
  // momentumX(14,27, 0-49)
    4.965813, 4.937301, 4.910845, 4.887145, 4.866809, 4.850321, 4.837995, 
    4.829924, 4.825934, 4.825562, 4.828056, 4.832419, 4.837465, 4.841897, 
    4.844372, 0, 5.018102, 5.023104, 5.028753, 5.033145, 5.034584, 5.021748, 
    5.006234, 4.985136, 4.959219, 4.928194, 4.892848, 4.854764, 4.817146, 
    4.782689, 4.757411, 4.731923, 4.71657, 4.711563, 4.716202, 4.729245, 
    4.749143, 4.774192, 4.802603, 4.832528, 4.862057, 4.88924, 4.912171, 
    4.929139, 4.938899, 4.940991, 4.93603, 4.925817, 4.913135, 4.901226,
  // momentumX(14,28, 0-49)
    4.969423, 4.940984, 4.914621, 4.891065, 4.870954, 4.854809, 4.842978, 
    4.835584, 4.832475, 4.833191, 4.836968, 4.842775, 4.849395, 4.855551, 
    4.860049, 0, 5.006672, 5.0121, 5.017801, 5.022041, 5.023263, 5.01228, 
    4.997938, 4.977812, 4.952632, 4.922198, 4.887433, 4.850056, 4.81334, 
    4.779905, 4.755203, 4.731562, 4.717834, 4.714186, 4.719908, 4.733754, 
    4.754178, 4.779477, 4.80786, 4.837467, 4.866374, 4.892624, 4.914323, 
    4.929817, 4.937974, 4.938513, 4.932271, 4.921261, 4.908408, 4.896985,
  // momentumX(14,29, 0-49)
    4.973598, 4.945132, 4.91878, 4.895313, 4.875417, 4.859663, 4.848455, 
    4.841969, 4.840096, 4.842386, 4.848045, 4.855969, 4.864852, 4.873392, 
    4.88053, 0, 4.991336, 4.997087, 5.002714, 5.006726, 5.007765, 4.999115, 
    4.986455, 4.96784, 4.943899, 4.91449, 4.880672, 4.844324, 4.808808, 
    4.776659, 4.752664, 4.731198, 4.719398, 4.717382, 4.724414, 4.739241, 
    4.760315, 4.785926, 4.81427, 4.84347, 4.871576, 4.896624, 4.916734, 
    4.930334, 4.936449, 4.935032, 4.927205, 4.915243, 4.902236, 4.891462,
  // momentumX(14,30, 0-49)
    4.978459, 4.950448, 4.924171, 4.90026, 4.879285, 4.861737, 4.848003, 
    4.838342, 4.832888, 4.831677, 4.83469, 4.841944, 4.853562, 4.869802, 
    4.890952, 4.937116, 4.960141, 4.981357, 4.999086, 5.011297, 5.016665, 
    5.010939, 4.99806, 4.977265, 4.949973, 4.916874, 4.879813, 4.841241, 
    4.804756, 4.772696, 4.748902, 4.729621, 4.719982, 4.719895, 4.728523, 
    4.744562, 4.766439, 4.792431, 4.820715, 4.84939, 4.876489, 4.900041, 
    4.918213, 4.929551, 4.93329, 4.929682, 4.920183, 4.907356, 4.894434, 
    4.88467,
  // momentumX(14,31, 0-49)
    4.983125, 4.955338, 4.929348, 4.905835, 4.885411, 4.868597, 4.85578, 
    4.847207, 4.842966, 4.843014, 4.847225, 4.855464, 4.867691, 4.884041, 
    4.904872, 4.935839, 4.949141, 4.969279, 4.984799, 4.994443, 4.997485, 
    4.991339, 4.978379, 4.958244, 4.932343, 4.901263, 4.86675, 4.83112, 
    4.797772, 4.768725, 4.747015, 4.731064, 4.72435, 4.726704, 4.737257, 
    4.754694, 4.777433, 4.803735, 4.831755, 4.85956, 4.885167, 4.906618, 
    4.922161, 4.930507, 4.931175, 4.92478, 4.913159, 4.899173, 4.886178, 
    4.877337,
  // momentumX(14,32, 0-49)
    4.987358, 4.959856, 4.934148, 4.91095, 4.890905, 4.874556, 4.862307, 
    4.854393, 4.850876, 4.851655, 4.85653, 4.865274, 4.877754, 4.894031, 
    4.914469, 4.932961, 4.939357, 4.958105, 4.971329, 4.978452, 4.979202, 
    4.972534, 4.959299, 4.939528, 4.914677, 4.885373, 4.853353, 4.820845, 
    4.790998, 4.765457, 4.746442, 4.73423, 4.730731, 4.735687, 4.748199, 
    4.766947, 4.790341, 4.816634, 4.843962, 4.870373, 4.893885, 4.912594, 
    4.924883, 4.929708, 4.926944, 4.917631, 4.904008, 4.889196, 4.876601, 
    4.869208,
  // momentumX(14,33, 0-49)
    4.99063, 4.963439, 4.938015, 4.915095, 4.895347, 4.879332, 4.867464, 
    4.859974, 4.856893, 4.858074, 4.863241, 4.872085, 4.88437, 4.900063, 
    4.919447, 4.928698, 4.931004, 4.947732, 4.958413, 4.962972, 4.961474, 
    4.954248, 4.940749, 4.921361, 4.897592, 4.870147, 4.840767, 4.811585, 
    4.785475, 4.763719, 4.747799, 4.739508, 4.739332, 4.746913, 4.761318, 
    4.78121, 4.804995, 4.83091, 4.85707, 4.88152, 4.902306, 4.917626, 
    4.926063, 4.926908, 4.920468, 4.908258, 4.892908, 4.877741, 4.866107, 
    4.860717,
  // momentumX(14,34, 0-49)
    4.992525, 4.96564, 4.940499, 4.917854, 4.898386, 4.882666, 4.871113, 
    4.863943, 4.86116, 4.862561, 4.867793, 4.876443, 4.888147, 4.902713, 
    4.920231, 4.923387, 4.923928, 4.937998, 4.945892, 4.947875, 4.944241, 
    4.936496, 4.92287, 4.90407, 4.881607, 4.856267, 4.829761, 4.804101, 
    4.781861, 4.764022, 4.751439, 4.747082, 4.750193, 4.760307, 4.776446, 
    4.797251, 4.821106, 4.846224, 4.870707, 4.892605, 4.910032, 4.921345, 
    4.92542, 4.921961, 4.911783, 4.896895, 4.880278, 4.865354, 4.855299, 
    4.852454,
  // momentumX(14,35, 0-49)
    4.99278, 4.96617, 4.941314, 4.91896, 4.899793, 4.884388, 4.873153, 
    4.866287, 4.863753, 4.865289, 4.87046, 4.87873, 4.889587, 4.902627, 
    4.917654, 4.917314, 4.917788, 4.928729, 4.933709, 4.933207, 4.927653, 
    4.919489, 4.905965, 4.888046, 4.867195, 4.844253, 4.820849, 4.798853, 
    4.780519, 4.766601, 4.757459, 4.756906, 4.763144, 4.775598, 4.793231, 
    4.814648, 4.838199, 4.862067, 4.884343, 4.903111, 4.916597, 4.923395, 
    4.922756, 4.914888, 4.901155, 4.884047, 4.866805, 4.85282, 4.844973, 
    4.84515,
  // momentumX(14,36, 0-49)
    4.991346, 4.964972, 4.940395, 4.918357, 4.899533, 4.884483, 4.873598, 
    4.867045, 4.864746, 4.866374, 4.871405, 4.879189, 4.889049, 4.900362, 
    4.912611, 4.910634, 4.912133, 4.919724, 4.921842, 4.919075, 4.911914, 
    4.903495, 4.890347, 4.873635, 4.854704, 4.834425, 4.814302, 4.79603, 
    4.781533, 4.77143, 4.765703, 4.768709, 4.777803, 4.792308, 4.811116, 
    4.832782, 4.855612, 4.877761, 4.897319, 4.912441, 4.921529, 4.923491, 
    4.918043, 4.905955, 4.889152, 4.870528, 4.853456, 4.841154, 4.836089, 
    4.839647,
  // momentumX(14,37, 0-49)
    4.988453, 4.962273, 4.937971, 4.916267, 4.897817, 4.883152, 4.872628, 
    4.866377, 4.864271, 4.865924, 4.870734, 4.877946, 4.88674, 4.896296, 
    4.905811, 4.903345, 4.906444, 4.910737, 4.910229, 4.90555, 4.897175, 
    4.888714, 4.876239, 4.86105, 4.844311, 4.826896, 4.810146, 4.795563, 
    4.784745, 4.778251, 4.77579, 4.782004, 4.793592, 4.809768, 4.829356, 
    4.850853, 4.87252, 4.892492, 4.908888, 4.919978, 4.924416, 4.921508, 
    4.911499, 4.895743, 4.87667, 4.857455, 4.841446, 4.831538, 4.829711, 
    4.836845,
  // momentumX(14,38, 0-49)
    4.984639, 4.958626, 4.934591, 4.913228, 4.895154, 4.880854, 4.870646, 
    4.86461, 4.862578, 4.864117, 4.868563, 4.875087, 4.882763, 4.890626, 
    4.897676, 4.89531, 4.900163, 4.901466, 4.898746, 4.892606, 4.88346, 
    4.875215, 4.863713, 4.850336, 4.836003, 4.821574, 4.808197, 4.797181, 
    4.789793, 4.786611, 4.787156, 4.796136, 4.809761, 4.82715, 4.84706, 
    4.867931, 4.887993, 4.905383, 4.918293, 4.92518, 4.925019, 4.917578, 
    4.903661, 4.885168, 4.864916, 4.846192, 4.832146, 4.825239, 4.826932, 
    4.837641,
  // momentumX(14,39, 0-49)
    4.980752, 4.95491, 4.931138, 4.910096, 4.892348, 4.878327, 4.868291, 
    4.862281, 4.86009, 4.861258, 4.865097, 4.870739, 4.877207, 4.88346, 
    4.888396, 4.886341, 4.892785, 4.891613, 4.887215, 4.88012, 4.87067, 
    4.862928, 4.852697, 4.841382, 4.829606, 4.818201, 4.808114, 4.800452, 
    4.796173, 4.795929, 4.799117, 4.810341, 4.825474, 4.843554, 4.863278, 
    4.883053, 4.901103, 4.915614, 4.924913, 4.927712, 4.92337, 4.912158, 
    4.895406, 4.875451, 4.855321, 4.838219, 4.826949, 4.82348, 4.828774, 
    4.842854,
  // momentumX(14,40, 0-49)
    4.977879, 4.952263, 4.928766, 4.908001, 4.890475, 4.876557, 4.866449, 
    4.860152, 4.857441, 4.857857, 4.860724, 4.86519, 4.87028, 4.874952, 
    4.878095, 4.876329, 4.883979, 4.880965, 4.875467, 4.867936, 4.858642, 
    4.851704, 4.843017, 4.833961, 4.824832, 4.816414, 4.809454, 4.804865, 
    4.80331, 4.805566, 4.810947, 4.823834, 4.839893, 4.8581, 4.87712, 
    4.895356, 4.911077, 4.92258, 4.928399, 4.927567, 4.919873, 4.906066, 
    4.88791, 4.868001, 4.849374, 4.834966, 4.827127, 4.827327, 4.836097, 
    4.853168,
  // momentumX(14,41, 0-49)
    4.977243, 4.951975, 4.928784, 4.908237, 4.890777, 4.876709, 4.866188, 
    4.859186, 4.855484, 4.854657, 4.856086, 4.858981, 4.862435, 4.865462, 
    4.867022, 4.865379, 4.873715, 4.869505, 4.863459, 4.855964, 4.84724, 
    4.841386, 4.834473, 4.827814, 4.821355, 4.81582, 4.811758, 4.8099, 
    4.810643, 4.814913, 4.82198, 4.835919, 4.852301, 4.870073, 4.8879, 
    4.904237, 4.91746, 4.92605, 4.928823, 4.925181, 4.915336, 4.900439, 
    4.882529, 4.864255, 4.848449, 4.837637, 4.833674, 4.837571, 4.849523, 
    4.869064,
  // momentumX(14,42, 0-49)
    4.980048, 4.955317, 4.932497, 4.912102, 4.894521, 4.880002, 4.868662, 
    4.860474, 4.855247, 4.852629, 4.852093, 4.852965, 4.854447, 4.855668, 
    4.855711, 4.853931, 4.862373, 4.857519, 4.851374, 4.844295, 4.836475, 
    4.831925, 4.826941, 4.822737, 4.818897, 4.816074, 4.814629, 4.815122, 
    4.817711, 4.823489, 4.831711, 4.846095, 4.862226, 4.879052, 4.895293, 
    4.909513, 4.92027, 4.926304, 4.926771, 4.921447, 4.910919, 4.896608, 
    4.88063, 4.865476, 4.85361, 4.847065, 4.847208, 4.854662, 4.869378, 
    4.89079,
  // momentumX(14,43, 0-49)
    4.987293, 4.963366, 4.941016, 4.920723, 4.902826, 4.887541, 4.874972, 
    4.865113, 4.857836, 4.852889, 4.849873, 4.848258, 4.847405, 4.846586, 
    4.845038, 4.842797, 4.850761, 4.845643, 4.839696, 4.833277, 4.826568, 
    4.82345, 4.820451, 4.818665, 4.817314, 4.816969, 4.817812, 4.820253, 
    4.824242, 4.831039, 4.839899, 4.854184, 4.869569, 4.885051, 4.89946, 
    4.911537, 4.920093, 4.924184, 4.923324, 4.917646, 4.908003, 4.895916, 
    4.88339, 4.872587, 4.865491, 4.863626, 4.867915, 4.878666, 4.895671, 
    4.918324,
  // momentumX(14,44, 0-49)
    4.999643, 4.97684, 4.955107, 4.934894, 4.916515, 4.900183, 4.886018, 
    4.874065, 4.864291, 4.85656, 4.850628, 4.846134, 4.842605, 4.839487, 
    4.83618, 4.833108, 4.840065, 4.83484, 4.82921, 4.823539, 4.818005, 
    4.81632, 4.815243, 4.815725, 4.816647, 4.818492, 4.821272, 4.825261, 
    4.830235, 4.837609, 4.846658, 4.8604, 4.874674, 4.888574, 4.901094, 
    4.911215, 4.918052, 4.921008, 4.91994, 4.915264, 4.907966, 4.899511, 
    4.891633, 4.886055, 4.884239, 4.887223, 4.895544, 4.909267, 4.928077, 
    4.951357,
  // momentumX(14,45, 0-49)
    5.017312, 4.996, 4.97507, 4.95496, 4.935992, 4.918405, 4.902376, 4.88803, 
    4.875444, 4.864624, 4.855481, 4.847826, 4.841365, 4.835716, 4.83044, 
    4.826169, 4.831665, 4.826299, 4.820926, 4.815934, 4.811489, 4.81111, 
    4.811764, 4.814254, 4.81716, 4.820862, 4.825219, 4.830384, 4.835991, 
    4.843586, 4.852475, 4.865373, 4.878339, 4.890605, 4.901376, 4.909918, 
    4.915675, 4.918389, 4.918215, 4.915745, 4.911979, 4.908191, 4.905741, 
    4.90587, 4.909535, 4.917328, 4.92946, 4.945801, 4.965949, 4.989285,
  // momentumX(14,46, 0-49)
    5.040022, 5.0206, 5.000702, 4.98078, 4.9612, 4.942265, 4.924236, 
    4.907354, 4.891817, 4.877773, 4.865296, 4.854357, 4.84483, 4.83649, 
    4.829052, 4.823248, 4.82694, 4.821243, 4.81594, 4.811431, 4.807864, 
    4.808546, 4.810627, 4.814773, 4.819308, 4.82451, 4.8301, 4.836121, 
    4.842098, 4.849669, 4.858179, 4.870093, 4.881728, 4.892483, 4.901812, 
    4.909278, 4.914648, 4.917972, 4.919623, 4.920277, 4.920839, 4.922309, 
    4.92564, 4.931595, 4.94067, 4.953065, 4.968709, 4.987298, 5.008345, 
    5.031216,
  // momentumX(14,47, 0-49)
    5.067022, 5.049904, 5.031317, 5.011751, 4.991643, 4.971396, 4.951393, 
    4.931998, 4.913552, 4.896341, 4.880581, 4.866395, 4.853802, 4.842718, 
    4.832986, 4.825392, 4.827056, 4.820758, 4.815261, 4.810961, 4.807976, 
    4.809393, 4.812525, 4.817905, 4.823682, 4.830026, 4.836539, 4.843167, 
    4.849349, 4.856772, 4.86482, 4.875768, 4.8862, 4.89571, 4.904, 4.910928, 
    4.916553, 4.921173, 4.925306, 4.929629, 4.934891, 4.941786, 4.950864, 
    4.962459, 4.976653, 4.993308, 5.012097, 5.032546, 5.05407, 5.075994,
  // momentumX(14,48, 0-49)
    5.097138, 5.082759, 5.065822, 5.046871, 5.026447, 5.005077, 4.983285, 
    4.961578, 4.940433, 4.920274, 4.901444, 4.884194, 4.868665, 4.854891, 
    4.842824, 4.833281, 4.832807, 4.825633, 4.819666, 4.81528, 4.812549, 
    4.814342, 4.818109, 4.824279, 4.830903, 4.838052, 4.845232, 4.852296, 
    4.858621, 4.86589, 4.873518, 4.883643, 4.893113, 4.901714, 4.90939, 
    4.916262, 4.922637, 4.928999, 4.935947, 4.944109, 4.954046, 4.966163, 
    4.980648, 4.997454, 5.016309, 5.036768, 5.058268, 5.080154, 5.101726, 
    5.122242,
  // momentumX(14,49, 0-49)
    5.131782, 5.121768, 5.107812, 5.090503, 5.070491, 5.048445, 5.025044, 
    5.000954, 4.976798, 4.953141, 4.93047, 4.909184, 4.889575, 4.87183, 
    4.856054, 4.844022, 4.848143, 4.838534, 4.83033, 4.824347, 4.820787, 
    4.825149, 4.832235, 4.842608, 4.852149, 4.861037, 4.868387, 4.874065, 
    4.877024, 4.881012, 4.885324, 4.894529, 4.902976, 4.910685, 4.917894, 
    4.925021, 4.93263, 4.941376, 4.951897, 4.964715, 4.980152, 4.99826, 
    5.018826, 5.04138, 5.065258, 5.08966, 5.113735, 5.1366, 5.15739, 5.175267,
  // momentumX(15,0, 0-49)
    5.116331, 5.087602, 5.057508, 5.02688, 4.99647, 4.966957, 4.938937, 
    4.912934, 4.889373, 4.86856, 4.850661, 4.835689, 4.823497, 4.813806, 
    4.806232, 4.800476, 4.797285, 4.793497, 4.79044, 4.787902, 4.785748, 
    4.784293, 4.783263, 4.78291, 4.783345, 4.784853, 4.787655, 4.791958, 
    4.797826, 4.805394, 4.814459, 4.825126, 4.83667, 4.848646, 4.860583, 
    4.872067, 4.882796, 4.892663, 4.901782, 4.910505, 4.919398, 4.929152, 
    4.940503, 4.954107, 4.970463, 4.989839, 5.012252, 5.037459, 5.064975, 
    5.094105,
  // momentumX(15,1, 0-49)
    5.096625, 5.067094, 5.036662, 5.006133, 4.976219, 4.94755, 4.920673, 
    4.896048, 4.874031, 4.854852, 4.838602, 4.825209, 4.81445, 4.805967, 
    4.799304, 4.794245, 4.792803, 4.788857, 4.785463, 4.782435, 4.779634, 
    4.777761, 4.776192, 4.775315, 4.77516, 4.776093, 4.778361, 4.782217, 
    4.787709, 4.795141, 4.804237, 4.815469, 4.827672, 4.840302, 4.852779, 
    4.864544, 4.87516, 4.884389, 4.892262, 4.899111, 4.905552, 4.912408, 
    4.920602, 4.931015, 4.944372, 4.961137, 4.981477, 5.005255, 5.032047, 
    5.061183,
  // momentumX(15,2, 0-49)
    5.078791, 5.048922, 5.018562, 4.988491, 4.95939, 4.931859, 4.906399, 
    4.883417, 4.863198, 4.845896, 4.831511, 4.819883, 4.810696, 4.803508, 
    4.797784, 4.793371, 4.793595, 4.789402, 4.78556, 4.781904, 4.778296, 
    4.775818, 4.773477, 4.771796, 4.770742, 4.770769, 4.772155, 4.775218, 
    4.780015, 4.787013, 4.795884, 4.807501, 4.820284, 4.833621, 4.846819, 
    4.859183, 4.870113, 4.879212, 4.886373, 4.891838, 4.89621, 4.900389, 
    4.905457, 4.912516, 4.922533, 4.936205, 4.953891, 4.975585, 5.000948, 
    5.029352,
  // momentumX(15,3, 0-49)
    5.06324, 5.033447, 5.003518, 4.974208, 4.946181, 4.920012, 4.896168, 
    4.875008, 4.856752, 4.841472, 4.829074, 4.819304, 4.811752, 4.805884, 
    4.801088, 4.797221, 4.798965, 4.794469, 4.790111, 4.78574, 4.781212, 
    4.777983, 4.774674, 4.771935, 4.769695, 4.768483, 4.768632, 4.770534, 
    4.774281, 4.780493, 4.788819, 4.800562, 4.81377, 4.827785, 4.841828, 
    4.855076, 4.866765, 4.876311, 4.883421, 4.888182, 4.891104, 4.893085, 
    4.895307, 4.899062, 4.905564, 4.915772, 4.93028, 4.949261, 4.972499, 
    4.999438,
  // momentumX(15,4, 0-49)
    5.050073, 5.020701, 4.9915, 4.963202, 4.936454, 4.911811, 4.889717, 
    4.87048, 4.854262, 4.841056, 4.830678, 4.822776, 4.81685, 4.812282, 
    4.808378, 4.804924, 4.807982, 4.803201, 4.798327, 4.79323, 4.787751, 
    4.783697, 4.779289, 4.77529, 4.771614, 4.768863, 4.767426, 4.767785, 
    4.770104, 4.775139, 4.782532, 4.794057, 4.807438, 4.822003, 4.836916, 
    4.851248, 4.864085, 4.874649, 4.88243, 4.887299, 4.88959, 4.890103, 
    4.890029, 4.890785, 4.89381, 4.900341, 4.911246, 4.92694, 4.947388, 
    4.972149,
  // momentumX(15,5, 0-49)
    5.039103, 5.010417, 4.982175, 4.95508, 4.929761, 4.906757, 4.886483, 
    4.869208, 4.855032, 4.843874, 4.835467, 4.829376, 4.825019, 4.821709, 
    4.818674, 4.815492, 4.819603, 4.814657, 4.809369, 4.803624, 4.797256, 
    4.792387, 4.786834, 4.781446, 4.776152, 4.771607, 4.768267, 4.766716, 
    4.767217, 4.770647, 4.77667, 4.787555, 4.800759, 4.81563, 4.831312, 
    4.846801, 4.861059, 4.873127, 4.882268, 4.888099, 4.8907, 4.89067, 
    4.889099, 4.887434, 4.887277, 4.890124, 4.89716, 4.909099, 4.926156, 
    4.948071,
  // momentumX(15,6, 0-49)
    5.029912, 5.00209, 4.974963, 4.949202, 4.925413, 4.904112, 4.885684, 
    4.870354, 4.85817, 4.848981, 4.84245, 4.838074, 4.835212, 4.833121, 
    4.830979, 4.827941, 4.832795, 4.827935, 4.822438, 4.816226, 4.809129, 
    4.803551, 4.796894, 4.790074, 4.783056, 4.776528, 4.771018, 4.767218, 
    4.765527, 4.766914, 4.771096, 4.780854, 4.793445, 4.80827, 4.824483, 
    4.841054, 4.856845, 4.870752, 4.88182, 4.889394, 4.893252, 4.893704, 
    4.891622, 4.888361, 4.885583, 4.885003, 4.888118, 4.895999, 4.909183, 
    4.927671,
  // momentumX(15,7, 0-49)
    5.021935, 4.99507, 4.96914, 4.944782, 4.922575, 4.902999, 4.886406, 
    4.872977, 4.862704, 4.855379, 4.850611, 4.847847, 4.846417, 4.845552, 
    4.844402, 4.841412, 4.846661, 4.84226, 4.836864, 4.83046, 4.822882, 
    4.816778, 4.809143, 4.800937, 4.792175, 4.783555, 4.775673, 4.769339, 
    4.765112, 4.764037, 4.765896, 4.774005, 4.785484, 4.799817, 4.816212, 
    4.833632, 4.850895, 4.866778, 4.880141, 4.89007, 4.896023, 4.897958, 
    4.896429, 4.892569, 4.887981, 4.884502, 4.88391, 4.887653, 4.896658, 
    4.911267,
  // momentumX(15,8, 0-49)
    5.014567, 4.988669, 4.963949, 4.941008, 4.920386, 4.902526, 4.887734, 
    4.876143, 4.867693, 4.862128, 4.859016, 4.857789, 4.857767, 4.858192, 
    4.858227, 4.855232, 4.860509, 4.857036, 4.852131, 4.845875, 4.838133, 
    4.83175, 4.82334, 4.813871, 4.803432, 4.792694, 4.782328, 4.773249, 
    4.766201, 4.762278, 4.76136, 4.767284, 4.777114, 4.790453, 4.806582, 
    4.824496, 4.842996, 4.860787, 4.876583, 4.889243, 4.897914, 4.902189, 
    4.902226, 4.898835, 4.893422, 4.887823, 4.884019, 4.883815, 4.888562, 
    4.899018,
  // momentumX(15,9, 0-49)
    5.007263, 4.982272, 4.958714, 4.937149, 4.918076, 4.901892, 4.888849, 
    4.879029, 4.872319, 4.868426, 4.866897, 4.867163, 4.868573, 4.870416, 
    4.871912, 4.868925, 4.873866, 4.87183, 4.867853, 4.862131, 4.854586, 
    4.848204, 4.83927, 4.828737, 4.816766, 4.803984, 4.791113, 4.779171, 
    4.76909, 4.762001, 4.7579, 4.761126, 4.768773, 4.780583, 4.795938, 
    4.813896, 4.833264, 4.85271, 4.870847, 4.886352, 4.898101, 4.905329, 
    4.907785, 4.905872, 4.900687, 4.893928, 4.887661, 4.883976, 4.884649, 
    4.890883,
  // momentumX(15,10, 0-49)
    4.999604, 4.975416, 4.952922, 4.932649, 4.915052, 4.900475, 4.889113, 
    4.880991, 4.875949, 4.873662, 4.873672, 4.875424, 4.878328, 4.881759, 
    4.885052, 4.882169, 4.886457, 4.886337, 4.883721, 4.878932, 4.87196, 
    4.865866, 4.856699, 4.845355, 4.832079, 4.817416, 4.802129, 4.787311, 
    4.774088, 4.7636, 4.755988, 4.756044, 4.760993, 4.770745, 4.784802, 
    4.802295, 4.822069, 4.84278, 4.862974, 4.881195, 4.896103, 4.906617, 
    4.912094, 4.912504, 4.908549, 4.901665, 4.893864, 4.887411, 4.884446, 
    4.886625,
  // momentumX(15,11, 0-49)
    4.991342, 4.967822, 4.946262, 4.927166, 4.910937, 4.897869, 4.8881, 
    4.881597, 4.878156, 4.877424, 4.878942, 4.882198, 4.886673, 4.891865, 
    4.897288, 4.89474, 4.898158, 4.900331, 4.899464, 4.895978, 4.889944, 
    4.88441, 4.875308, 4.863452, 4.849164, 4.832879, 4.815373, 4.797784, 
    4.781417, 4.767402, 4.756055, 4.752538, 4.754327, 4.761522, 4.773763, 
    4.790272, 4.809944, 4.831436, 4.853266, 4.873887, 4.891792, 4.905651, 
    4.914472, 4.917807, 4.915928, 4.909914, 4.901585, 4.893248, 4.8873, 
    4.885808,
  // momentumX(15,12, 0-49)
    4.982402, 4.959404, 4.938636, 4.920569, 4.905574, 4.893891, 4.885602, 
    4.880623, 4.878705, 4.879471, 4.882472, 4.887239, 4.893341, 4.900425, 
    4.908225, 4.906451, 4.908953, 4.913633, 4.914804, 4.91294, 4.908176, 
    4.903432, 4.894686, 4.88264, 4.867683, 4.850114, 4.830691, 4.810552, 
    4.791155, 4.773605, 4.758424, 4.751015, 4.749251, 4.753448, 4.763399, 
    4.778428, 4.797483, 4.819242, 4.842208, 4.86478, 4.885344, 4.90237, 
    4.914593, 4.92119, 4.922007, 4.917713, 4.90983, 4.900563, 4.892437, 
    4.887838,
  // momentumX(15,13, 0-49)
    4.972854, 4.950241, 4.930109, 4.912913, 4.898992, 4.888544, 4.881598, 
    4.87802, 4.877524, 4.879713, 4.884143, 4.890391, 4.89812, 4.907125, 
    4.917382, 4.917123, 4.918903, 4.926107, 4.929477, 4.929471, 4.926257, 
    4.922477, 4.914348, 4.90243, 4.887171, 4.868714, 4.847758, 4.825398, 
    4.803198, 4.782228, 4.763248, 4.751732, 4.746114, 4.746946, 4.7542, 
    4.767303, 4.785262, 4.806781, 4.830365, 4.854382, 4.877144, 4.897, 
    4.912463, 4.922406, 4.926286, 4.924352, 4.917756, 4.908478, 4.899033, 
    4.892014,
  // momentumX(15,14, 0-49)
    4.96287, 4.940514, 4.920871, 4.904384, 4.891365, 4.881975, 4.876204, 
    4.873875, 4.874665, 4.878159, 4.883919, 4.89156, 4.900823, 4.911641, 
    4.924194, 4.926576, 4.928138, 4.937673, 4.943261, 4.945259, 4.943804, 
    4.941094, 4.933791, 4.922291, 4.907089, 4.888156, 4.866101, 4.841918, 
    4.817236, 4.793077, 4.770475, 4.754752, 4.745088, 4.742292, 4.746523, 
    4.757329, 4.773777, 4.7946, 4.818307, 4.843254, 4.867715, 4.889956, 
    4.908341, 4.921505, 4.928574, 4.929399, 4.924733, 4.916243, 4.906309, 
    4.897605,
  // momentumX(15,15, 0-49)
    4.952686, 4.930484, 4.911194, 4.895252, 4.88295, 4.874424, 4.869629, 
    4.868354, 4.870248, 4.874878, 4.881808, 4.890677, 4.901279, 4.913642, 
    4.92807, 4.93463, 4.936832, 4.948342, 4.95604, 4.960089, 4.960528, 
    4.958922, 4.952585, 4.941731, 4.926888, 4.907864, 4.885134, 4.85956, 
    4.832775, 4.80575, 4.779841, 4.759933, 4.746149, 4.739574, 4.740567, 
    4.748801, 4.763408, 4.783151, 4.806544, 4.831944, 4.857608, 4.881755, 
    4.90265, 4.918758, 4.928937, 4.932689, 4.930367, 4.923283, 4.913586, 
    4.903914,
  // momentumX(15,16, 0-49)
    4.942564, 4.920435, 4.90138, 4.885822, 4.874048, 4.866168, 4.862118, 
    4.86166, 4.864422, 4.869958, 4.877826, 4.887679, 4.899335, 4.912846, 
    4.92854, 4.941131, 4.945195, 4.958213, 4.967833, 4.973904, 4.976303, 
    4.975766, 4.970457, 4.960384, 4.946107, 4.927279, 4.904236, 4.877665, 
    4.849168, 4.819665, 4.790876, 4.766929, 4.749082, 4.738706, 4.736363, 
    4.741861, 4.7544, 4.77277, 4.795497, 4.820938, 4.847348, 4.872924, 
    4.89588, 4.91456, 4.92762, 4.934264, 4.934485, 4.929224, 4.920336, 
    4.910336,
  // momentumX(15,17, 0-49)
    4.932777, 4.910663, 4.891735, 4.876411, 4.864961, 4.857486, 4.853906, 
    4.853971, 4.857299, 4.863437, 4.871946, 4.88248, 4.894852, 4.909085, 
    4.925418, 4.945959, 4.953385, 4.967457, 4.978798, 4.986842, 4.991218, 
    4.991667, 4.987359, 4.978087, 4.964433, 4.945938, 4.922795, 4.895525, 
    4.865663, 4.834091, 4.80294, 4.77522, 4.753508, 4.739446, 4.733802, 
    4.736515, 4.746866, 4.76367, 4.785466, 4.810616, 4.837379, 4.863954, 
    4.888523, 4.909357, 4.924963, 4.934315, 4.937086, 4.933866, 4.926193, 
    4.916392,
  // momentumX(15,18, 0-49)
    4.923589, 4.901454, 4.882562, 4.867312, 4.855964, 4.848607, 4.845161, 
    4.845378, 4.848886, 4.855247, 4.864042, 4.874938, 4.887739, 4.902402, 
    4.918972, 4.949069, 4.961415, 4.976269, 4.989225, 4.999232, 5.005604, 
    5.006928, 5.003522, 4.994929, 4.981759, 4.963496, 4.940249, 4.9124, 
    4.881422, 4.848179, 4.815248, 4.784146, 4.758912, 4.741425, 4.732646, 
    4.732654, 4.740804, 4.755947, 4.776639, 4.801248, 4.828047, 4.855239, 
    4.881002, 4.903563, 4.921335, 4.933104, 4.938289, 4.93716, 4.930946, 
    4.921741,
  // momentumX(15,19, 0-49)
    4.915263, 4.893085, 4.874133, 4.858778, 4.847258, 4.839663, 4.83592, 
    4.835809, 4.838999, 4.845114, 4.853805, 4.864809, 4.877959, 4.89312, 
    4.910018, 4.950513, 4.968981, 4.984726, 4.999439, 5.011564, 5.02004, 
    5.022157, 5.019508, 5.011316, 4.998226, 4.979774, 4.956087, 4.927523, 
    4.895533, 4.860983, 4.826902, 4.792949, 4.764691, 4.744195, 4.732588, 
    4.730083, 4.736119, 4.749599, 4.769093, 4.792991, 4.819576, 4.847066, 
    4.873648, 4.897533, 4.917068, 4.93091, 4.938273, 4.939157, 4.934505, 
    4.926172,
  // momentumX(15,20, 0-49)
    4.908185, 4.886056, 4.867468, 4.852916, 4.84274, 4.837077, 4.835821, 
    4.838592, 4.844738, 4.853366, 4.863411, 4.873747, 4.883327, 4.89133, 
    4.897302, 0, 4.994577, 4.999668, 5.005548, 5.011305, 5.016126, 5.015633, 
    5.013115, 5.006968, 4.997258, 4.982792, 4.962961, 4.937488, 4.907465, 
    4.873701, 4.839848, 4.803802, 4.772908, 4.749545, 4.735105, 4.72999, 
    4.733762, 4.745383, 4.763453, 4.786373, 4.812434, 4.839869, 4.866875, 
    4.891658, 4.912527, 4.928051, 4.937283, 4.939999, 4.936891, 4.929584,
  // momentumX(15,21, 0-49)
    4.90235, 4.880386, 4.861916, 4.847402, 4.837146, 4.831253, 4.829581, 
    4.831733, 4.837054, 4.844685, 4.853627, 4.862837, 4.871323, 4.878238, 
    4.882979, 0, 5.004196, 5.009486, 5.015777, 5.021951, 5.027033, 5.024549, 
    5.020569, 5.013208, 5.002763, 4.988084, 4.968498, 4.943565, 4.914167, 
    4.880956, 4.847917, 4.810899, 4.778774, 4.753971, 4.737977, 4.73131, 
    4.733636, 4.743992, 4.761029, 4.783178, 4.80876, 4.836029, 4.863201, 
    4.888492, 4.910194, 4.926821, 4.937312, 4.941274, 4.939192, 4.932497,
  // momentumX(15,22, 0-49)
    4.897773, 4.875886, 4.857458, 4.842922, 4.832562, 4.826463, 4.824469, 
    4.826171, 4.830924, 4.837883, 4.846084, 4.854511, 4.862186, 4.868207, 
    4.871812, 0, 5.010537, 5.015932, 5.022656, 5.029411, 5.035066, 5.0311, 
    5.026239, 5.01824, 5.007516, 4.992895, 4.973616, 4.949099, 4.920087, 
    4.887161, 4.854692, 4.816629, 4.78334, 4.757275, 4.739974, 4.732033, 
    4.73318, 4.742507, 4.758702, 4.78022, 4.805398, 4.83251, 4.859784, 
    4.885447, 4.907785, 4.925273, 4.936773, 4.941762, 4.940569, 4.934464,
  // momentumX(15,23, 0-49)
    4.894632, 4.872791, 4.854372, 4.839801, 4.829348, 4.823086, 4.820855, 
    4.822244, 4.826617, 4.833141, 4.840868, 4.848798, 4.855937, 4.861334, 
    4.864092, 0, 5.014832, 5.020237, 5.02725, 5.034447, 5.040577, 5.035399, 
    5.029847, 5.021343, 5.010375, 4.995757, 4.976672, 4.952449, 4.923741, 
    4.891075, 4.859142, 4.82031, 4.786209, 4.75929, 4.741114, 4.732311, 
    4.73266, 4.741292, 4.75692, 4.778018, 4.802937, 4.829955, 4.857316, 
    4.883248, 4.906034, 4.924124, 4.93632, 4.94202, 4.941433, 4.935718,
  // momentumX(15,24, 0-49)
    4.89303, 4.871227, 4.852822, 4.83823, 4.827715, 4.821345, 4.818963, 
    4.820161, 4.824309, 4.830588, 4.838061, 4.845731, 4.8526, 4.857682, 4.86, 
    0, 5.017446, 5.022851, 5.03004, 5.037525, 5.043984, 5.038036, 5.032043, 
    5.023195, 5.012022, 4.997339, 4.978312, 4.954233, 4.925709, 4.893244, 
    4.861749, 4.822506, 4.787988, 4.760626, 4.741983, 4.732702, 4.732585, 
    4.740788, 4.756044, 4.776845, 4.801548, 4.828448, 4.855792, 4.881816, 
    4.904807, 4.9232, 4.935774, 4.941876, 4.941653, 4.936192,
  // momentumX(15,25, 0-49)
    4.892978, 4.871228, 4.852853, 4.838268, 4.827735, 4.821324, 4.818879, 
    4.820003, 4.824073, 4.830282, 4.8377, 4.84534, 4.852205, 4.857303, 
    4.859646, 0, 5.017977, 5.023447, 5.030755, 5.038391, 5.045011, 5.03886, 
    5.032743, 5.023767, 5.012475, 4.997696, 4.978612, 4.954521, 4.926036, 
    4.893661, 4.862384, 4.823091, 4.788538, 4.761134, 4.742421, 4.733041, 
    4.732802, 4.74087, 4.755989, 4.776659, 4.801252, 4.828063, 4.855346, 
    4.881342, 4.904335, 4.922764, 4.935397, 4.941571, 4.941417, 4.935998,
  // momentumX(15,26, 0-49)
    4.894406, 4.87272, 4.854392, 4.839842, 4.829338, 4.822953, 4.820543, 
    4.82172, 4.82587, 4.832198, 4.839781, 4.84764, 4.854785, 4.860251, 
    4.863098, 0, 5.016332, 5.021949, 5.029336, 5.036996, 5.043603, 5.037862, 
    5.031976, 5.023129, 5.011848, 4.996982, 4.977752, 4.953513, 4.924929, 
    4.892527, 4.861219, 4.822248, 4.78804, 4.760976, 4.742573, 4.733451, 
    4.733408, 4.741605, 4.756795, 4.777483, 4.802044, 4.828778, 4.855942, 
    4.881776, 4.904565, 4.922753, 4.935126, 4.941044, 4.940664, 4.935086,
  // momentumX(15,27, 0-49)
    4.89715, 4.875522, 4.857244, 4.842745, 4.83231, 4.826026, 4.823761, 
    4.825141, 4.829566, 4.836245, 4.84426, 4.852632, 4.860379, 4.866575, 
    4.870389, 0, 5.012642, 5.018445, 5.025831, 5.033369, 5.039788, 5.035005, 
    5.029674, 5.021203, 5.01006, 4.995123, 4.97568, 4.951184, 4.922391, 
    4.889878, 4.858337, 4.820057, 4.786572, 4.760231, 4.74251, 4.733994, 
    4.734449, 4.743031, 4.758483, 4.779317, 4.80391, 4.830564, 4.857533, 
    4.883053, 4.905414, 4.923075, 4.934859, 4.940183, 4.939286, 4.933345,
  // momentumX(15,28, 0-49)
    4.900956, 4.87935, 4.861095, 4.846647, 4.83631, 4.830202, 4.828211, 
    4.829986, 4.834939, 4.842281, 4.851081, 4.860333, 4.869051, 4.876345, 
    4.881514, 0, 5.007342, 5.013274, 5.020514, 5.02774, 5.033801, 5.030379, 
    5.02587, 5.017995, 5.00712, 4.992149, 4.972463, 4.947652, 4.918607, 
    4.885978, 4.854132, 4.816909, 4.784528, 4.759285, 4.742601, 4.735004, 
    4.736219, 4.745374, 4.761208, 4.782232, 4.806831, 4.833304, 4.85991, 
    4.884882, 4.906523, 4.923325, 4.934174, 4.938588, 4.936932, 4.93051,
  // momentumX(15,29, 0-49)
    4.905488, 4.883822, 4.865526, 4.851095, 4.840873, 4.835017, 4.833459, 
    4.83588, 4.841707, 4.850139, 4.860193, 4.870795, 4.8809, 4.889626, 
    4.896388, 0, 5.000063, 5.005975, 5.012874, 5.019604, 5.025175, 5.023331, 
    5.019852, 5.012797, 5.002379, 4.987502, 4.967638, 4.942543, 4.913272, 
    4.880569, 4.848407, 4.812506, 4.781537, 4.757733, 4.742431, 4.736076, 
    4.738331, 4.748291, 4.764679, 4.786003, 4.810646, 4.836909, 4.86304, 
    4.887277, 4.907935, 4.923557, 4.933121, 4.936285, 4.933587, 4.926498,
  // momentumX(15,30, 0-49)
    4.910488, 4.888827, 4.870213, 4.855021, 4.843503, 4.83578, 4.831827, 
    4.831496, 4.834548, 4.840704, 4.849711, 4.861379, 4.875586, 4.892223, 
    4.911034, 4.954827, 4.973868, 4.991736, 5.008694, 5.022947, 5.033298, 
    5.035358, 5.033057, 5.025144, 5.012241, 4.993824, 4.97003, 4.941264, 
    4.909084, 4.874454, 4.840883, 4.805935, 4.77645, 4.754404, 4.74091, 
    4.73623, 4.739908, 4.750978, 4.768137, 4.789886, 4.814612, 4.84061, 
    4.866129, 4.889415, 4.908816, 4.922949, 4.930926, 4.932596, 4.928713, 
    4.920949,
  // momentumX(15,31, 0-49)
    4.915942, 4.89447, 4.876083, 4.861194, 4.850078, 4.842865, 4.83952, 
    4.839871, 4.843635, 4.850474, 4.860056, 4.872119, 4.886497, 4.903143, 
    4.922074, 4.95497, 4.968733, 4.986028, 5.00144, 5.013679, 5.021948, 
    5.023351, 5.020294, 5.011942, 4.998954, 4.980783, 4.957542, 4.929637, 
    4.898599, 4.865321, 4.832775, 4.800514, 4.773793, 4.754419, 4.743352, 
    4.740744, 4.746068, 4.758324, 4.776205, 4.798216, 4.822738, 4.848071, 
    4.872464, 4.894181, 4.911629, 4.923537, 4.929198, 4.928702, 4.923073, 
    4.914211,
  // momentumX(15,32, 0-49)
    4.921215, 4.899942, 4.881758, 4.8671, 4.856259, 4.849372, 4.846404, 
    4.847165, 4.851349, 4.858582, 4.868499, 4.880802, 4.895323, 4.912056, 
    4.93118, 4.954336, 4.96384, 4.98057, 4.994486, 5.004793, 5.011045, 
    5.011725, 5.007792, 4.99875, 4.985291, 4.966941, 4.943911, 4.916705, 
    4.886889, 4.855299, 4.824359, 4.795338, 4.771907, 4.755643, 4.747331, 
    4.746997, 4.754054, 4.767476, 4.785954, 4.808, 4.832004, 4.856267, 
    4.879059, 4.898688, 4.913652, 4.922843, 4.925797, 4.9229, 4.91548, 
    4.905674,
  // momentumX(15,33, 0-49)
    4.92593, 4.904881, 4.886914, 4.872478, 4.861875, 4.855245, 4.852547, 
    4.853583, 4.858017, 4.865453, 4.875493, 4.887812, 4.902227, 4.91875, 
    4.937635, 4.952839, 4.959489, 4.975294, 4.98753, 4.995835, 5.000043, 
    4.999904, 4.99502, 4.985198, 4.971148, 4.952522, 4.929667, 4.903242, 
    4.874849, 4.845289, 4.816482, 4.7911, 4.771321, 4.758461, 4.753111, 
    4.755168, 4.763979, 4.778497, 4.797407, 4.819228, 4.842355, 4.865105, 
    4.885779, 4.902761, 4.914688, 4.920676, 4.920567, 4.915102, 4.905936, 
    4.895429,
  // momentumX(15,34, 0-49)
    4.929762, 4.908973, 4.891263, 4.877086, 4.866748, 4.860384, 4.857946, 
    4.859209, 4.863815, 4.871333, 4.881327, 4.893431, 4.907422, 4.923276, 
    4.941233, 4.950496, 4.955647, 4.969988, 4.980257, 4.986433, 4.988561, 
    4.987503, 4.981656, 4.971096, 4.956528, 4.937751, 4.915259, 4.889861, 
    4.86318, 4.836005, 4.809812, 4.788346, 4.772446, 4.763155, 4.760866, 
    4.765345, 4.775867, 4.791358, 4.810493, 4.831789, 4.853648, 4.874407, 
    4.892422, 4.906191, 4.914549, 4.916904, 4.913468, 4.905375, 4.89462, 
    4.883753,
  // momentumX(15,35, 0-49)
    4.932462, 4.911976, 4.894581, 4.880731, 4.870724, 4.864684, 4.862538, 
    4.864038, 4.868792, 4.87632, 4.886137, 4.897826, 4.911088, 4.925822, 
    4.942156, 4.947344, 4.952077, 4.964399, 4.972419, 4.976362, 4.976421, 
    4.974379, 4.967628, 4.95648, 4.941605, 4.922957, 4.901151, 4.877123, 
    4.852477, 4.828023, 4.80485, 4.787461, 4.77554, 4.769867, 4.77063, 
    4.777473, 4.789596, 4.805881, 4.824989, 4.845424, 4.865595, 4.883875, 
    4.898703, 4.908737, 4.913075, 4.911485, 4.904602, 4.893983, 4.881938, 
    4.87114,
  // momentumX(15,36, 0-49)
    4.933903, 4.91376, 4.896746, 4.883297, 4.873699, 4.86805, 4.866251, 
    4.868015, 4.872907, 4.880397, 4.889943, 4.901053, 4.91335, 4.926611, 
    4.940794, 4.943399, 4.948446, 4.958294, 4.963863, 4.965548, 4.963623, 
    4.960588, 4.953065, 4.941565, 4.926686, 4.908533, 4.887803, 4.865521, 
    4.843225, 4.821772, 4.801928, 4.788659, 4.780696, 4.778567, 4.782275, 
    4.791337, 4.804873, 4.821717, 4.840497, 4.85971, 4.87777, 4.893103, 
    4.904272, 4.910153, 4.91017, 4.904511, 4.894277, 4.881431, 4.868542, 
    4.858325,
  // momentumX(15,37, 0-49)
    4.934103, 4.914344, 4.897767, 4.884783, 4.875652, 4.870442, 4.86902, 
    4.871055, 4.876065, 4.883467, 4.892656, 4.903069, 4.914239, 4.925816, 
    4.937567, 4.938635, 4.944391, 4.951484, 4.954533, 4.954038, 4.950295, 
    4.946325, 4.938226, 4.926672, 4.912144, 4.894886, 4.875633, 4.855452, 
    4.83577, 4.817514, 4.801187, 4.791965, 4.787823, 4.789057, 4.795502, 
    4.806548, 4.821237, 4.838345, 4.856464, 4.874076, 4.889618, 4.9016, 
    4.908755, 4.910237, 4.905857, 4.896271, 4.883037, 4.868485, 4.855347, 
    4.846265,
  // momentumX(15,38, 0-49)
    4.933275, 4.913924, 4.897812, 4.885321, 4.876671, 4.871897, 4.870824, 
    4.873085, 4.878146, 4.88538, 4.894122, 4.903744, 4.913695, 4.923514, 
    4.932799, 4.932977, 4.93955, 4.943816, 4.944435, 4.941947, 4.936632, 
    4.93186, 4.923436, 4.912159, 4.898354, 4.882379, 4.864967, 4.847182, 
    4.8303, 4.815341, 4.802587, 4.797229, 4.79666, 4.800972, 4.809848, 
    4.822561, 4.83807, 4.855095, 4.872189, 4.887829, 4.900504, 4.908844, 
    4.911808, 4.908888, 4.900332, 4.88727, 4.871682, 4.85616, 4.843473, 
    4.836088,
  // momentumX(15,39, 0-49)
    4.931844, 4.912904, 4.897245, 4.885211, 4.876986, 4.87256, 4.871725, 
    4.874079, 4.879056, 4.885987, 4.894164, 4.902904, 4.911595, 4.919686, 
    4.926654, 4.926291, 4.933585, 4.935168, 4.933599, 4.929408, 4.922832, 
    4.91746, 4.909001, 4.898345, 4.885618, 4.871275, 4.856004, 4.840826, 
    4.826837, 4.815162, 4.805911, 4.804132, 4.80679, 4.813807, 4.824722, 
    4.838705, 4.85464, 4.871191, 4.88689, 4.900232, 4.909787, 4.914362, 
    4.913201, 4.906186, 4.894016, 4.878262, 4.861233, 4.845648, 4.834178, 
    4.828999,
  // momentumX(15,40, 0-49)
    4.930457, 4.911899, 4.896629, 4.884946, 4.876993, 4.872725, 4.87191, 
    4.874125, 4.878788, 4.885204, 4.892647, 4.900396, 4.907799, 4.914251, 
    4.919162, 4.918425, 4.926207, 4.925446, 4.92205, 4.916519, 4.909047, 
    4.903338, 4.895158, 4.885455, 4.874131, 4.861706, 4.848792, 4.836337, 
    4.825235, 4.816731, 4.810798, 4.812224, 4.817683, 4.826947, 4.839435, 
    4.854232, 4.870153, 4.885829, 4.899788, 4.910583, 4.91692, 4.917839, 
    4.912915, 4.902449, 4.887573, 4.870214, 4.852869, 4.838229, 4.828725, 
    4.826172,
  // momentumX(15,41, 0-49)
    4.929952, 4.911724, 4.896721, 4.885202, 4.877274, 4.872872, 4.871749, 
    4.873485, 4.877499, 4.883104, 4.889571, 4.896175, 4.902244, 4.907153, 
    4.910297, 4.909247, 4.917224, 4.914587, 4.909807, 4.903347, 4.895372, 
    4.889627, 4.882048, 4.873604, 4.863957, 4.853662, 4.843232, 4.833522, 
    4.825214, 4.819678, 4.816773, 4.820962, 4.828731, 4.839725, 4.853273, 
    4.868386, 4.883842, 4.898261, 4.910213, 4.918354, 4.921581, 4.919222, 
    4.911222, 4.898285, 4.881907, 4.864242, 4.847815, 4.835123, 4.828254, 
    4.828617,
  // momentumX(15,42, 0-49)
    4.931294, 4.913325, 4.898424, 4.886817, 4.878589, 4.873669, 4.871818, 
    4.872636, 4.875574, 4.879983, 4.885159, 4.890398, 4.895037, 4.898464, 
    4.900094, 4.898733, 4.906603, 4.902615, 4.896917, 4.88995, 4.881868, 
    4.876405, 4.86973, 4.862811, 4.855051, 4.847018, 4.839118, 4.832088, 
    4.826405, 4.823557, 4.823317, 4.829775, 4.83932, 4.851501, 4.865571, 
    4.880503, 4.89507, 4.907923, 4.917725, 4.923294, 4.923772, 4.918811, 
    4.908726, 4.894571, 4.878089, 4.861507, 4.847205, 4.837363, 4.833653, 
    4.837076,
  // momentumX(15,43, 0-49)
    4.935475, 4.917697, 4.902711, 4.890727, 4.881828, 4.875952, 4.872892, 
    4.872292, 4.873665, 4.876423, 4.879921, 4.883506, 4.886554, 4.888489, 
    4.888772, 4.887052, 4.894532, 4.889695, 4.883519, 4.876438, 4.868618, 
    4.863738, 4.85823, 4.853035, 4.847303, 4.841592, 4.836183, 4.831695, 
    4.828406, 4.827918, 4.829926, 4.83814, 4.84892, 4.86174, 4.875812, 
    4.89011, 4.90344, 4.914546, 4.922236, 4.925542, 4.923896, 4.917282, 
    4.906342, 4.892384, 4.877251, 4.863077, 4.851962, 4.845681, 4.845468, 
    4.851949,
  // momentumX(15,44, 0-49)
    4.943389, 4.925753, 4.910508, 4.897867, 4.887924, 4.880651, 4.875891, 
    4.873359, 4.872651, 4.87327, 4.874662, 4.876251, 4.877479, 4.87783, 
    4.876827, 4.87465, 4.881481, 4.876204, 4.869909, 4.863044, 4.855793, 
    4.851745, 4.847598, 4.844251, 4.840609, 4.837198, 4.834173, 4.832032, 
    4.830871, 4.832383, 4.836201, 4.845671, 4.857166, 4.870117, 4.883736, 
    4.897036, 4.908914, 4.918256, 4.924076, 4.925666, 4.922758, 4.91564, 
    4.905199, 4.892863, 4.880429, 4.869793, 4.862683, 4.860432, 4.863861, 
    4.873267,
  // momentumX(15,45, 0-49)
    4.955724, 4.938224, 4.922591, 4.909056, 4.897744, 4.88868, 4.881776, 
    4.876834, 4.873561, 4.871572, 4.870428, 4.86966, 4.868797, 4.867399, 
    4.865062, 4.862271, 4.868221, 4.862769, 4.856599, 4.850181, 4.843715, 
    4.840663, 4.837982, 4.836504, 4.834927, 4.833717, 4.832911, 4.832884, 
    4.833569, 4.836724, 4.841933, 4.852195, 4.863946, 4.876606, 4.889421, 
    4.901495, 4.911865, 4.919618, 4.924015, 4.924632, 4.921483, 4.915091, 
    4.906478, 4.897058, 4.888436, 4.882178, 4.879595, 4.881592, 4.888622, 
    4.900716,
  // momentumX(15,46, 0-49)
    4.972857, 4.955551, 4.939471, 4.924886, 4.911969, 4.900812, 4.891409, 
    4.883674, 4.877432, 4.872438, 4.868383, 4.864922, 4.861692, 4.858339, 
    4.854538, 4.850924, 4.855777, 4.850251, 4.844319, 4.838459, 4.832879, 
    4.830882, 4.82966, 4.82997, 4.830338, 4.831164, 4.832362, 4.834197, 
    4.836456, 4.840928, 4.847151, 4.857822, 4.869471, 4.881536, 4.893338, 
    4.904113, 4.913095, 4.919608, 4.923187, 4.923685, 4.921351, 4.916856, 
    4.911235, 4.905757, 4.901744, 4.900376, 4.902549, 4.908782, 4.91922, 
    4.933684,
  // momentumX(15,47, 0-49)
    4.994822, 4.977833, 4.961337, 4.945648, 4.931002, 4.917567, 4.905441, 
    4.894656, 4.885172, 4.87689, 4.869647, 4.863233, 4.857401, 4.851891, 
    4.846448, 4.841775, 4.845335, 4.839686, 4.833971, 4.828657, 4.82394, 
    4.822939, 4.823054, 4.824963, 4.827073, 4.829704, 4.832666, 4.836111, 
    4.839708, 4.845225, 4.85217, 4.862968, 4.874279, 4.885587, 4.896322, 
    4.905891, 4.913754, 4.9195, 4.922939, 4.92417, 4.923613, 4.921988, 
    4.920238, 4.919398, 4.920445, 4.924166, 4.931067, 4.941337, 4.954875, 
    4.971336,
  // momentumX(15,48, 0-49)
    5.021287, 5.004817, 4.988027, 4.971284, 4.954903, 4.939142, 4.92421, 
    4.910266, 4.897417, 4.885714, 4.875143, 4.865629, 4.857044, 4.849217, 
    4.841962, 4.835991, 4.838085, 4.832155, 4.826528, 4.821638, 4.817649, 
    4.817477, 4.818703, 4.821928, 4.825503, 4.829668, 4.834137, 4.838961, 
    4.843709, 4.850078, 4.857544, 4.868315, 4.879192, 4.88973, 4.899494, 
    4.908081, 4.915195, 4.920693, 4.92464, 4.927336, 4.929301, 4.931226, 
    4.933884, 4.938024, 4.944261, 4.953, 4.964405, 4.978386, 4.994637, 5.01268,
  // momentumX(15,49, 0-49)
    5.058356, 5.043217, 5.026606, 5.00895, 4.990648, 4.972076, 4.953585, 
    4.935503, 4.918123, 4.901687, 4.886375, 4.872292, 4.859453, 4.847805, 
    4.837231, 4.829314, 4.83676, 4.82897, 4.82178, 4.815975, 4.811789, 
    4.814678, 4.819662, 4.827548, 4.834721, 4.8415, 4.847211, 4.851875, 
    4.854626, 4.859023, 4.86429, 4.875, 4.885332, 4.89494, 4.903584, 
    4.911133, 4.917612, 4.923219, 4.928326, 4.933444, 4.939155, 4.946041, 
    4.9546, 4.965176, 4.977912, 4.992743, 5.009426, 5.027546, 5.046576, 
    5.065892,
  // momentumX(16,0, 0-49)
    5.010379, 4.983305, 4.957535, 4.933589, 4.911873, 4.89267, 4.876139, 
    4.862313, 4.851107, 4.842322, 4.835676, 4.830809, 4.827321, 4.824801, 
    4.82285, 4.821224, 4.82087, 4.8188, 4.816489, 4.813863, 4.810887, 
    4.80795, 4.804797, 4.801712, 4.798837, 4.796524, 4.795112, 4.794984, 
    4.796442, 4.799865, 4.805302, 4.813079, 4.822648, 4.833603, 4.845372, 
    4.857257, 4.868512, 4.878438, 4.88649, 4.892384, 4.896164, 4.898243, 
    4.899375, 4.90057, 4.90296, 4.907646, 4.915551, 4.92732, 4.943265, 
    4.963357,
  // momentumX(16,1, 0-49)
    4.998121, 4.971027, 4.945522, 4.922115, 4.901196, 4.88303, 4.86775, 
    4.855347, 4.845687, 4.838506, 4.833449, 4.830081, 4.827929, 4.826505, 
    4.825345, 4.824247, 4.825438, 4.823134, 4.820419, 4.817234, 4.813533, 
    4.810053, 4.806176, 4.802295, 4.798471, 4.795121, 4.792607, 4.79137, 
    4.791726, 4.794225, 4.798886, 4.806432, 4.81596, 4.827044, 4.839068, 
    4.851271, 4.86282, 4.87292, 4.880921, 4.886435, 4.889426, 4.890259, 
    4.889693, 4.888795, 4.888814, 4.891007, 4.896475, 4.906033, 4.920139, 
    4.938877,
  // momentumX(16,2, 0-49)
    4.988944, 4.96211, 4.937086, 4.914367, 4.894336, 4.877245, 4.863204, 
    4.852176, 4.84398, 4.838302, 4.834718, 4.832727, 4.831792, 4.831364, 
    4.830914, 4.830249, 4.832897, 4.830378, 4.827298, 4.8236, 4.819216, 
    4.815224, 4.810616, 4.805884, 4.801012, 4.796468, 4.792636, 4.790017, 
    4.788951, 4.790158, 4.793639, 4.800545, 4.809657, 4.82056, 4.832631, 
    4.845079, 4.857021, 4.867584, 4.876018, 4.881814, 4.884809, 4.885249, 
    4.883801, 4.88151, 4.879666, 4.879637, 4.882692, 4.889841, 4.901728, 
    4.918592,
  // momentumX(16,3, 0-49)
    4.98254, 4.95621, 4.931844, 4.90993, 4.890845, 4.874831, 4.861982, 
    4.852237, 4.845376, 4.841043, 4.838762, 4.837986, 4.838121, 4.838571, 
    4.838752, 4.838411, 4.842396, 4.83975, 4.836403, 4.832302, 4.827349, 
    4.822939, 4.817657, 4.812073, 4.806106, 4.800255, 4.794926, 4.790676, 
    4.787887, 4.787426, 4.789301, 4.795124, 4.80339, 4.813739, 4.82558, 
    4.838131, 4.850492, 4.86174, 4.871041, 4.877756, 4.88156, 4.882516, 
    4.881122, 4.878296, 4.87528, 4.873495, 4.874341, 4.879025, 4.888411, 
    4.902944,
  // momentumX(16,4, 0-49)
    4.978348, 4.952726, 4.929165, 4.908149, 4.890049, 4.875096, 4.863371, 
    4.854793, 4.849114, 4.845946, 4.844783, 4.845037, 4.846092, 4.847313, 
    4.848078, 4.847959, 4.853121, 4.85051, 4.847063, 4.842731, 4.837382, 
    4.832712, 4.826875, 4.8205, 4.813451, 4.806242, 4.799288, 4.793202, 
    4.788418, 4.785934, 4.785778, 4.790048, 4.797011, 4.806389, 4.817661, 
    4.830092, 4.842803, 4.854854, 4.865345, 4.873514, 4.878854, 4.881207, 
    4.880831, 4.878424, 4.875085, 4.872192, 4.871225, 4.873564, 4.880309, 
    4.89215,
  // momentumX(16,5, 0-49)
    4.975636, 4.950883, 4.928251, 4.908212, 4.891126, 4.877218, 4.866553, 
    4.859032, 4.85439, 4.852214, 4.851986, 4.853107, 4.85495, 4.856871, 
    4.858217, 4.858232, 4.864367, 4.862026, 4.858702, 4.854363, 4.848849, 
    4.844121, 4.837903, 4.830859, 4.822809, 4.814256, 4.805618, 4.797554, 
    4.790562, 4.785738, 4.78315, 4.785407, 4.790595, 4.798553, 4.808867, 
    4.820886, 4.833784, 4.84663, 4.858483, 4.868478, 4.87593, 4.880437, 
    4.881971, 4.880943, 4.878209, 4.875005, 4.872805, 4.87311, 4.877246, 
    4.886169,
  // momentumX(16,6, 0-49)
    4.97359, 4.949832, 4.92823, 4.909238, 4.893208, 4.880342, 4.870695, 
    4.864148, 4.860424, 4.859102, 4.859666, 4.861528, 4.864074, 4.866668, 
    4.868656, 4.868736, 4.875587, 4.873809, 4.870874, 4.866787, 4.861371, 
    4.856816, 4.85043, 4.842885, 4.83398, 4.824172, 4.81387, 4.803766, 
    4.794423, 4.787009, 4.781643, 4.781456, 4.784411, 4.790498, 4.799439, 
    4.810699, 4.823528, 4.837036, 4.850263, 4.862264, 4.872192, 4.87941, 
    4.883584, 4.884794, 4.883579, 4.880935, 4.878224, 4.876989, 4.878732, 
    4.884682,
  // momentumX(16,7, 0-49)
    4.971429, 4.948754, 4.928265, 4.910394, 4.895467, 4.883669, 4.87503, 
    4.869415, 4.866539, 4.865985, 4.867253, 4.869784, 4.872997, 4.876294, 
    4.879041, 4.879138, 4.8864, 4.885508, 4.883248, 4.879677, 4.874628, 
    4.870487, 4.864169, 4.856335, 4.846771, 4.835867, 4.824009, 4.811897, 
    4.800161, 4.789993, 4.781582, 4.778574, 4.778876, 4.782658, 4.789808, 
    4.799926, 4.812365, 4.826291, 4.840752, 4.85474, 4.86728, 4.877518, 
    4.884831, 4.888952, 4.890053, 4.888813, 4.886382, 4.88424, 4.883992, 
    4.887099,
  // momentumX(16,8, 0-49)
    4.9685, 4.946961, 4.927648, 4.910966, 4.897206, 4.886523, 4.878919, 
    4.874241, 4.872197, 4.872381, 4.874321, 4.877502, 4.881399, 4.885472, 
    4.889145, 4.889234, 4.896564, 4.896873, 4.895561, 4.892765, 4.888341, 
    4.884839, 4.878826, 4.870933, 4.860958, 4.849187, 4.835968, 4.82198, 
    4.807916, 4.794942, 4.783319, 4.777194, 4.774482, 4.775564, 4.780519, 
    4.789104, 4.800787, 4.814806, 4.83023, 4.846014, 4.861082, 4.874398, 
    4.885083, 4.892534, 4.896551, 4.897444, 4.896061, 4.893718, 4.892021, 
    4.892599,
  // momentumX(16,9, 0-49)
    4.964339, 4.943954, 4.92586, 4.910425, 4.897897, 4.888393, 4.88188, 
    4.878181, 4.876997, 4.87794, 4.88057, 4.88443, 4.889064, 4.894015, 
    4.898808, 4.898908, 4.90595, 4.907724, 4.907599, 4.905803, 4.90224, 
    4.89956, 4.894073, 4.886361, 4.876246, 4.863895, 4.849592, 4.833972, 
    4.817759, 4.802047, 4.787168, 4.777723, 4.771718, 4.769764, 4.772158, 
    4.778826, 4.789371, 4.803106, 4.81913, 4.836383, 4.853708, 4.869932, 
    4.883956, 4.894887, 4.902172, 4.905732, 4.906059, 4.904214, 4.901698, 
    4.900219,
  // momentumX(16,10, 0-49)
    4.958708, 4.939458, 4.922597, 4.908445, 4.897206, 4.888947, 4.88359, 
    4.880938, 4.880676, 4.882433, 4.885808, 4.890401, 4.895841, 4.901774, 
    4.907865, 4.908079, 4.914513, 4.917924, 4.919169, 4.918551, 4.916037, 
    4.914315, 4.909543, 4.902239, 4.892272, 4.879665, 4.864626, 4.847709, 
    4.829641, 4.811388, 4.793344, 4.780487, 4.770998, 4.76575, 4.765265, 
    4.769666, 4.77869, 4.791737, 4.807944, 4.826241, 4.845419, 4.864198, 
    4.881311, 4.895623, 4.906263, 4.912791, 4.915321, 4.914591, 4.911907, 
    4.908954,
  // momentumX(16,11, 0-49)
    4.951579, 4.933411, 4.917763, 4.904904, 4.894985, 4.88802, 4.883884, 
    4.882345, 4.883079, 4.88572, 4.889904, 4.895293, 4.901602, 4.9086, 
    4.916114, 4.916668, 4.922263, 4.927371, 4.930091, 4.930777, 4.929453, 
    4.928766, 4.924852, 4.918157, 4.908612, 4.89609, 4.88071, 4.862903, 
    4.84337, 4.822893, 4.801913, 4.785665, 4.77261, 4.763888, 4.760275, 
    4.762101, 4.769247, 4.781209, 4.797158, 4.816027, 4.836568, 4.857426, 
    4.877209, 4.894594, 4.908454, 4.918019, 4.923042, 4.923909, 4.92166, 
    4.917865,
  // momentumX(16,12, 0-49)
    4.94311, 4.925941, 4.911447, 4.899851, 4.89125, 4.885598, 4.882725, 
    4.882352, 4.884141, 4.887729, 4.892781, 4.899015, 4.906228, 4.914317, 
    4.923285, 4.924597, 4.929274, 4.936002, 4.940219, 4.942276, 4.942241, 
    4.942596, 4.939634, 4.933708, 4.924829, 4.912722, 4.897404, 4.879156, 
    4.858614, 4.836325, 4.812768, 4.793261, 4.776662, 4.764382, 4.757468, 
    4.756468, 4.761423, 4.771923, 4.787184, 4.80614, 4.827521, 4.849919, 
    4.871853, 4.891866, 4.908628, 4.921103, 4.928713, 4.931497, 4.930191, 
    4.926173,
  // momentumX(16,13, 0-49)
    4.933587, 4.917305, 4.903876, 4.893475, 4.886146, 4.881787, 4.880175, 
    4.88099, 4.883869, 4.888443, 4.894396, 4.901491, 4.909599, 4.918728, 
    4.929043, 4.931781, 4.935657, 4.943816, 4.94947, 4.952912, 4.954217, 
    4.955572, 4.953596, 4.948547, 4.940525, 4.92912, 4.914241, 4.895998, 
    4.874925, 4.8513, 4.825628, 4.803096, 4.783074, 4.767251, 4.756944, 
    4.752938, 4.755445, 4.764153, 4.778327, 4.796912, 4.81862, 4.842006, 
    4.865535, 4.887653, 4.906889, 4.921998, 4.932122, 4.936985, 4.937004, 
    4.933322,
  // momentumX(16,14, 0-49)
    4.923371, 4.90785, 4.895366, 4.886055, 4.879909, 4.876776, 4.87638, 
    4.87836, 4.882319, 4.887879, 4.894729, 4.902659, 4.9116, 4.921633, 
    4.933037, 4.938135, 4.941565, 4.95087, 4.957839, 4.962636, 4.965298, 
    4.967563, 4.966561, 4.962437, 4.955395, 4.944908, 4.93078, 4.912937, 
    4.891786, 4.867318, 4.84006, 4.814806, 4.791577, 4.772316, 4.758617, 
    4.751506, 4.751376, 4.758027, 4.770776, 4.788579, 4.810141, 4.833998, 
    4.858574, 4.882263, 4.903494, 4.920869, 4.933316, 4.940278, 4.941876, 
    4.938986,
  // momentumX(16,15, 0-49)
    4.912854, 4.897959, 4.88628, 4.877921, 4.87283, 4.870809, 4.871537, 
    4.874606, 4.87959, 4.886088, 4.893784, 4.90248, 4.912133, 4.922858, 
    4.93496, 4.94358, 4.947157, 4.957278, 4.965407, 4.971506, 4.97552, 
    4.978578, 4.978491, 4.975286, 4.969269, 4.959824, 4.946657, 4.929514, 
    4.908661, 4.883808, 4.855515, 4.827887, 4.801735, 4.779232, 4.762231, 
    4.752002, 4.749129, 4.753531, 4.764589, 4.781275, 4.80229, 4.826159, 
    4.851291, 4.876046, 4.898795, 4.918036, 4.932535, 4.941511, 4.944815, 
    4.943059,
  // momentumX(16,16, 0-49)
    4.902413, 4.888007, 4.876982, 4.869414, 4.865215, 4.864151, 4.865855, 
    4.869885, 4.87578, 4.883116, 4.891562, 4.900916, 4.911123, 4.922285, 
    4.934649, 4.948032, 4.952551, 4.96318, 4.972324, 4.979673, 4.985033, 
    4.98876, 4.989505, 4.98716, 4.982129, 4.973736, 4.961613, 4.945337, 
    4.92504, 4.900175, 4.871372, 4.841729, 4.81299, 4.787511, 4.767387, 
    4.75412, 4.748487, 4.750541, 4.759723, 4.775039, 4.795194, 4.818704, 
    4.843974, 4.86935, 4.893178, 4.913892, 4.930142, 4.940972, 4.946005, 
    4.945608,
  // momentumX(16,17, 0-49)
    4.892386, 4.878341, 4.867813, 4.860855, 4.857354, 4.857041, 4.859523, 
    4.864323, 4.870955, 4.878976, 4.88804, 4.897923, 4.908541, 4.919922, 
    4.932185, 4.951418, 4.957764, 4.968699, 4.978784, 4.987378, 4.994099, 
    4.998383, 4.999869, 4.998282, 4.994113, 4.986661, 4.975505, 4.960099, 
    4.940459, 4.915834, 4.886974, 4.855661, 4.824695, 4.796576, 4.773589, 
    4.757456, 4.749144, 4.748833, 4.756054, 4.769843, 4.78891, 4.811782, 
    4.836864, 4.862501, 4.88703, 4.908854, 4.926551, 4.939031, 4.945736, 
    4.946805,
  // momentumX(16,18, 0-49)
    4.883057, 4.86925, 4.859056, 4.852509, 4.849472, 4.849656, 4.852646, 
    4.857956, 4.865088, 4.873597, 4.88313, 4.893447, 4.904416, 4.91596, 
    4.927983, 4.95368, 4.962641, 4.973895, 4.984979, 4.994907, 5.003065, 
    5.007842, 5.009997, 5.009035, 5.005515, 4.998745, 4.988299, 4.973565, 
    4.954499, 4.930216, 4.901648, 4.868981, 4.836173, 4.805798, 4.780288, 
    4.761552, 4.750729, 4.748141, 4.753402, 4.76559, 4.783442, 4.805486, 
    4.83014, 4.855759, 4.880685, 4.903311, 4.922166, 4.936076, 4.944336, 
    4.946891,
  // momentumX(16,19, 0-49)
    4.874649, 4.860956, 4.850918, 4.844546, 4.841686, 4.842038, 4.845186, 
    4.850657, 4.857982, 4.866745, 4.876626, 4.887396, 4.898871, 4.910821, 
    4.922827, 4.954803, 4.966801, 4.978681, 4.991045, 5.002561, 5.012359, 
    5.017647, 5.020454, 5.019977, 5.016799, 5.010279, 5.000051, 4.985547, 
    4.966752, 4.942739, 4.9147, 4.880971, 4.846727, 4.814543, 4.786932, 
    4.765944, 4.752872, 4.748176, 4.751559, 4.76216, 4.778742, 4.799853, 
    4.823924, 4.849325, 4.874414, 4.897583, 4.917346, 4.932465, 4.942127, 
    4.946119,
  // momentumX(16,20, 0-49)
    4.867816, 4.854584, 4.845321, 4.840126, 4.838893, 4.841312, 4.846864, 
    4.85486, 4.864492, 4.874896, 4.885221, 4.894706, 4.902756, 4.909014, 
    4.913389, 0, 4.987489, 4.991956, 4.99765, 5.003873, 5.010102, 5.012218, 
    5.01397, 5.014071, 5.012827, 5.009157, 5.002196, 4.990902, 4.974914, 
    4.953116, 4.927007, 4.893116, 4.858006, 4.824359, 4.79484, 4.771689, 
    4.756392, 4.749557, 4.751001, 4.759923, 4.775121, 4.79516, 4.818483, 
    4.843477, 4.868512, 4.891992, 4.912422, 4.928527, 4.93941, 4.944731,
  // momentumX(16,21, 0-49)
    4.861976, 4.848943, 4.839874, 4.834837, 4.833697, 4.836112, 4.841539, 
    4.849289, 4.858567, 4.868547, 4.878441, 4.887538, 4.895265, 4.901219, 
    4.905196, 0, 4.992397, 4.997305, 5.003582, 5.010384, 5.017054, 5.017688, 
    5.018337, 5.017498, 5.015707, 5.011953, 5.005382, 4.994881, 4.979984, 
    4.959462, 4.935041, 4.90137, 4.866254, 4.832252, 4.801982, 4.777731, 
    4.761089, 4.752796, 4.752783, 4.760341, 4.774326, 4.793342, 4.815856, 
    4.840277, 4.864996, 4.888429, 4.909086, 4.925674, 4.937243, 4.943362,
  // momentumX(16,22, 0-49)
    4.857375, 4.844437, 4.83546, 4.830493, 4.82939, 4.83179, 4.837147, 
    4.844765, 4.853857, 4.863614, 4.873266, 4.882125, 4.889603, 4.895244, 
    4.898731, 0, 4.995681, 5.000916, 5.007755, 5.015225, 5.022527, 5.022017, 
    5.021948, 5.020552, 5.018504, 5.014805, 5.008574, 4.99863, 4.984444, 
    4.964725, 4.941484, 4.907679, 4.872356, 4.837974, 4.807092, 4.781999, 
    4.764341, 4.754937, 4.753801, 4.760295, 4.773324, 4.791523, 4.813382, 
    4.837328, 4.86177, 4.885137, 4.905946, 4.922899, 4.935011, 4.941789,
  // momentumX(16,23, 0-49)
    4.854089, 4.841188, 4.83224, 4.82729, 4.82618, 4.828554, 4.833859, 
    4.841405, 4.850407, 4.860065, 4.869614, 4.878358, 4.885695, 4.891115, 
    4.894202, 0, 4.998227, 5.003655, 5.010888, 5.018858, 5.026659, 5.025187, 
    5.024527, 5.02266, 5.020362, 5.016635, 5.010581, 5.000975, 4.98724, 
    4.968055, 4.945672, 4.911668, 4.876164, 4.841541, 4.810292, 4.784687, 
    4.76639, 4.756265, 4.754383, 4.760154, 4.772521, 4.790148, 4.811541, 
    4.835138, 4.85936, 4.882646, 4.903519, 4.920674, 4.933112, 4.940302,
  // momentumX(16,24, 0-49)
    4.852131, 4.839238, 4.830288, 4.825319, 4.824179, 4.826513, 4.831777, 
    4.839285, 4.848259, 4.8579, 4.867444, 4.876188, 4.88351, 4.888863, 
    4.891764, 0, 5.000336, 5.005877, 5.013352, 5.021645, 5.029784, 5.027698, 
    5.026659, 5.024476, 5.021976, 5.018165, 5.01214, 5.002656, 4.989122, 
    4.970199, 4.948319, 4.914134, 4.878489, 4.843718, 4.812261, 4.786366, 
    4.767694, 4.757131, 4.754774, 4.760069, 4.771986, 4.789208, 4.810258, 
    4.833585, 4.857615, 4.880801, 4.901666, 4.918907, 4.931514, 4.938937,
  // momentumX(16,25, 0-49)
    4.85146, 4.838564, 4.829591, 4.824589, 4.823408, 4.825703, 4.830941, 
    4.838443, 4.847441, 4.857141, 4.866776, 4.875635, 4.883084, 4.888557, 
    4.891555, 0, 5.001617, 5.00724, 5.014842, 5.023288, 5.03158, 5.02933, 
    5.02819, 5.025898, 5.02329, 5.019381, 5.01327, 5.003716, 4.990139, 
    4.971201, 4.949409, 4.915092, 4.87936, 4.844524, 4.813005, 4.787022, 
    4.768224, 4.757499, 4.754951, 4.760036, 4.771738, 4.788752, 4.809611, 
    4.83277, 4.856662, 4.879742, 4.900535, 4.917737, 4.930336, 4.937777,
  // momentumX(16,26, 0-49)
    4.851977, 4.839075, 4.830077, 4.825035, 4.82382, 4.826095, 4.831341, 
    4.838893, 4.847992, 4.857843, 4.867679, 4.876782, 4.884514, 4.890315, 
    4.893711, 0, 5.001983, 5.007671, 5.015292, 5.023718, 5.031972, 5.030043, 
    5.029104, 5.026941, 5.024355, 5.020361, 5.014077, 5.004286, 4.990434, 
    4.971213, 4.949087, 4.914718, 4.878968, 4.844158, 4.812709, 4.786823, 
    4.768129, 4.757494, 4.755009, 4.760123, 4.771822, 4.788801, 4.809599, 
    4.832676, 4.856466, 4.87942, 4.900066, 4.917099, 4.929512, 4.936756,
  // momentumX(16,27, 0-49)
    4.853549, 4.84063, 4.831599, 4.826528, 4.825302, 4.827601, 4.832926, 
    4.840624, 4.849943, 4.860089, 4.870278, 4.879788, 4.887972, 4.894296, 
    4.898354, 0, 5.001553, 5.007257, 5.014753, 5.022965, 5.030978, 5.02979, 
    5.029314, 5.027491, 5.025039, 5.020969, 5.014422, 5.00423, 4.989888, 
    4.970133, 4.947292, 4.912957, 4.877278, 4.842611, 4.811395, 4.785818, 
    4.767478, 4.757198, 4.755036, 4.760416, 4.772312, 4.789418, 4.810269, 
    4.833325, 4.857021, 4.879806, 4.900201, 4.916908, 4.928932, 4.935752,
  // momentumX(16,28, 0-49)
    4.855995, 4.843037, 4.833967, 4.828879, 4.827681, 4.830082, 4.835604, 
    4.843608, 4.853339, 4.863991, 4.874754, 4.884873, 4.89369, 4.900697, 
    4.905574, 0, 5.000744, 5.006339, 5.013515, 5.021286, 5.028846, 5.028683, 
    5.02886, 5.027533, 5.025298, 5.021149, 5.014251, 5.003506, 4.988485, 
    4.967993, 4.944139, 4.909925, 4.874425, 4.840048, 4.809262, 4.78423, 
    4.766501, 4.756835, 4.75523, 4.761073, 4.773315, 4.790642, 4.811593, 
    4.834626, 4.858176, 4.88069, 4.900694, 4.916894, 4.928325, 4.934512,
  // momentumX(16,29, 0-49)
    4.859104, 4.846059, 4.836926, 4.831833, 4.830725, 4.833347, 4.839246, 
    4.847798, 4.858232, 4.869702, 4.881335, 4.892307, 4.901924, 4.909692, 
    4.91538, 0, 4.999225, 5.004516, 5.011139, 5.018236, 5.025145, 5.026101, 
    5.027013, 5.026284, 5.024335, 5.02012, 5.012819, 5.001411, 4.985559, 
    4.964156, 4.939056, 4.904996, 4.869781, 4.835892, 4.805812, 4.781667, 
    4.764914, 4.756218, 4.755496, 4.762076, 4.774881, 4.792583, 4.813718, 
    4.836743, 4.86009, 4.882205, 4.90162, 4.917064, 4.927612, 4.93287,
  // momentumX(16,30, 0-49)
    4.862476, 4.849107, 4.839384, 4.833349, 4.830894, 4.831782, 4.835658, 
    4.842111, 4.850717, 4.861089, 4.872904, 4.885905, 4.899866, 4.914509, 
    4.92938, 4.966947, 4.978901, 4.992922, 5.007429, 5.020907, 5.032383, 
    5.037577, 5.040587, 5.040208, 5.037008, 5.03027, 5.019615, 5.004519, 
    4.98509, 4.960538, 4.932539, 4.897691, 4.862357, 4.828973, 4.799906, 
    4.777106, 4.761838, 4.754601, 4.75519, 4.762854, 4.776481, 4.794729, 
    4.81613, 4.839152, 4.862225, 4.883802, 4.902434, 4.91689, 4.926324, 
    4.930448,
  // momentumX(16,31, 0-49)
    4.866781, 4.853611, 4.844128, 4.83839, 4.836299, 4.837609, 4.84195, 
    4.848881, 4.857934, 4.868675, 4.880737, 4.893844, 4.9078, 4.922468, 
    4.937697, 4.967824, 4.977847, 4.991458, 5.004806, 5.016727, 5.02653, 
    5.031267, 5.033574, 5.032618, 5.028995, 5.021968, 5.011114, 4.995862, 
    4.976276, 4.951561, 4.923069, 4.889333, 4.855425, 4.823767, 4.796635, 
    4.775844, 4.762507, 4.756995, 4.759011, 4.767756, 4.782095, 4.800686, 
    4.822061, 4.844687, 4.867003, 4.887477, 4.904691, 4.917486, 4.925124, 
    4.927476,
  // momentumX(16,32, 0-49)
    4.871303, 4.858335, 4.849073, 4.843582, 4.841766, 4.843366, 4.848002, 
    4.855215, 4.864517, 4.875458, 4.887661, 4.900854, 4.91489, 4.929732, 
    4.945438, 4.968321, 4.976445, 4.989829, 5.002178, 5.012691, 5.02094, 
    5.025236, 5.026824, 5.025161, 5.020825, 5.013091, 5.001563, 4.985727, 
    4.965698, 4.940761, 4.912001, 4.879725, 4.847709, 4.81828, 4.793566, 
    4.775197, 4.764112, 4.760547, 4.764117, 4.773983, 4.788996, 4.807811, 
    4.82897, 4.850946, 4.872193, 4.891208, 4.906636, 4.917415, 4.922964, 
    4.92335,
  // momentumX(16,33, 0-49)
    4.875925, 4.863193, 4.854173, 4.84893, 4.847354, 4.84918, 4.854009, 
    4.861369, 4.870765, 4.881741, 4.893917, 4.907042, 4.921004, 4.935845, 
    4.951768, 4.968263, 4.974986, 4.988035, 4.999339, 5.008449, 5.015163, 
    5.01895, 5.019767, 5.017297, 5.012066, 5.003394, 4.99095, 4.974339, 
    4.95378, 4.928711, 4.900013, 4.869541, 4.839824, 4.813044, 4.791133, 
    4.775503, 4.766909, 4.765444, 4.770644, 4.78163, 4.797239, 4.816132, 
    4.836852, 4.857888, 4.877718, 4.894889, 4.908136, 4.916543, 4.919724, 
    4.917984,
  // momentumX(16,34, 0-49)
    4.880545, 4.868095, 4.859358, 4.854384, 4.85305, 4.855068, 4.860024, 
    4.867435, 4.876794, 4.887642, 4.899608, 4.912449, 4.926073, 4.940565, 
    4.956202, 4.967526, 4.973517, 4.985917, 4.996002, 5.003626, 5.008771, 
    5.011938, 5.011914, 5.00858, 5.002374, 4.992685, 4.979272, 4.961896, 
    4.940898, 4.915932, 4.887727, 4.859404, 4.832354, 4.80857, 4.789754, 
    4.777088, 4.771133, 4.771847, 4.778687, 4.790736, 4.806821, 4.825599, 
    4.845624, 4.865399, 4.883441, 4.89837, 4.909048, 4.914743, 4.915324, 
    4.911375,
  // momentumX(16,35, 0-49)
    4.885081, 4.87296, 4.864542, 4.85986, 4.858766, 4.86095, 4.865981, 
    4.873355, 4.882562, 4.893137, 4.904713, 4.917045, 4.930042, 4.943787, 
    4.95856, 4.96601, 4.971895, 4.98324, 4.991876, 4.997907, 5.001445, 
    5.003863, 5.002946, 4.998738, 4.991569, 4.980916, 4.966636, 4.948666, 
    4.927465, 4.902946, 4.87573, 4.849896, 4.825834, 4.805314, 4.78979, 
    4.780211, 4.776949, 4.779835, 4.788252, 4.801247, 4.817632, 4.836062, 
    4.855099, 4.87327, 4.889144, 4.901443, 4.909194, 4.911911, 4.909752, 
    4.903614,
  // momentumX(16,36, 0-49)
    4.889462, 4.877706, 4.869629, 4.86524, 4.864367, 4.866679, 4.871722, 
    4.878978, 4.887927, 4.898099, 4.909123, 4.920747, 4.932858, 4.9455, 
    4.958887, 4.963627, 4.969875, 4.979753, 4.986724, 4.99107, 4.992982, 
    4.994537, 4.992704, 4.987673, 4.979637, 4.968187, 4.95327, 4.935, 
    4.913944, 4.890288, 4.86458, 4.841549, 4.820729, 4.803648, 4.791512, 
    4.78504, 4.784429, 4.789392, 4.799244, 4.812998, 4.82945, 4.847256, 
    4.864984, 4.881196, 4.894536, 4.903861, 4.908413, 4.907989, 4.90308, 
    4.894912,
  // momentumX(16,37, 0-49)
    4.893633, 4.882252, 4.874506, 4.870379, 4.869679, 4.872052, 4.877029, 
    4.88408, 4.892673, 4.902333, 4.912676, 4.923434, 4.934464, 4.94574, 
    4.957366, 4.960308, 4.967186, 4.975255, 4.980393, 4.983005, 4.983312, 
    4.983918, 4.981193, 4.975446, 4.966719, 4.954725, 4.939501, 4.921314, 
    4.900814, 4.878473, 4.854766, 4.834799, 4.817393, 4.803834, 4.79508, 
    4.791636, 4.793539, 4.800397, 4.811465, 4.825723, 4.841955, 4.858814, 
    4.87489, 4.888796, 4.899277, 4.905368, 4.906568, 4.902996, 4.895502, 
    4.885627,
  // momentumX(16,38, 0-49)
    4.897552, 4.886523, 4.879058, 4.875122, 4.874506, 4.876844, 4.881657, 
    4.888404, 4.896548, 4.905604, 4.915175, 4.924968, 4.934794, 4.944555, 
    4.954224, 4.956, 4.963574, 4.969604, 4.972828, 4.973719, 4.972487, 
    4.972108, 4.968562, 4.962262, 4.953082, 4.940866, 4.925722, 4.908052, 
    4.888546, 4.867952, 4.846678, 4.82996, 4.816054, 4.805999, 4.800521, 
    4.799932, 4.804125, 4.812616, 4.824606, 4.83905, 4.854722, 4.870285, 
    4.884364, 4.895648, 4.903024, 4.905744, 4.903603, 4.897072, 4.887355, 
    4.876265,
  // momentumX(16,39, 0-49)
    4.901218, 4.89047, 4.88319, 4.879328, 4.878665, 4.880836, 4.885359, 
    4.891698, 4.899304, 4.907685, 4.916423, 4.925197, 4.933774, 4.94198, 
    4.94967, 4.950666, 4.958837, 4.962734, 4.964062, 4.96331, 4.960653, 
    4.959311, 4.955066, 4.948422, 4.939073, 4.926993, 4.912344, 4.89563, 
    4.877538, 4.859074, 4.840569, 4.827199, 4.81678, 4.810116, 4.807721, 
    4.809731, 4.815915, 4.825707, 4.838266, 4.852526, 4.867264, 4.881167, 
    4.892925, 4.901339, 4.905478, 4.904854, 4.89959, 4.890512, 4.879136, 
    4.86748,
  // momentumX(16,40, 0-49)
    4.904684, 4.894101, 4.886861, 4.882905, 4.882024, 4.883858, 4.887946, 
    4.893749, 4.900727, 4.90837, 4.916239, 4.923985, 4.931323, 4.938021, 
    4.943837, 4.94427, 4.952819, 4.954637, 4.954183, 4.951932, 4.948014, 
    4.94579, 4.941018, 4.934273, 4.925064, 4.913489, 4.89974, 4.884389, 
    4.868077, 4.852043, 4.83653, 4.826512, 4.819475, 4.816006, 4.816424, 
    4.820711, 4.828525, 4.839235, 4.851963, 4.865639, 4.879057, 4.89096, 
    4.900132, 4.905531, 4.906458, 4.902721, 4.89478, 4.883789, 4.871507, 
    4.860053,
  // momentumX(16,41, 0-49)
    4.908092, 4.897519, 4.89013, 4.885876, 4.884562, 4.88586, 4.889328, 
    4.894451, 4.90069, 4.907524, 4.914495, 4.921216, 4.927366, 4.932658, 
    4.93679, 4.93676, 4.945415, 4.945338, 4.943303, 4.939752, 4.934779, 
    4.93182, 4.926731, 4.920149, 4.911396, 4.900678, 4.888195, 4.874551, 
    4.86031, 4.846904, 4.834485, 4.827735, 4.823891, 4.823347, 4.826247, 
    4.832436, 4.841479, 4.852689, 4.86517, 4.87786, 4.889602, 4.899222, 
    4.905647, 4.908044, 4.905981, 4.899584, 4.889641, 4.877569, 4.865269, 
    4.854838,
  // momentumX(16,42, 0-49)
    4.911717, 4.900965, 4.893209, 4.888418, 4.886428, 4.886953, 4.889586, 
    4.893843, 4.899196, 4.905123, 4.911144, 4.91684, 4.921854, 4.925863, 
    4.928534, 4.928086, 4.936563, 4.934877, 4.931522, 4.926918, 4.92114, 
    4.917643, 4.912477, 4.906325, 4.89833, 4.888782, 4.877871, 4.866199, 
    4.854226, 4.843546, 4.834213, 4.830557, 4.829648, 4.831701, 4.836706, 
    4.84439, 4.854242, 4.865532, 4.877361, 4.888703, 4.898479, 4.905645, 
    4.909317, 4.908913, 4.904303, 4.895933, 4.88486, 4.872675, 4.861303, 
    4.852696,
  // momentumX(16,43, 0-49)
    4.915979, 4.904849, 4.896491, 4.890907, 4.887977, 4.887463, 4.889009, 
    4.892169, 4.896441, 4.901309, 4.90628, 4.910909, 4.914815, 4.91765, 
    4.919073, 4.918221, 4.926271, 4.923316, 4.918942, 4.91356, 4.907251, 
    4.903452, 4.898461, 4.892997, 4.886028, 4.877912, 4.868806, 4.859283, 
    4.849682, 4.841722, 4.835365, 4.834563, 4.836274, 4.840557, 4.847266, 
    4.856031, 4.866275, 4.877251, 4.888074, 4.897788, 4.905428, 4.910126, 
    4.911233, 4.908454, 4.901965, 4.892494, 4.881298, 4.870026, 4.860497, 
    4.854419,
  // momentumX(16,44, 0-49)
    4.921442, 4.909743, 4.900558, 4.893926, 4.889781, 4.887942, 4.888114, 
    4.889902, 4.892839, 4.89643, 4.900186, 4.903648, 4.906418, 4.90814, 
    4.908477, 4.907215, 4.914638, 4.910761, 4.905677, 4.899805, 4.89325, 
    4.8894, 4.884832, 4.880281, 4.874562, 4.868074, 4.860928, 4.853642, 
    4.846432, 4.841105, 4.837529, 4.839285, 4.843264, 4.849389, 4.857398, 
    4.866843, 4.877102, 4.887429, 4.896988, 4.90492, 4.910418, 4.912833, 
    4.911785, 4.907272, 4.89976, 4.890192, 4.879921, 4.87054, 4.863652, 
    4.860648,
  // momentumX(16,45, 0-49)
    4.928774, 4.916354, 4.906143, 4.89823, 4.892606, 4.889152, 4.887639, 
    4.887737, 4.889032, 4.891066, 4.893369, 4.895489, 4.897025, 4.897626, 
    4.89697, 4.895264, 4.901911, 4.897421, 4.891912, 4.885824, 4.879295, 
    4.875637, 4.871709, 4.868249, 4.863946, 4.85921, 4.854095, 4.849058, 
    4.844183, 4.84133, 4.840287, 4.844272, 4.850154, 4.857734, 4.866662, 
    4.876428, 4.886393, 4.895836, 4.903998, 4.910158, 4.913705, 4.914233, 
    4.911644, 4.906223, 4.898661, 4.890035, 4.881682, 4.875031, 4.871395, 
    4.871812,
  // momentumX(16,46, 0-49)
    4.93868, 4.925437, 4.914054, 4.904667, 4.897326, 4.891982, 4.888477, 
    4.886553, 4.885867, 4.886013, 4.886566, 4.887105, 4.88724, 4.886635, 
    4.884993, 4.88277, 4.888525, 4.883657, 4.877955, 4.871884, 4.865617, 
    4.862357, 4.859235, 4.856978, 4.854181, 4.851244, 4.848159, 4.845309, 
    4.842661, 4.842082, 4.843284, 4.849162, 4.856587, 4.865265, 4.874779, 
    4.88458, 4.894042, 4.902493, 4.909286, 4.913868, 4.915846, 4.915076, 
    4.911729, 4.906325, 4.899712, 4.892994, 4.887399, 4.884111, 4.884117, 
    4.888099,
  // momentumX(16,47, 0-49)
    4.951799, 4.937706, 4.925067, 4.914071, 4.904827, 4.897355, 4.891575, 
    4.887312, 4.884302, 4.88222, 4.880702, 4.879376, 4.87789, 4.875928, 
    4.873226, 4.870365, 4.875134, 4.870023, 4.864284, 4.858397, 4.852556, 
    4.849838, 4.847615, 4.846592, 4.845309, 4.844142, 4.843019, 4.842241, 
    4.841671, 4.843141, 4.846299, 4.853746, 4.862389, 4.871863, 4.881702, 
    4.891355, 4.900224, 4.907723, 4.913341, 4.916712, 4.917672, 4.916331, 
    4.913086, 4.908631, 4.903881, 4.899878, 4.897662, 4.89813, 4.901938, 
    4.909441,
  // momentumX(16,48, 0-49)
    4.968619, 4.953721, 4.939814, 4.927141, 4.915872, 4.906098, 4.897817, 
    4.890945, 4.885314, 4.880691, 4.876794, 4.873322, 4.869973, 4.866468, 
    4.862566, 4.858901, 4.862593, 4.857264, 4.85155, 4.845926, 4.840598, 
    4.838478, 4.837162, 4.837315, 4.837472, 4.837968, 4.838675, 4.839813, 
    4.841158, 4.844455, 4.849295, 4.858031, 4.867624, 4.877662, 4.887666, 
    4.897097, 4.905418, 4.912148, 4.916932, 4.919597, 4.920197, 4.91906, 
    4.916761, 4.914085, 4.911936, 4.911226, 4.912759, 4.917141, 4.92471, 
    4.935537,
  // momentumX(16,49, 0-49)
    4.997341, 4.981748, 4.96641, 4.95162, 4.937616, 4.924573, 4.9126, 
    4.901742, 4.89198, 4.883229, 4.875348, 4.868152, 4.861418, 4.854907, 
    4.848384, 4.843278, 4.852906, 4.845834, 4.83861, 4.832042, 4.8264, 
    4.827126, 4.82929, 4.833854, 4.837558, 4.840845, 4.843235, 4.844953, 
    4.845376, 4.847987, 4.852074, 4.862319, 4.872993, 4.88364, 4.893794, 
    4.902972, 4.910752, 4.916822, 4.921046, 4.923507, 4.924527, 4.92465, 
    4.9246, 4.925184, 4.927189, 4.931278, 4.93792, 4.947337, 4.959503, 
    4.974175,
  // momentumX(17,0, 0-49)
    4.932086, 4.910845, 4.892358, 4.876889, 4.864563, 4.855368, 4.849143, 
    4.845583, 4.844279, 4.84473, 4.846404, 4.84877, 4.851345, 4.853716, 
    4.855547, 4.85666, 4.858193, 4.857396, 4.855773, 4.853347, 4.850139, 
    4.846555, 4.84232, 4.837674, 4.832701, 4.827689, 4.822936, 4.818818, 
    4.815685, 4.813998, 4.813952, 4.81605, 4.819995, 4.825649, 4.832704, 
    4.840699, 4.849057, 4.857137, 4.864295, 4.869975, 4.873768, 4.8755, 
    4.875279, 4.87353, 4.870981, 4.868604, 4.867512, 4.868828, 4.873548, 
    4.882422,
  // momentumX(17,1, 0-49)
    4.927293, 4.906449, 4.888511, 4.873724, 4.862199, 4.853904, 4.848652, 
    4.846119, 4.845862, 4.847353, 4.850029, 4.853331, 4.856744, 4.859819, 
    4.862175, 4.863629, 4.866576, 4.865678, 4.863865, 4.861151, 4.857523, 
    4.853695, 4.849001, 4.843752, 4.837935, 4.831862, 4.825829, 4.820256, 
    4.815511, 4.812222, 4.810579, 4.811505, 4.814435, 4.819283, 4.825787, 
    4.83351, 4.841879, 4.850229, 4.85787, 4.864164, 4.868599, 4.870879, 
    4.870985, 4.869229, 4.866257, 4.863015, 4.860652, 4.860381, 4.863338, 
    4.87043,
  // momentumX(17,2, 0-49)
    4.925047, 4.904743, 4.887443, 4.873371, 4.862625, 4.855145, 4.85073, 
    4.849032, 4.849593, 4.851871, 4.855292, 4.859291, 4.863336, 4.866961, 
    4.86975, 4.871462, 4.875763, 4.874875, 4.873009, 4.870171, 4.866305, 
    4.862421, 4.857438, 4.851728, 4.845177, 4.838098, 4.830777, 4.823665, 
    4.817146, 4.812004, 4.80843, 4.807797, 4.809296, 4.812929, 4.81851, 
    4.825661, 4.833847, 4.842411, 4.850638, 4.857832, 4.863382, 4.866856, 
    4.868075, 4.867185, 4.864679, 4.861393, 4.858432, 4.857043, 4.85846, 
    4.863751,
  // momentumX(17,3, 0-49)
    4.924704, 4.905055, 4.888456, 4.875116, 4.865107, 4.858351, 4.854629, 
    4.85358, 4.85474, 4.85757, 4.861506, 4.865989, 4.870497, 4.874556, 
    4.877724, 4.879621, 4.88518, 4.884454, 4.882708, 4.879936, 4.876042, 
    4.872316, 4.867249, 4.861258, 4.854124, 4.846151, 4.837596, 4.828926, 
    4.820539, 4.813347, 4.807551, 4.805, 4.804668, 4.806671, 4.810932, 
    4.817171, 4.824917, 4.833555, 4.842372, 4.850632, 4.85764, 4.862832, 
    4.865854, 4.866643, 4.865483, 4.863023, 4.860238, 4.858329, 4.858582, 
    4.862187,
  // momentumX(17,4, 0-49)
    4.925554, 4.906652, 4.890803, 4.878195, 4.868879, 4.862763, 4.859605, 
    4.859044, 4.860619, 4.863809, 4.868073, 4.87288, 4.877728, 4.882148, 
    4.885689, 4.887709, 4.894379, 4.894003, 4.892564, 4.890065, 4.886366, 
    4.88302, 4.878093, 4.872019, 4.8645, 4.855797, 4.846127, 4.835956, 
    4.825689, 4.816328, 4.808094, 4.803315, 4.800786, 4.800761, 4.803308, 
    4.808267, 4.815266, 4.823757, 4.833058, 4.842415, 4.85107, 4.858335, 
    4.863684, 4.866829, 4.867804, 4.867007, 4.865207, 4.863475, 4.863067, 
    4.865251,
  // momentumX(17,5, 0-49)
    4.926895, 4.908814, 4.893754, 4.881882, 4.873228, 4.86768, 4.86499, 
    4.864796, 4.866652, 4.870066, 4.874532, 4.879558, 4.884674, 4.889433, 
    4.893384, 4.89547, 4.903042, 4.903224, 4.902287, 4.900254, 4.896966, 
    4.894212, 4.889642, 4.883701, 4.87602, 4.866802, 4.856206, 4.844675, 
    4.832611, 4.821059, 4.810258, 4.803021, 4.79799, 4.795586, 4.796041, 
    4.799346, 4.805257, 4.813318, 4.822897, 4.833249, 4.843571, 4.853073, 
    4.861067, 4.867047, 4.870778, 4.872372, 4.872322, 4.871489, 4.871013, 
    4.872166,
  // momentumX(17,6, 0-49)
    4.928093, 4.910898, 4.896666, 4.885541, 4.877535, 4.872518, 4.870237, 
    4.870338, 4.872396, 4.875957, 4.880558, 4.885754, 4.891115, 4.89623, 
    4.900664, 4.902766, 4.910966, 4.911911, 4.911652, 4.910261, 4.907574, 
    4.905591, 4.901582, 4.895983, 4.888383, 4.878903, 4.867634, 4.85497, 
    4.841294, 4.827643, 4.814258, 4.804423, 4.796666, 4.791592, 4.789618, 
    4.790914, 4.795382, 4.802684, 4.812258, 4.823384, 4.835237, 4.84695, 
    4.857692, 4.866757, 4.873649, 4.878177, 4.88052, 4.881258, 4.881336, 
    4.881945,
  // momentumX(17,7, 0-49)
    4.928635, 4.912382, 4.89902, 4.888669, 4.88132, 4.87683, 4.874942, 
    4.875315, 4.877554, 4.88124, 4.88596, 4.891318, 4.896939, 4.902454, 
    4.907468, 4.909537, 4.918041, 4.919922, 4.920493, 4.919884, 4.91795, 
    4.916876, 4.913595, 4.908529, 4.901253, 4.891789, 4.880151, 4.866659, 
    4.851659, 4.836112, 4.820251, 4.80779, 4.797184, 4.789228, 4.78455, 
    4.783514, 4.786196, 4.792386, 4.801616, 4.813207, 4.826326, 4.840052, 
    4.853444, 4.865614, 4.875832, 4.883608, 4.8888, 4.891662, 4.892874, 
    4.893465,
  // momentumX(17,8, 0-49)
    4.928143, 4.912886, 4.900441, 4.890904, 4.884245, 4.880311, 4.878841, 
    4.87951, 4.88195, 4.885783, 4.890644, 4.89619, 4.902103, 4.908071, 
    4.913764, 4.915773, 4.92422, 4.927168, 4.928677, 4.928949, 4.927879, 
    4.927794, 4.925365, 4.920992, 4.914267, 4.905104, 4.893435, 4.879482, 
    4.863534, 4.846408, 4.828302, 4.813304, 4.799834, 4.788882, 4.781299, 
    4.777662, 4.778239, 4.782969, 4.791487, 4.803172, 4.817198, 4.83261, 
    4.848373, 4.863461, 4.876935, 4.88804, 4.896313, 4.901678, 4.904503, 
    4.905589,
  // momentumX(17,9, 0-49)
    4.926387, 4.91217, 4.900692, 4.892024, 4.88611, 4.882786, 4.881791, 
    4.882813, 4.88551, 4.889541, 4.894586, 4.900361, 4.906602, 4.913068, 
    4.919524, 4.921489, 4.929521, 4.933596, 4.936105, 4.937315, 4.937177, 
    4.938101, 4.936598, 4.933035, 4.927056, 4.918464, 4.90711, 4.893102, 
    4.876647, 4.85835, 4.838352, 4.821018, 4.804783, 4.790828, 4.780226, 
    4.773788, 4.771987, 4.774931, 4.782368, 4.793742, 4.808257, 4.824928, 
    4.84266, 4.860311, 4.876772, 4.891061, 4.902427, 4.910475, 4.915247, 
    4.917273,
  // momentumX(17,10, 0-49)
    4.923273, 4.910128, 4.899665, 4.891922, 4.886822, 4.884184, 4.883743, 
    4.885196, 4.888224, 4.892519, 4.897807, 4.903848, 4.910443, 4.917434, 
    4.924696, 4.92671, 4.934017, 4.939202, 4.942721, 4.944888, 4.945706, 
    4.947608, 4.947049, 4.944363, 4.939278, 4.931495, 4.920787, 4.907132, 
    4.890639, 4.871647, 4.850207, 4.83084, 4.812048, 4.795187, 4.781552, 
    4.772192, 4.767801, 4.768667, 4.774671, 4.785334, 4.799887, 4.817338, 
    4.836549, 4.856289, 4.875316, 4.892464, 4.906739, 4.917458, 4.924351, 
    4.92766,
  // momentumX(17,11, 0-49)
    4.918819, 4.906762, 4.897353, 4.890594, 4.886381, 4.884509, 4.884711, 
    4.886684, 4.890129, 4.89476, 4.90034, 4.906679, 4.913639, 4.921144, 
    4.929193, 4.931473, 4.937835, 4.944029, 4.948521, 4.951626, 4.953395, 
    4.95619, 4.956545, 4.954758, 4.950663, 4.943872, 4.934094, 4.921172, 
    4.905105, 4.885919, 4.863553, 4.842531, 4.821484, 4.801915, 4.785327, 
    4.773007, 4.765884, 4.764438, 4.768693, 4.778259, 4.792406, 4.810146, 
    4.830305, 4.851591, 4.872667, 4.89222, 4.909069, 4.922284, 4.931321, 
    4.936136,
  // momentumX(17,12, 0-49)
    4.913151, 4.902174, 4.89384, 4.888111, 4.884847, 4.883822, 4.884756, 
    4.887339, 4.891278, 4.896312, 4.90223, 4.908882, 4.91619, 4.924158, 
    4.932895, 4.935816, 4.941145, 4.948177, 4.953555, 4.957557, 4.960253, 
    4.96382, 4.965019, 4.964102, 4.961035, 4.955356, 4.946728, 4.934856, 
    4.919626, 4.900735, 4.877989, 4.855725, 4.832791, 4.810797, 4.791426, 
    4.776199, 4.766277, 4.762349, 4.764593, 4.772719, 4.786045, 4.803592, 
    4.82417, 4.846443, 4.869005, 4.890441, 4.90943, 4.924849, 4.935921, 
    4.942349,
  // momentumX(17,13, 0-49)
    4.906466, 4.896542, 4.889278, 4.884605, 4.882339, 4.882226, 4.883963, 
    4.887234, 4.891738, 4.897228, 4.903514, 4.91048, 4.918095, 4.926425, 
    4.93566, 4.939777, 4.944144, 4.951789, 4.95794, 4.962779, 4.966364, 
    4.970561, 4.972504, 4.972393, 4.970335, 4.96582, 4.958477, 4.947888, 
    4.933827, 4.915659, 4.893061, 4.869974, 4.845552, 4.821473, 4.799566, 
    4.781562, 4.768855, 4.762346, 4.762383, 4.768782, 4.78092, 4.797838, 
    4.818337, 4.841057, 4.864547, 4.887329, 4.907979, 4.925239, 4.938151, 
    4.946199,
  // momentumX(17,14, 0-49)
    4.899024, 4.89009, 4.883871, 4.880249, 4.879004, 4.879846, 4.882438, 
    4.886447, 4.891568, 4.897552, 4.90422, 4.911483, 4.919337, 4.927886, 
    4.937351, 4.943377, 4.947018, 4.955034, 4.961828, 4.967443, 4.971882, 
    4.976558, 4.979132, 4.979733, 4.97862, 4.975255, 4.969245, 4.960069, 
    4.947399, 4.930287, 4.908312, 4.884778, 4.859268, 4.833473, 4.809331, 
    4.788751, 4.773347, 4.764234, 4.761935, 4.766388, 4.777039, 4.792955, 
    4.812939, 4.835619, 4.859524, 4.883137, 4.904978, 4.923697, 4.9382, 
    4.947796,
  // momentumX(17,15, 0-49)
    4.891112, 4.883087, 4.877852, 4.875248, 4.875012, 4.876813, 4.880279, 
    4.885053, 4.890813, 4.897305, 4.904356, 4.911882, 4.919893, 4.928493, 
    4.93788, 4.946609, 4.949912, 4.958069, 4.965397, 4.97174, 4.97701, 
    4.982026, 4.985116, 4.986323, 4.986053, 4.983757, 4.979042, 4.971297, 
    4.960118, 4.944283, 4.923313, 4.899639, 4.873401, 4.84626, 4.820212, 
    4.797309, 4.779364, 4.767699, 4.763014, 4.76538, 4.774317, 4.788934, 
    4.808044, 4.830278, 4.854156, 4.87815, 4.900752, 4.920557, 4.936386, 
    4.947409,
  // momentumX(17,16, 0-49)
    4.883029, 4.875806, 4.871468, 4.869812, 4.870532, 4.873254, 4.877571, 
    4.883094, 4.889482, 4.896476, 4.903892, 4.911646, 4.919736, 4.928235, 
    4.937255, 4.949426, 4.952873, 4.96102, 4.968817, 4.975876, 4.981983, 
    4.987225, 4.990734, 4.992444, 4.992887, 4.991526, 4.987975, 4.981569, 
    4.971848, 4.957378, 4.937684, 4.914083, 4.887414, 4.859268, 4.831649, 
    4.806712, 4.786437, 4.772339, 4.765296, 4.765512, 4.772596, 4.785703, 
    4.803671, 4.825141, 4.84864, 4.872643, 4.89564, 4.916207, 4.933103, 
    4.945402,
  // momentumX(17,17, 0-49)
    4.875055, 4.868514, 4.864955, 4.864135, 4.86571, 4.869261, 4.87435, 
    4.880558, 4.88753, 4.89499, 4.902754, 4.910722, 4.918859, 4.927171, 
    4.935653, 4.951737, 4.955822, 4.963933, 4.972224, 4.980051, 4.987048, 
    4.992446, 4.996313, 4.998434, 4.999444, 4.99883, 4.99623, 4.990953, 
    4.982525, 4.969369, 4.951089, 4.927674, 4.900793, 4.871935, 4.843071, 
    4.816412, 4.794065, 4.777717, 4.768412, 4.766494, 4.771667, 4.783143, 
    4.799794, 4.820279, 4.843141, 4.866875, 4.889984, 4.911039, 4.928771, 
    4.942188,
  // momentumX(17,18, 0-49)
    4.867438, 4.861432, 4.858498, 4.858359, 4.860627, 4.864854, 4.870573, 
    4.87735, 4.884819, 4.892704, 4.900818, 4.909043, 4.917301, 4.925497, 
    4.93346, 4.953443, 4.958536, 4.966762, 4.975693, 4.984436, 4.992451, 
    4.997995, 5.002215, 5.004687, 5.006111, 5.006001, 5.004041, 4.999564, 
    4.992125, 4.980086, 4.963223, 4.940009, 4.913056, 4.88373, 4.853928, 
    4.825867, 4.801744, 4.783382, 4.771981, 4.768018, 4.771304, 4.781112, 
    4.796357, 4.815728, 4.83779, 4.861065, 4.884079, 4.905415, 4.923792, 
    4.938173,
  // momentumX(17,19, 0-49)
    4.860362, 4.854715, 4.852209, 4.85253, 4.855262, 4.859932, 4.866065, 
    4.87323, 4.881079, 4.889356, 4.89789, 4.906549, 4.915184, 4.923564, 
    4.931289, 4.954461, 4.960647, 4.969331, 4.979218, 4.989158, 4.998429, 
    5.004205, 5.008854, 5.011667, 5.013352, 5.01345, 5.011711, 5.007554, 
    5.000636, 4.989366, 4.973771, 4.950686, 4.92374, 4.894152, 4.863704, 
    4.834578, 4.809007, 4.788918, 4.775646, 4.769795, 4.771284, 4.77946, 
    4.793291, 4.811497, 4.83268, 4.855388, 4.878173, 4.899641, 4.918513, 
    4.933718,
  // momentumX(17,20, 0-49)
    4.854655, 4.849918, 4.84861, 4.850455, 4.855026, 4.861779, 4.870096, 
    4.879328, 4.888843, 4.898059, 4.906477, 4.913717, 4.919533, 4.923843, 
    4.926725, 0, 4.976701, 4.980468, 4.985542, 4.99134, 4.997496, 5.000072, 
    5.003079, 5.005518, 5.008004, 5.009818, 5.010391, 5.008807, 5.004483, 
    4.995662, 4.982596, 4.960472, 4.934066, 4.904542, 4.873656, 4.843603, 
    4.816685, 4.794946, 4.779853, 4.772143, 4.771838, 4.778371, 4.790754, 
    4.807751, 4.827991, 4.850053, 4.872515, 4.894001, 4.913239, 4.929135,
  // momentumX(17,21, 0-49)
    4.849359, 4.844958, 4.844018, 4.846222, 4.851108, 4.858102, 4.866564, 
    4.875849, 4.885345, 4.89451, 4.90289, 4.910137, 4.916014, 4.920402, 
    4.923314, 0, 4.978804, 4.983113, 4.98882, 4.995245, 5.001908, 5.003341, 
    5.005481, 5.007151, 5.009163, 5.010862, 5.011708, 5.010763, 5.007414, 
    4.999859, 4.988595, 4.967202, 4.941577, 4.912706, 4.882171, 4.852049, 
    4.824604, 4.801916, 4.785548, 4.776368, 4.774518, 4.77953, 4.790494, 
    4.806223, 4.825388, 4.846598, 4.868461, 4.889622, 4.908823, 4.924966,
  // momentumX(17,22, 0-49)
    4.84491, 4.840719, 4.840024, 4.842488, 4.847629, 4.854852, 4.863504, 
    4.872935, 4.882536, 4.891777, 4.900223, 4.907533, 4.913461, 4.917856, 
    4.920673, 0, 4.980448, 4.985187, 4.991485, 4.998569, 5.005846, 5.006361, 
    5.007894, 5.009054, 5.010793, 5.012468, 5.013533, 5.01302, 5.010294, 
    5.003533, 4.9935, 4.972336, 4.947056, 4.918531, 4.888209, 4.858057, 
    4.830273, 4.806931, 4.789643, 4.779356, 4.776308, 4.780115, 4.789931, 
    4.804622, 4.822892, 4.843383, 4.864727, 4.885594, 4.904738, 4.921063,
  // momentumX(17,23, 0-49)
    4.841343, 4.837268, 4.836722, 4.839362, 4.844692, 4.852111, 4.860959, 
    4.870574, 4.880348, 4.889748, 4.898341, 4.905778, 4.911798, 4.916217, 
    4.918941, 0, 4.982242, 4.987259, 4.993968, 5.001531, 5.009266, 5.00898, 
    5.009981, 5.010692, 5.012161, 5.013753, 5.014909, 5.014637, 5.012286, 
    5.006017, 4.996813, 4.975653, 4.950515, 4.922195, 4.892049, 4.861947, 
    4.834018, 4.810307, 4.792441, 4.781416, 4.77753, 4.780464, 4.789426, 
    4.803322, 4.820889, 4.840794, 4.86169, 4.882262, 4.901279, 4.917653,
  // momentumX(17,24, 0-49)
    4.838642, 4.834622, 4.834155, 4.836901, 4.842365, 4.849943, 4.858972, 
    4.868788, 4.878774, 4.888392, 4.897195, 4.904826, 4.911006, 4.915524, 
    4.918251, 0, 4.984415, 4.98959, 4.996536, 5.004384, 5.012406, 5.011586, 
    5.012234, 5.012639, 5.013902, 5.015387, 5.016535, 5.016338, 5.014139, 
    5.008089, 4.999325, 4.978053, 4.952898, 4.924624, 4.894527, 4.864416, 
    4.836373, 4.812413, 4.794162, 4.782639, 4.778178, 4.7805, 4.788852, 
    4.80217, 4.819218, 4.838678, 4.859221, 4.879544, 4.898427, 4.914783,
  // momentumX(17,25, 0-49)
    4.836769, 4.832759, 4.832325, 4.83513, 4.840688, 4.8484, 4.857604, 
    4.867634, 4.877865, 4.887749, 4.896824, 4.904718, 4.911138, 4.915858, 
    4.918736, 0, 4.986551, 4.991792, 4.998822, 5.006766, 5.014881, 5.013883, 
    5.014416, 5.014708, 5.015873, 5.017272, 5.018345, 5.018085, 5.015834, 
    5.009744, 5.001011, 4.979569, 4.954289, 4.925926, 4.895759, 4.865575, 
    4.83743, 4.813322, 4.794866, 4.783079, 4.778309, 4.780292, 4.788291, 
    4.801262, 4.817979, 4.837139, 4.85742, 4.877531, 4.89625, 4.912501,
  // momentumX(17,26, 0-49)
    4.835672, 4.83165, 4.831218, 4.834058, 4.839693, 4.847535, 4.856926, 
    4.867199, 4.877722, 4.887929, 4.897342, 4.905571, 4.912312, 4.917341, 
    4.920526, 0, 4.988527, 4.993752, 5.000716, 5.008561, 5.016568, 5.015782, 
    5.016457, 5.016857, 5.018059, 5.019417, 5.020375, 5.019933, 5.017445, 
    5.011068, 5.001957, 4.980327, 4.954838, 4.92627, 4.895921, 4.865594, 
    4.837351, 4.813177, 4.794672, 4.782838, 4.778008, 4.779906, 4.787796, 
    4.800632, 4.817194, 4.836185, 4.856286, 4.876206, 4.894732, 4.910787,
  // momentumX(17,27, 0-49)
    4.835305, 4.831254, 4.830816, 4.833688, 4.83941, 4.847407, 4.857031, 
    4.86761, 4.878496, 4.889104, 4.898934, 4.907572, 4.914705, 4.920119, 
    4.923718, 0, 4.990418, 4.995515, 5.002238, 5.00977, 5.01746, 5.017213, 
    5.018252, 5.01895, 5.020303, 5.021653, 5.022446, 5.021699, 5.018786, 
    5.011879, 5.002003, 4.980161, 4.954391, 4.925523, 4.894915, 4.864421, 
    4.836125, 4.812012, 4.793656, 4.782018, 4.777392, 4.779467, 4.787487, 
    4.800394, 4.816962, 4.835893, 4.855869, 4.875599, 4.893869, 4.909608,
  // momentumX(17,28, 0-49)
    4.835628, 4.831538, 4.831094, 4.834014, 4.839862, 4.848079, 4.85802, 
    4.869009, 4.880377, 4.891504, 4.90185, 4.910967, 4.91853, 4.924347, 
    4.928369, 0, 4.992599, 4.997404, 5.003668, 5.010651, 5.017807, 5.018314, 
    5.019859, 5.020988, 5.022568, 5.023917, 5.02448, 5.023301, 5.019778, 
    5.01211, 5.00112, 4.979014, 4.952876, 4.923621, 4.892708, 4.862062, 
    4.833807, 4.809922, 4.791938, 4.780753, 4.776589, 4.779086, 4.787449, 
    4.8006, 4.817302, 4.836254, 4.856133, 4.875648, 4.893589, 4.908889,
  // momentumX(17,29, 0-49)
    4.836607, 4.832465, 4.832018, 4.835017, 4.841056, 4.849597, 4.859998, 
    4.871566, 4.883592, 4.8954, 4.906381, 4.916035, 4.924014, 4.930147, 
    4.934448, 0, 4.994762, 4.999057, 5.004619, 5.010811, 5.01722, 5.01852, 
    5.020604, 5.022212, 5.02405, 5.025388, 5.025658, 5.023925, 5.019612, 
    5.010951, 4.998516, 4.976011, 4.949397, 4.919718, 4.888555, 4.857924, 
    4.829979, 4.806665, 4.789436, 4.779088, 4.77575, 4.778986, 4.787952, 
    4.80154, 4.818505, 4.837532, 4.857296, 4.876508, 4.89396, 4.908601,
  // momentumX(17,30, 0-49)
    4.837832, 4.833149, 4.831962, 4.833973, 4.838768, 4.84586, 4.854743, 
    4.86493, 4.875998, 4.887613, 4.899509, 4.911485, 4.923332, 4.93478, 
    4.945404, 4.975517, 4.979926, 4.9902, 5.001615, 5.01291, 5.023316, 
    5.028723, 5.033325, 5.036073, 5.037669, 5.037555, 5.035443, 5.030748, 
    5.023216, 5.011344, 4.995587, 4.971336, 4.943355, 4.912786, 4.881282, 
    4.850867, 4.823629, 4.801392, 4.785451, 4.776451, 4.77439, 4.778745, 
    4.788615, 4.802867, 4.820241, 4.839418, 4.859073, 4.87792, 4.894762, 
    4.908581,
  // momentumX(17,31, 0-49)
    4.840512, 4.836057, 4.835127, 4.837435, 4.842564, 4.85002, 4.85927, 
    4.869801, 4.881155, 4.892956, 4.904926, 4.916868, 4.928643, 4.940125, 
    4.951134, 4.976396, 4.981072, 4.990958, 5.001443, 5.011515, 5.020609, 
    5.025819, 5.029953, 5.032291, 5.033554, 5.033181, 5.03083, 5.025838, 
    5.017842, 5.005279, 4.988306, 4.964038, 4.936157, 4.905926, 4.875092, 
    4.845701, 4.81979, 4.799075, 4.784719, 4.777233, 4.77651, 4.781954, 
    4.792624, 4.80736, 4.824892, 4.843892, 4.863036, 4.881039, 4.896733, 
    4.90915,
  // momentumX(17,32, 0-49)
    4.84394, 4.839687, 4.838961, 4.84147, 4.8468, 4.854445, 4.863869, 
    4.874544, 4.886004, 4.897867, 4.909857, 4.921802, 4.933619, 4.9453, 
    4.956847, 4.976905, 4.981479, 4.991234, 5.00101, 5.010061, 5.018018, 
    5.023118, 5.026866, 5.028792, 5.02958, 5.028664, 5.025671, 5.019921, 
    5.011018, 4.997434, 4.979104, 4.954812, 4.927166, 4.897542, 4.867736, 
    4.839773, 4.815597, 4.796778, 4.784322, 4.7786, 4.779403, 4.786065, 
    4.797607, 4.812852, 4.830517, 4.849267, 4.867775, 4.88477, 4.899115, 
    4.909908,
  // momentumX(17,33, 0-49)
    4.848188, 4.844136, 4.843581, 4.846228, 4.851653, 4.859349, 4.868777, 
    4.879411, 4.890791, 4.902544, 4.914413, 4.926251, 4.938032, 4.949833, 
    4.961806, 4.976944, 4.981427, 4.991122, 5.000261, 5.008378, 5.015282, 
    5.02028, 5.023657, 5.025142, 5.025333, 5.023657, 5.019734, 5.012911, 
    5.002809, 4.988014, 4.968327, 4.944061, 4.916827, 4.88808, 4.859641, 
    4.83347, 4.811376, 4.794761, 4.784458, 4.780696, 4.783165, 4.791138, 
    4.803601, 4.819355, 4.837107, 4.855516, 4.87325, 4.889057, 4.901842, 
    4.910791,
  // momentumX(17,34, 0-49)
    4.853289, 4.849438, 4.849027, 4.851749, 4.857172, 4.864788, 4.874062, 
    4.88448, 4.895594, 4.907053, 4.91862, 4.930174, 4.941731, 4.953428, 
    4.965522, 4.976438, 4.981064, 4.990592, 4.999053, 5.006239, 5.012118, 
    5.01695, 5.019924, 5.020919, 5.020409, 5.017825, 5.01279, 5.004707, 
    4.993249, 4.9772, 4.956297, 4.932189, 4.905595, 4.878024, 4.85128, 
    4.827223, 4.8075, 4.793324, 4.785354, 4.783679, 4.787896, 4.797219, 
    4.810601, 4.826828, 4.844588, 4.862535, 4.879337, 4.893764, 4.904784, 
    4.911689,
  // momentumX(17,35, 0-49)
    4.859222, 4.855562, 4.855252, 4.857974, 4.863289, 4.870693, 4.879658, 
    4.889689, 4.900362, 4.911344, 4.922421, 4.933497, 4.944608, 4.955915, 
    4.967728, 4.975316, 4.980386, 4.989532, 4.997201, 5.003416, 5.00826, 
    5.012824, 5.015333, 5.015789, 5.014503, 5.010921, 5.004682, 4.995273, 
    4.982435, 4.965222, 4.943371, 4.919636, 4.893962, 4.867884, 4.843148, 
    4.82148, 4.804347, 4.792766, 4.787225, 4.787683, 4.793653, 4.804296, 
    4.81854, 4.835147, 4.852794, 4.870125, 4.885816, 4.898671, 4.907736, 
    4.912441,
  // momentumX(17,36, 0-49)
    4.865902, 4.862398, 4.862123, 4.86475, 4.869839, 4.876892, 4.885399, 
    4.894885, 4.904952, 4.915292, 4.925711, 4.936127, 4.946576, 4.957216, 
    4.968345, 4.973502, 4.979285, 4.987776, 4.994511, 4.999691, 5.003481, 
    5.007654, 5.009626, 5.009497, 5.007393, 5.002791, 4.995346, 4.984653, 
    4.97054, 4.952381, 4.929957, 4.90688, 4.882451, 4.858187, 4.835741, 
    4.816682, 4.802279, 4.793364, 4.790259, 4.792812, 4.800456, 4.812315, 
    4.827287, 4.844121, 4.861478, 4.877997, 4.892375, 4.903469, 4.910425, 
    4.912837,
  // momentumX(17,37, 0-49)
    4.873171, 4.869758, 4.869428, 4.871847, 4.876582, 4.883149, 4.891055, 
    4.899855, 4.909174, 4.918733, 4.928355, 4.93796, 4.947573, 4.957314, 
    4.967422, 4.970922, 4.977585, 4.98515, 4.990809, 4.994896, 4.997612, 
    5.001259, 5.002623, 5.001882, 4.998955, 4.993373, 4.984812, 4.972988, 
    4.957819, 4.939039, 4.916505, 4.894428, 4.871589, 4.849447, 4.829532, 
    4.813232, 4.801623, 4.795353, 4.794603, 4.799121, 4.808279, 4.821166, 
    4.836657, 4.853489, 4.870317, 4.885788, 4.898634, 4.907787, 4.91253, 
    4.912643,
  // momentumX(17,38, 0-49)
    4.880799, 4.877385, 4.876884, 4.878968, 4.88322, 4.889169, 4.896352, 
    4.904349, 4.912816, 4.921493, 4.930215, 4.938902, 4.947552, 4.956231, 
    4.965086, 4.967517, 4.975098, 4.981501, 4.985966, 4.988914, 4.990543, 
    4.993541, 4.994239, 4.992883, 4.989176, 4.982718, 4.973215, 4.960507, 
    4.944603, 4.925617, 4.903484, 4.88278, 4.861875, 4.842131, 4.824929, 
    4.811468, 4.802634, 4.798907, 4.800348, 4.806618, 4.817043, 4.830686, 
    4.846407, 4.862938, 4.878937, 4.893082, 4.904164, 4.911223, 4.913716, 
    4.911637,
  // momentumX(17,39, 0-49)
    4.8885, 4.884964, 4.884163, 4.885783, 4.889422, 4.894643, 4.901007, 
    4.908122, 4.915665, 4.923398, 4.931163, 4.938869, 4.946483, 4.95401, 
    4.961489, 4.963247, 4.971654, 4.976719, 4.979917, 4.981703, 4.982242, 
    4.984488, 4.984486, 4.982543, 4.978146, 4.970976, 4.960778, 4.947517, 
    4.931282, 4.912557, 4.891349, 4.872391, 4.853734, 4.836616, 4.822244, 
    4.811627, 4.805473, 4.804114, 4.807503, 4.815238, 4.826606, 4.840658, 
    4.856246, 4.87211, 4.886935, 4.899451, 4.908543, 4.913409, 4.913702, 
    4.909656,
  // momentumX(17,40, 0-49)
    4.895968, 4.892166, 4.890924, 4.891946, 4.894863, 4.899263, 4.90474, 
    4.910928, 4.917522, 4.924296, 4.931087, 4.937795, 4.944351, 4.950702, 
    4.956784, 4.958094, 4.967124, 4.970757, 4.972659, 4.973285, 4.972751, 
    4.974173, 4.973469, 4.971002, 4.966048, 4.958385, 4.947799, 4.934374, 
    4.918255, 4.900277, 4.880496, 4.863629, 4.847486, 4.833153, 4.821659, 
    4.813825, 4.810189, 4.810955, 4.815989, 4.824837, 4.836764, 4.850812, 
    4.865849, 4.880637, 4.893913, 4.904496, 4.911415, 4.914057, 4.912313, 
    4.906664,
  // momentumX(17,41, 0-49)
    4.902921, 4.898695, 4.89686, 4.897158, 4.899249, 4.902759, 4.907311, 
    4.91256, 4.918214, 4.924046, 4.929891, 4.935626, 4.941149, 4.946351, 
    4.951089, 4.952054, 4.96143, 4.963621, 4.964247, 4.963741, 4.962173, 
    4.962739, 4.96137, 4.958476, 4.95314, 4.945245, 4.934614, 4.921438, 
    4.905893, 4.88913, 4.871221, 4.856738, 4.843309, 4.831854, 4.823215, 
    4.818036, 4.816703, 4.819304, 4.825633, 4.835196, 4.847248, 4.860843, 
    4.874875, 4.888161, 4.899525, 4.907917, 4.912551, 4.913051, 4.909559, 
    4.9028,
  // momentumX(17,42, 0-49)
    4.909159, 4.904336, 4.901761, 4.901208, 4.902383, 4.904947, 4.90855, 
    4.912868, 4.917612, 4.922549, 4.9275, 4.932313, 4.936859, 4.940983, 
    4.944482, 4.945125, 4.954541, 4.955351, 4.954765, 4.953189, 4.95065, 
    4.950379, 4.948419, 4.945224, 4.939711, 4.931865, 4.921547, 4.909028, 
    4.894497, 4.879364, 4.863691, 4.851813, 4.841222, 4.832664, 4.826799, 
    4.8241, 4.824811, 4.828923, 4.836165, 4.846019, 4.857746, 4.870423, 
    4.883003, 4.894386, 4.903529, 4.90956, 4.911921, 4.910494, 4.905684, 
    4.898421,
  // momentumX(17,43, 0-49)
    4.914628, 4.909033, 4.905563, 4.904037, 4.904203, 4.905764, 4.908397, 
    4.91179, 4.915656, 4.919752, 4.923867, 4.927831, 4.931473, 4.934608, 
    4.936998, 4.937302, 4.946457, 4.946009, 4.944318, 4.94176, 4.938349, 
    4.937307, 4.934862, 4.93152, 4.926051, 4.91854, 4.908878, 4.897394, 
    4.884263, 4.871099, 4.857931, 4.848797, 4.84109, 4.835384, 4.832156, 
    4.83172, 4.834194, 4.839475, 4.847241, 4.856964, 4.867921, 4.879242, 
    4.889966, 4.899126, 4.905847, 4.909483, 4.909735, 4.906756, 4.901185, 
    4.894104,
  // momentumX(17,44, 0-49)
    4.919461, 4.912925, 4.908408, 4.905779, 4.904836, 4.90532, 4.90694, 
    4.909394, 4.912395, 4.915678, 4.919009, 4.92218, 4.924991, 4.92723, 
    4.928645, 4.928577, 4.937214, 4.935669, 4.933005, 4.929586, 4.925431, 
    4.923725, 4.920937, 4.917611, 4.91241, 4.905505, 4.896807, 4.88668, 
    4.875265, 4.864319, 4.85382, 4.847488, 4.84264, 4.839678, 4.838911, 
    4.8405, 4.844442, 4.850554, 4.858476, 4.867672, 4.877462, 4.887057, 
    4.895621, 4.902356, 4.906611, 4.907991, 4.906475, 4.902468, 4.896797, 
    4.890616,
  // momentumX(17,45, 0-49)
    4.924008, 4.916375, 4.910664, 4.906796, 4.904622, 4.903929, 4.904456, 
    4.905918, 4.908018, 4.910478, 4.913033, 4.91544, 4.91747, 4.918889, 
    4.919441, 4.918964, 4.926886, 4.924419, 4.920935, 4.916797, 4.912052, 
    4.909824, 4.906849, 4.903707, 4.898986, 4.892923, 4.885447, 4.876929, 
    4.86746, 4.858889, 4.851131, 4.847575, 4.845493, 4.84512, 4.846608, 
    4.849974, 4.855102, 4.861737, 4.869482, 4.877822, 4.886137, 4.893749, 
    4.899987, 4.904269, 4.906194, 4.90565, 4.902875, 4.898486, 4.893424, 
    4.888831,
  // momentumX(17,46, 0-49)
    4.928825, 4.919962, 4.912918, 4.90767, 4.904126, 4.902122, 4.90143, 
    4.901784, 4.902892, 4.904456, 4.906185, 4.907807, 4.909061, 4.909698, 
    4.909465, 4.908536, 4.915604, 4.912388, 4.908238, 4.903537, 4.898368, 
    4.895784, 4.892784, 4.88998, 4.885921, 4.880892, 4.874827, 4.868092, 
    4.860718, 4.854588, 4.849548, 4.848677, 4.849215, 4.851243, 4.854764, 
    4.859663, 4.865725, 4.87262, 4.879941, 4.887194, 4.89385, 4.899375, 
    4.903301, 4.905291, 4.905223, 4.903256, 4.899861, 4.895799, 4.892039, 
    4.889628,
  // momentumX(17,47, 0-49)
    4.934628, 4.924436, 4.915936, 4.909171, 4.904103, 4.900622, 4.898542, 
    4.897622, 4.897577, 4.898103, 4.89889, 4.899638, 4.900064, 4.899903, 
    4.898912, 4.897471, 4.903601, 4.899779, 4.895105, 4.889996, 4.884573, 
    4.881795, 4.878922, 4.876583, 4.873326, 4.869465, 4.864933, 4.860072, 
    4.85486, 4.851156, 4.848743, 4.850405, 4.853375, 4.857594, 4.862926, 
    4.869143, 4.875928, 4.882905, 4.889649, 4.895721, 4.900694, 4.904212, 
    4.906034, 4.906089, 4.904534, 4.901772, 4.898455, 4.895413, 4.893567, 
    4.893793,
  // momentumX(17,48, 0-49)
    4.942206, 4.930628, 4.920584, 4.912177, 4.905432, 4.900293, 4.896624, 
    4.894217, 4.892807, 4.892093, 4.891754, 4.891472, 4.890954, 4.889923, 
    4.888144, 4.886106, 4.891249, 4.886915, 4.881835, 4.876449, 4.870919, 
    4.868098, 4.865475, 4.863686, 4.861314, 4.858688, 4.855734, 4.852766, 
    4.84971, 4.848352, 4.848417, 4.852421, 4.857611, 4.863803, 4.870745, 
    4.878098, 4.885471, 4.89244, 4.898585, 4.903532, 4.906981, 4.908762, 
    4.908873, 4.907512, 4.905091, 4.902219, 4.899659, 4.898243, 4.898774, 
    4.901918,
  // momentumX(17,49, 0-49)
    4.959617, 4.946238, 4.934052, 4.923233, 4.913883, 4.906022, 4.89959, 
    4.894449, 4.890389, 4.887144, 4.884412, 4.881876, 4.879222, 4.876143, 
    4.872361, 4.869101, 4.880398, 4.874001, 4.866947, 4.860031, 4.853502, 
    4.852767, 4.852791, 4.85458, 4.855067, 4.854731, 4.853221, 4.850918, 
    4.847435, 4.846223, 4.846673, 4.853611, 4.861576, 4.870242, 4.879228, 
    4.888075, 4.896299, 4.903437, 4.909089, 4.912979, 4.914989, 4.915207, 
    4.913942, 4.911713, 4.909215, 4.907247, 4.906631, 4.908108, 4.91226, 
    4.919442,
  // momentumX(18,0, 0-49)
    4.884809, 4.871144, 4.860725, 4.853534, 4.849423, 4.848121, 4.849251, 
    4.852354, 4.856926, 4.862458, 4.868456, 4.874484, 4.880164, 4.885192, 
    4.88933, 4.892411, 4.895638, 4.896484, 4.896322, 4.895182, 4.893073, 
    4.890365, 4.886718, 4.882278, 4.87701, 4.871042, 4.864499, 4.857598, 
    4.850573, 4.843819, 4.837571, 4.832456, 4.82845, 4.825788, 4.824625, 
    4.825011, 4.826875, 4.830015, 4.834108, 4.838731, 4.843399, 4.84762, 
    4.850959, 4.853108, 4.853957, 4.853652, 4.852622, 4.851551, 4.851324, 
    4.852911,
  // momentumX(18,1, 0-49)
    4.884934, 4.871832, 4.862022, 4.855465, 4.85199, 4.851309, 4.853025, 
    4.856676, 4.861752, 4.867746, 4.874176, 4.880609, 4.886672, 4.892051, 
    4.896487, 4.899747, 4.904272, 4.905182, 4.905079, 4.903979, 4.901849, 
    4.899334, 4.895684, 4.891092, 4.885404, 4.878729, 4.871161, 4.862932, 
    4.854278, 4.845744, 4.837555, 4.830768, 4.825129, 4.820971, 4.818543, 
    4.817976, 4.819256, 4.822213, 4.826527, 4.831753, 4.837351, 4.842746, 
    4.847396, 4.850862, 4.852898, 4.853511, 4.853005, 4.851987, 4.851309, 
    4.851967,
  // momentumX(18,2, 0-49)
    4.886409, 4.873914, 4.864717, 4.858756, 4.855839, 4.85566, 4.857812, 
    4.861832, 4.867219, 4.87348, 4.880151, 4.886819, 4.893123, 4.898752, 
    4.903427, 4.906798, 4.912543, 4.913613, 4.913682, 4.912762, 4.910775, 
    4.908639, 4.905188, 4.900646, 4.894743, 4.887562, 4.879149, 4.869736, 
    4.859549, 4.849249, 4.839058, 4.830468, 4.823002, 4.817106, 4.813138, 
    4.811329, 4.811743, 4.814265, 4.818604, 4.82431, 4.830813, 4.837478, 
    4.84367, 4.848833, 4.852573, 4.854734, 4.855453, 4.855189, 4.854686, 
    4.854899,
  // momentumX(18,3, 0-49)
    4.888647, 4.876785, 4.868192, 4.862783, 4.86035, 4.860566, 4.863028, 
    4.867271, 4.872816, 4.879192, 4.885966, 4.892745, 4.899195, 4.905011, 
    4.909902, 4.913323, 4.920159, 4.921499, 4.921853, 4.921245, 4.919561, 
    4.917976, 4.914915, 4.910623, 4.904731, 4.897276, 4.888249, 4.877862, 
    4.866318, 4.854356, 4.842188, 4.831735, 4.822308, 4.814471, 4.808708, 
    4.805367, 4.804612, 4.806405, 4.810504, 4.816482, 4.823758, 4.831663, 
    4.839493, 4.846585, 4.852404, 4.856616, 4.859165, 4.860306, 4.860612, 
    4.860924,
  // momentumX(18,4, 0-49)
    4.89114, 4.879928, 4.871926, 4.867028, 4.865009, 4.865537, 4.868205, 
    4.872565, 4.878159, 4.884547, 4.891326, 4.898142, 4.904681, 4.910653, 
    4.915773, 4.919184, 4.926921, 4.92865, 4.929398, 4.929215, 4.927966, 
    4.927078, 4.924573, 4.920717, 4.91506, 4.907583, 4.898214, 4.887125, 
    4.874485, 4.861058, 4.847029, 4.834742, 4.823296, 4.813377, 4.805604, 
    4.800458, 4.798227, 4.798971, 4.802519, 4.808488, 4.816317, 4.825317, 
    4.834739, 4.843832, 4.851933, 4.858536, 4.863369, 4.866457, 4.868152, 
    4.869117,
  // momentumX(18,5, 0-49)
    4.893487, 4.882936, 4.875515, 4.871094, 4.869439, 4.870214, 4.873019, 
    4.877421, 4.882993, 4.889328, 4.89606, 4.90287, 4.909472, 4.915598, 
    4.920979, 4.924315, 4.932712, 4.934937, 4.936172, 4.936502, 4.935794, 
    4.935705, 4.933889, 4.930626, 4.925414, 4.918171, 4.908759, 4.897293, 
    4.883885, 4.869284, 4.853611, 4.839611, 4.826176, 4.814109, 4.80417, 
    4.796988, 4.792989, 4.792358, 4.795018, 4.800653, 4.808738, 4.818592, 
    4.829433, 4.840447, 4.85086, 4.860002, 4.867395, 4.872821, 4.876379, 
    4.878513,
  // momentumX(18,6, 0-49)
    4.895404, 4.88553, 4.878681, 4.874718, 4.873394, 4.874374, 4.877271, 
    4.881673, 4.887185, 4.893434, 4.900091, 4.906876, 4.913533, 4.919827, 
    4.925513, 4.928716, 4.937472, 4.940289, 4.942079, 4.942984, 4.942886, 
    4.94365, 4.942612, 4.940061, 4.935476, 4.928711, 4.919563, 4.908076, 
    4.894294, 4.878877, 4.861876, 4.846375, 4.831077, 4.816886, 4.8047, 
    4.795306, 4.789286, 4.78697, 4.788401, 4.79335, 4.801349, 4.811738, 
    4.823725, 4.836451, 4.849043, 4.860695, 4.870737, 4.878716, 4.884475, 
    4.888203,
  // momentumX(18,7, 0-49)
    4.896717, 4.887537, 4.881267, 4.877753, 4.876744, 4.877908, 4.880875, 
    4.885259, 4.890693, 4.896843, 4.903419, 4.910171, 4.916884, 4.92336, 
    4.929397, 4.932419, 4.941206, 4.944678, 4.947065, 4.948576, 4.949125, 
    4.950751, 4.950533, 4.948766, 4.944954, 4.938883, 4.930294, 4.919146, 
    4.905412, 4.889598, 4.871658, 4.854958, 4.838015, 4.821816, 4.807391, 
    4.795682, 4.787444, 4.783171, 4.783046, 4.786955, 4.794499, 4.80506, 
    4.81785, 4.831971, 4.846484, 4.860461, 4.873067, 4.88364, 4.891777, 
    4.897409,
  // momentumX(18,8, 0-49)
    4.897334, 4.888876, 4.8832, 4.880144, 4.879449, 4.880795, 4.88383, 
    4.888193, 4.893551, 4.899602, 4.906095, 4.912813, 4.919581, 4.926244, 
    4.932665, 4.935491, 4.943973, 4.948122, 4.951126, 4.953247, 4.954448, 
    4.956897, 4.957495, 4.956541, 4.953597, 4.948393, 4.940624, 4.930164, 
    4.916898, 4.901135, 4.882703, 4.865164, 4.846878, 4.828883, 4.812316, 
    4.798274, 4.78769, 4.78124, 4.779273, 4.781801, 4.788523, 4.798871, 
    4.812071, 4.82721, 4.843288, 4.859285, 4.874232, 4.887288, 4.897826, 
    4.905539,
  // momentumX(18,9, 0-49)
    4.897227, 4.889523, 4.884467, 4.881888, 4.881528, 4.883073, 4.886189, 
    4.890546, 4.895837, 4.901796, 4.908204, 4.914883, 4.921696, 4.928542, 
    4.935356, 4.938022, 4.945889, 4.950691, 4.9543, 4.957017, 4.958854, 
    4.962049, 4.963417, 4.963258, 4.96123, 4.957014, 4.950277, 4.940805, 
    4.928404, 4.913132, 4.894676, 4.876698, 4.85743, 4.837928, 4.819408, 
    4.803104, 4.790129, 4.78135, 4.777303, 4.778151, 4.783701, 4.793451, 
    4.806657, 4.822395, 4.839628, 4.857264, 4.874227, 4.889527, 4.902359, 
    4.912195,
  // momentumX(18,10, 0-49)
    4.896404, 4.88949, 4.885093, 4.883026, 4.883033, 4.884808, 4.888037, 
    4.892411, 4.897654, 4.903532, 4.909855, 4.916485, 4.923323, 4.930325, 
    4.937502, 4.940127, 4.947123, 4.952506, 4.956683, 4.959964, 4.962405, 
    4.966238, 4.968298, 4.968881, 4.967768, 4.964606, 4.959049, 4.950807, 
    4.939605, 4.925227, 4.90721, 4.889191, 4.869336, 4.848673, 4.828465, 
    4.810056, 4.79473, 4.783552, 4.777253, 4.776168, 4.780232, 4.789024, 
    4.80184, 4.817754, 4.835709, 4.854557, 4.873146, 4.890373, 4.905285, 
    4.917168,
  // momentumX(18,11, 0-49)
    4.894901, 4.888815, 4.885118, 4.88361, 4.884029, 4.886082, 4.889462, 
    4.893889, 4.899112, 4.904922, 4.911164, 4.917727, 4.924558, 4.931664, 
    4.939128, 4.941932, 4.947885, 4.95373, 4.958413, 4.962218, 4.965225, 
    4.969569, 4.972219, 4.97346, 4.973217, 4.971121, 4.966827, 4.95998, 
    4.950234, 4.937087, 4.91993, 4.90224, 4.882188, 4.860743, 4.839166, 
    4.818886, 4.801331, 4.787762, 4.779115, 4.775909, 4.778225, 4.785737, 
    4.797791, 4.813478, 4.831725, 4.851353, 4.87115, 4.889936, 4.906639, 
    4.920398,
  // momentumX(18,12, 0-49)
    4.892765, 4.88754, 4.884587, 4.88369, 4.884581, 4.886966, 4.890554, 
    4.89508, 4.900316, 4.906077, 4.912237, 4.918715, 4.925493, 4.932621, 
    4.940238, 4.94356, 4.948406, 4.954556, 4.959667, 4.963951, 4.967489, 
    4.972205, 4.97533, 4.977124, 4.977676, 4.976608, 4.973598, 4.968228, 
    4.960105, 4.94844, 4.9325, 4.915447, 4.895557, 4.873702, 4.851109, 
    4.829243, 4.809653, 4.793781, 4.782765, 4.777319, 4.777685, 4.783647, 
    4.794613, 4.809704, 4.827843, 4.847833, 4.868425, 4.888381, 4.906549, 
    4.921947,
  // momentumX(18,13, 0-49)
    4.890054, 4.885715, 4.88355, 4.883318, 4.884742, 4.887525, 4.891382, 
    4.89606, 4.901348, 4.907085, 4.913165, 4.919536, 4.926205, 4.93325, 
    4.940831, 4.945117, 4.948902, 4.955187, 4.960639, 4.96536, 4.969398, 
    4.97435, 4.977834, 4.980072, 4.981319, 4.981205, 4.979434, 4.975549, 
    4.969117, 4.959093, 4.944644, 4.928452, 4.909022, 4.887101, 4.86384, 
    4.840705, 4.81933, 4.801309, 4.787976, 4.780247, 4.778527, 4.782729, 
    4.792338, 4.806513, 4.824186, 4.844155, 4.865149, 4.885897, 4.905189, 
    4.921952,
  // momentumX(18,14, 0-49)
    4.886841, 4.883399, 4.882051, 4.882535, 4.884551, 4.887797, 4.891985, 
    4.896872, 4.902257, 4.907996, 4.914003, 4.920245, 4.926744, 4.933584, 
    4.940909, 4.94667, 4.949551, 4.95581, 4.961526, 4.966652, 4.971175, 
    4.976239, 4.979972, 4.982547, 4.984378, 4.98511, 4.984487, 4.982019, 
    4.977257, 4.968933, 4.956161, 4.94096, 4.922206, 4.900504, 4.876897, 
    4.852814, 4.829932, 4.809971, 4.794442, 4.784451, 4.780582, 4.782882, 
    4.790926, 4.803923, 4.820827, 4.840441, 4.861489, 4.882676, 4.90276, 
    4.920603,
  // momentumX(18,15, 0-49)
    4.883207, 4.880651, 4.880136, 4.881371, 4.884029, 4.887794, 4.892372, 
    4.897519, 4.903045, 4.908817, 4.914763, 4.920861, 4.927134, 4.93365, 
    4.940502, 4.948238, 4.950455, 4.956568, 4.962499, 4.96802, 4.973034, 
    4.978105, 4.982003, 4.984821, 4.987122, 4.988574, 4.988962, 4.987782, 
    4.984583, 4.977922, 4.966918, 4.952744, 4.934793, 4.913519, 4.889838, 
    4.865107, 4.84101, 4.819353, 4.801796, 4.789631, 4.783615, 4.783937, 
    4.790273, 4.801894, 4.817789, 4.836773, 4.857575, 4.878895, 4.899468, 
    4.918118,
  // momentumX(18,16, 0-49)
    4.879242, 4.87754, 4.87785, 4.879844, 4.883172, 4.887492, 4.892501, 
    4.897952, 4.903658, 4.909498, 4.915406, 4.921362, 4.92738, 4.933488, 
    4.939705, 4.949776, 4.951613, 4.95754, 4.963687, 4.969635, 4.975175, 
    4.98018, 4.984186, 4.987179, 4.989842, 4.991875, 4.993103, 4.993021, 
    4.991203, 4.986084, 4.976843, 4.963641, 4.946527, 4.925811, 4.902266, 
    4.877148, 4.852115, 4.829021, 4.809649, 4.795449, 4.787349, 4.785682, 
    4.790234, 4.800347, 4.815056, 4.8332, 4.853517, 4.874714, 4.895517, 
    4.914725,
  // momentumX(18,17, 0-49)
    4.875041, 4.874127, 4.875218, 4.87795, 4.881939, 4.886819, 4.892274, 
    4.898053, 4.903974, 4.909922, 4.915837, 4.921696, 4.927484, 4.933181, 
    4.938707, 4.951196, 4.952917, 4.958723, 4.965165, 4.971624, 4.977774, 
    4.982686, 4.986784, 4.989913, 4.992849, 4.995311, 4.997171, 4.997947, 
    4.997252, 4.993465, 4.9859, 4.973534, 4.95721, 4.937099, 4.913828, 
    4.888538, 4.862826, 4.838557, 4.817604, 4.801552, 4.791484, 4.787878, 
    4.790633, 4.799174, 4.812584, 4.829738, 4.849395, 4.870271, 4.891096, 
    4.910655,
  // momentumX(18,18, 0-49)
    4.870688, 4.87046, 4.872247, 4.875643, 4.880235, 4.885635, 4.891515, 
    4.897624, 4.90379, 4.909906, 4.91592, 4.921796, 4.927487, 4.932893, 
    4.937829, 4.952391, 4.954152, 4.960028, 4.966936, 4.974069, 4.980973, 
    4.985815, 4.99005, 4.993322, 4.99646, 4.999198, 5.001451, 5.002779, 
    5.002877, 5.000129, 4.994055, 4.982319, 4.966665, 4.947137, 4.924218, 
    4.898921, 4.872756, 4.847573, 4.825289, 4.807601, 4.795727, 4.790283, 
    4.791286, 4.798248, 4.810311, 4.826389, 4.84527, 4.865687, 4.886379, 
    4.906126,
  // momentumX(18,19, 0-49)
    4.86625, 4.86655, 4.868883, 4.872808, 4.877879, 4.883698, 4.889936, 
    4.896357, 4.902807, 4.909202, 4.915492, 4.921624, 4.927492, 4.932897, 
    4.937518, 4.953274, 4.955041, 4.961284, 4.968928, 4.976991, 4.984876, 
    4.989754, 4.994244, 4.997727, 5.001033, 5.003887, 5.006248, 5.007756, 
    5.008227, 5.006122, 5.001248, 4.98988, 4.974717, 4.955695, 4.933158, 
    4.907983, 4.881572, 4.855722, 4.832371, 4.813286, 4.799805, 4.792671, 
    4.792016, 4.797443, 4.808165, 4.823141, 4.841189, 4.861065, 4.881521, 
    4.901341,
  // momentumX(18,20, 0-49)
    4.862615, 4.864183, 4.867981, 4.873559, 4.880429, 4.888097, 4.896105, 
    4.904039, 4.91155, 4.918352, 4.924236, 4.929071, 4.932817, 4.935514, 
    4.937287, 0, 4.967083, 4.970193, 4.974487, 4.979447, 4.9848, 4.986744, 
    4.989418, 4.992031, 4.995424, 4.999174, 5.003032, 5.006403, 5.008925, 
    5.008933, 5.006418, 4.996209, 4.982046, 4.963815, 4.941799, 4.916811, 
    4.8902, 4.86374, 4.83939, 4.818989, 4.803974, 4.79521, 4.792936, 
    4.796848, 4.806228, 4.820079, 4.837255, 4.856534, 4.87668, 4.896485,
  // momentumX(18,21, 0-49)
    4.858526, 4.860593, 4.864909, 4.870983, 4.878288, 4.886311, 4.89458, 
    4.902694, 4.910328, 4.917231, 4.923228, 4.928211, 4.932137, 4.935033, 
    4.936998, 0, 4.96749, 4.971151, 4.976059, 4.981626, 4.987492, 4.988534, 
    4.990527, 4.992525, 4.995533, 4.999171, 5.003212, 5.007048, 5.010316, 
    5.011328, 5.010325, 5.000771, 4.987464, 4.970185, 4.949078, 4.924807, 
    4.898589, 4.872103, 4.847268, 4.82596, 4.809701, 4.799472, 4.795639, 
    4.798006, 4.805933, 4.818489, 4.834568, 4.852976, 4.872499, 4.891943,
  // momentumX(18,22, 0-49)
    4.854605, 4.857058, 4.861805, 4.868328, 4.876069, 4.884493, 4.893115, 
    4.901526, 4.909408, 4.916522, 4.922707, 4.927864, 4.931949, 4.93498, 
    4.937038, 0, 4.968196, 4.972306, 4.977769, 4.98394, 4.990365, 4.990649, 
    4.992125, 4.993677, 4.996429, 5.000011, 5.004191, 5.008338, 5.01208, 
    5.013722, 5.013745, 5.004387, 4.991473, 4.974729, 4.954206, 4.930459, 
    4.904589, 4.878174, 4.853073, 4.831153, 4.813982, 4.802622, 4.797538, 
    4.798625, 4.805327, 4.816769, 4.831888, 4.849522, 4.86848, 4.887581,
  // momentumX(18,23, 0-49)
    4.850917, 4.853661, 4.858761, 4.865675, 4.873829, 4.882668, 4.891686, 
    4.900468, 4.908682, 4.916094, 4.922538, 4.927917, 4.932185, 4.935344, 
    4.93747, 0, 4.969583, 4.973991, 4.979832, 4.98642, 4.993236, 4.992826, 
    4.993824, 4.99496, 4.99745, 5.000928, 5.005152, 5.009469, 5.013495, 
    5.015525, 5.016229, 5.006853, 4.994095, 4.977653, 4.95752, 4.934175, 
    4.908624, 4.882356, 4.857164, 4.834885, 4.817104, 4.804931, 4.798903, 
    4.798989, 4.804698, 4.81521, 4.8295, 4.846437, 4.864852, 4.883585,
  // momentumX(18,24, 0-49)
    4.847519, 4.850479, 4.85586, 4.863112, 4.871647, 4.880895, 4.890332, 
    4.899526, 4.908134, 4.915905, 4.92267, 4.928324, 4.932813, 4.936135, 
    4.938357, 0, 4.971826, 4.976392, 4.982431, 4.989242, 4.996271, 4.995375, 
    4.996037, 4.996878, 4.999168, 5.002536, 5.006739, 5.011106, 5.015255, 
    5.017463, 5.018531, 5.009044, 4.996279, 4.979924, 4.959941, 4.936765, 
    4.911347, 4.885115, 4.859817, 4.837259, 4.819028, 4.806264, 4.799543, 
    4.798884, 4.803843, 4.813639, 4.827281, 4.843661, 4.86163, 4.880041,
  // momentumX(18,25, 0-49)
    4.84447, 4.847589, 4.853196, 4.860741, 4.869628, 4.879272, 4.889136, 
    4.898769, 4.907809, 4.915988, 4.923122, 4.929097, 4.933853, 4.937385, 
    4.939763, 0, 4.974479, 4.979081, 4.985147, 4.991983, 4.999034, 4.997939, 
    4.99846, 4.999179, 5.001375, 5.00467, 5.008821, 5.013151, 5.017279, 
    5.019472, 5.020578, 5.010951, 4.998077, 4.981641, 4.961603, 4.938382, 
    4.91291, 4.88659, 4.861147, 4.838369, 4.819839, 4.806698, 4.799538, 
    4.7984, 4.802862, 4.81217, 4.825348, 4.841312, 4.858924, 4.877048,
  // momentumX(18,26, 0-49)
    4.841846, 4.845082, 4.850876, 4.858679, 4.867893, 4.877924, 4.888223, 
    4.898314, 4.907815, 4.916437, 4.923976, 4.930305, 4.935359, 4.939139, 
    4.941726, 0, 4.977385, 4.981901, 4.98783, 4.994493, 5.001371, 5.000391, 
    5.000994, 5.001788, 5.004019, 5.007303, 5.01139, 5.015614, 5.019589, 
    5.021584, 5.022406, 5.012643, 4.999584, 4.982924, 4.962636, 4.939158, 
    4.913439, 4.886895, 4.861254, 4.838302, 4.819606, 4.806296, 4.798949, 
    4.797599, 4.801824, 4.810872, 4.823782, 4.839473, 4.856821, 4.874699,
  // momentumX(18,27, 0-49)
    4.839744, 4.843068, 4.84902, 4.857059, 4.866587, 4.877005, 4.887747, 
    4.898317, 4.908307, 4.917399, 4.925366, 4.932062, 4.937419, 4.941448, 
    4.944248, 0, 4.980576, 4.984866, 4.990472, 4.996755, 5.003257, 5.002659, 
    5.003529, 5.004568, 5.006943, 5.01026, 5.014267, 5.018305, 5.021995, 
    5.023608, 5.023826, 5.013915, 5.000586, 4.983556, 4.962839, 4.938921, 
    4.912803, 4.885948, 4.860112, 4.837081, 4.818402, 4.805168, 4.797915, 
    4.796639, 4.800896, 4.809918, 4.822744, 4.838297, 4.855458, 4.873108,
  // momentumX(18,28, 0-49)
    4.838279, 4.841671, 4.847761, 4.856022, 4.86586, 4.876674, 4.887884, 
    4.898968, 4.909482, 4.919071, 4.927473, 4.934519, 4.940135, 4.94435, 
    4.94729, 0, 4.984393, 4.988278, 4.993347, 4.999027, 5.004954, 5.004905, 
    5.006158, 5.007552, 5.010141, 5.013506, 5.017393, 5.021155, 5.024417, 
    5.025462, 5.024777, 5.014656, 5.000932, 4.983361, 4.962024, 4.937493, 
    4.910855, 4.883649, 4.857671, 4.834711, 4.816276, 4.803395, 4.796536, 
    4.795633, 4.800196, 4.80943, 4.82236, 4.837905, 4.854949, 4.872379,
  // momentumX(18,29, 0-49)
    4.837578, 4.841016, 4.847223, 4.855696, 4.865859, 4.8771, 4.888828, 
    4.900484, 4.911574, 4.921689, 4.930514, 4.937848, 4.943614, 4.94786, 
    4.950751, 0, 4.988549, 4.991818, 4.996123, 5.000973, 5.006124, 5.006631, 
    5.00827, 5.010037, 5.012847, 5.016247, 5.019962, 5.023355, 5.02604, 
    5.026312, 5.024417, 5.013925, 4.999619, 4.981328, 4.959243, 4.93405, 
    4.906947, 4.879553, 4.853701, 4.831154, 4.813352, 4.801226, 4.795144, 
    4.794957, 4.800112, 4.80978, 4.822963, 4.83858, 4.855508, 4.872646,
  // momentumX(18,30, 0-49)
    4.837201, 4.839952, 4.84534, 4.852841, 4.861905, 4.872, 4.882656, 
    4.893489, 4.904216, 4.914642, 4.924639, 4.934104, 4.942914, 4.950874, 
    4.957664, 4.980512, 4.978384, 4.985451, 4.993881, 5.002621, 5.011064, 
    5.015289, 5.019503, 5.022801, 5.026014, 5.028763, 5.03095, 5.032186, 
    5.032328, 5.02988, 5.02498, 5.012665, 4.996644, 4.97683, 4.95351, 
    4.927465, 4.899968, 4.872666, 4.847361, 4.825732, 4.809091, 4.798231, 
    4.793395, 4.794331, 4.800419, 4.81079, 4.824425, 4.840233, 4.8571, 
    4.873925,
  // momentumX(18,31, 0-49)
    4.838711, 4.841673, 4.847275, 4.855004, 4.864307, 4.874646, 4.885531, 
    4.896559, 4.907419, 4.917896, 4.927857, 4.937228, 4.945951, 4.953948, 
    4.961065, 4.980995, 4.980417, 4.987096, 4.994756, 5.002519, 5.00993, 
    5.014159, 5.018117, 5.021186, 5.024208, 5.026828, 5.028913, 5.029993, 
    5.029801, 5.02675, 5.020671, 5.008065, 4.991631, 4.971384, 4.94774, 
    4.9216, 4.89433, 4.86762, 4.843251, 4.822825, 4.807539, 4.798059, 
    4.794508, 4.796546, 4.803485, 4.814416, 4.828295, 4.844025, 4.860487, 
    4.876597,
  // momentumX(18,32, 0-49)
    4.841342, 4.844412, 4.850084, 4.857855, 4.867183, 4.877531, 4.888418, 
    4.899436, 4.910273, 4.920713, 4.930632, 4.93998, 4.948754, 4.956964, 
    4.964594, 4.980965, 4.981505, 4.988069, 4.995195, 5.002202, 5.00878, 
    5.013144, 5.016983, 5.019907, 5.02272, 5.025066, 5.026776, 5.02734, 
    5.026409, 5.022374, 5.014822, 5.001704, 4.984722, 4.964009, 4.940114, 
    4.914057, 4.88728, 4.861488, 4.838411, 4.819547, 4.80595, 4.798151, 
    4.796151, 4.799515, 4.807491, 4.819123, 4.833344, 4.849035, 4.865076, 
    4.880392,
  // momentumX(18,33, 0-49)
    4.845201, 4.848296, 4.853919, 4.861576, 4.870737, 4.880888, 4.891561, 
    4.902365, 4.912999, 4.923262, 4.933043, 4.942318, 4.951126, 4.959552, 
    4.967697, 4.980441, 4.981912, 4.988523, 4.995258, 5.001646, 5.007523, 
    5.012081, 5.015876, 5.018697, 5.021259, 5.023195, 5.024305, 5.02406, 
    5.022061, 5.016749, 5.007536, 4.993733, 4.976113, 4.954939, 4.930896, 
    4.905118, 4.879101, 4.85454, 4.833084, 4.816096, 4.804484, 4.798627, 
    4.798405, 4.803288, 4.812459, 4.824915, 4.839553, 4.855231, 4.870821, 
    4.885258,
  // momentumX(18,34, 0-49)
    4.850313, 4.853356, 4.858818, 4.866215, 4.875041, 4.884804, 4.895066, 
    4.905462, 4.915716, 4.925641, 4.935148, 4.944232, 4.952967, 4.961494, 
    4.970001, 4.979457, 4.981847, 4.98854, 4.994935, 5.000776, 5.006025, 
    5.010772, 5.014541, 5.01726, 5.019513, 5.020917, 5.02124, 5.019953, 
    5.016633, 5.00984, 4.998881, 4.98429, 4.966008, 4.944437, 4.920403, 
    4.895131, 4.870153, 4.847122, 4.82758, 4.812739, 4.803346, 4.799632, 
    4.801355, 4.8079, 4.818378, 4.831736, 4.846831, 4.862496, 4.877587, 
    4.891049,
  // momentumX(18,35, 0-49)
    4.85662, 4.859527, 4.864711, 4.871711, 4.880044, 4.889249, 4.898926, 
    4.908741, 4.918445, 4.927876, 4.936965, 4.94572, 4.954232, 4.962675, 
    4.971297, 4.978046, 4.981433, 4.988136, 4.99417, 4.999484, 5.004143, 
    5.009024, 5.012743, 5.015333, 5.017207, 5.017971, 5.017355, 5.014852, 
    5.01003, 5.001642, 4.988949, 4.973538, 4.954648, 4.932821, 4.909005, 
    4.884502, 4.860847, 4.839624, 4.822244, 4.809759, 4.80275, 4.801305, 
    4.805072, 4.813345, 4.825176, 4.839457, 4.855005, 4.870616, 4.885136, 
    4.89752,
  // momentumX(18,36, 0-49)
    4.863973, 4.866647, 4.871443, 4.877914, 4.885613, 4.894113, 4.903052, 
    4.912133, 4.921141, 4.929941, 4.938475, 4.946762, 4.954895, 4.963057, 
    4.971507, 4.97621, 4.980695, 4.987263, 4.992869, 4.997642, 5.001723, 
    5.006649, 5.010259, 5.012672, 5.014094, 5.014126, 5.01246, 5.008624, 
    5.0022, 4.992191, 4.977875, 4.961699, 4.942339, 4.920467, 4.897135, 
    4.87369, 4.85164, 4.83247, 4.817447, 4.807454, 4.802914, 4.80378, 
    4.809597, 4.819584, 4.832732, 4.847884, 4.863813, 4.879286, 4.893135, 
    4.904335,
  // momentumX(18,37, 0-49)
    4.872146, 4.874485, 4.878777, 4.884603, 4.891544, 4.899216, 4.907293, 
    4.91552, 4.923715, 4.931767, 4.939631, 4.947328, 4.954942, 4.962633, 
    4.970646, 4.973928, 4.979574, 4.985822, 4.990914, 4.995116, 4.99861, 
    5.003463, 5.006887, 5.00906, 5.009962, 5.009189, 5.006405, 5.001185, 
    4.993144, 4.981586, 4.965855, 4.949062, 4.929453, 4.907815, 4.885276, 
    4.863191, 4.843011, 4.8261, 4.813562, 4.806119, 4.804044, 4.807168, 
    4.814948, 4.826537, 4.840876, 4.856761, 4.872931, 4.888124, 4.901169, 
    4.911073,
  // momentumX(18,38, 0-49)
    4.880842, 4.882741, 4.886423, 4.891498, 4.897586, 4.904336, 4.911465, 
    4.918751, 4.926048, 4.933264, 4.940367, 4.947376, 4.954354, 4.961426, 
    4.968778, 4.971156, 4.977955, 4.983696, 4.988179, 4.991767, 4.994656, 
    4.999306, 5.002451, 5.004314, 5.004631, 5.003013, 4.999096, 4.992517, 
    4.982934, 4.969998, 4.953146, 4.935975, 4.916419, 4.895351, 4.873941, 
    4.853517, 4.83544, 4.820933, 4.810941, 4.806021, 4.806313, 4.811546, 
    4.821102, 4.834083, 4.849388, 4.86578, 4.881971, 4.896688, 4.908768, 
    4.917272,
  // momentumX(18,39, 0-49)
    4.889717, 4.891066, 4.894044, 4.898291, 4.903454, 4.909225, 4.915352, 
    4.921652, 4.927999, 4.934326, 4.940608, 4.946858, 4.953117, 4.959458, 
    4.965996, 4.96784, 4.975702, 4.980766, 4.984552, 4.987484, 4.989732, 
    4.99404, 4.996809, 4.998293, 4.997983, 4.995514, 4.990504, 4.982667, 
    4.971714, 4.957668, 4.940073, 4.922842, 4.903699, 4.883575, 4.863635, 
    4.84515, 4.829363, 4.817347, 4.809879, 4.807374, 4.809848, 4.816947, 
    4.827996, 4.842059, 4.858009, 4.874594, 4.890515, 4.904504, 4.915439, 
    4.922453,
  // momentumX(18,40, 0-49)
    4.8984, 4.899097, 4.90129, 4.904646, 4.908849, 4.913617, 4.91873, 
    4.924032, 4.929419, 4.934838, 4.940274, 4.945725, 4.951211, 4.956755, 
    4.96239, 4.963936, 4.972683, 4.976931, 4.979949, 4.982178, 4.983747, 
    4.987577, 4.989875, 4.990921, 4.989964, 4.98668, 4.98068, 4.971765, 
    4.959704, 4.944898, 4.927004, 4.910091, 4.891764, 4.872965, 4.854824, 
    4.838517, 4.825151, 4.815638, 4.810602, 4.81032, 4.814709, 4.823346, 
    4.835516, 4.850266, 4.866456, 4.882841, 4.898137, 4.911113, 4.920713, 
    4.926178,
  // momentumX(18,41, 0-49)
    4.906529, 4.906476, 4.907814, 4.910242, 4.91347, 4.917244, 4.921369, 
    4.925701, 4.930154, 4.934687, 4.939281, 4.94393, 4.948625, 4.953344, 
    4.958044, 4.959407, 4.968792, 4.97213, 4.974324, 4.975806, 4.976653, 
    4.979882, 4.981626, 4.98219, 4.980597, 4.976579, 4.969752, 4.960011, 
    4.947186, 4.932035, 4.914319, 4.898144, 4.881041, 4.863939, 4.847887, 
    4.833943, 4.823065, 4.816005, 4.813236, 4.814918, 4.820882, 4.830656, 
    4.843504, 4.858468, 4.874428, 4.890163, 4.904439, 4.916101, 4.924196, 
    4.928107,
  // momentumX(18,42, 0-49)
    4.913782, 4.912883, 4.913308, 4.914782, 4.917043, 4.919858, 4.923043, 
    4.926467, 4.93005, 4.933751, 4.937549, 4.941423, 4.945343, 4.949245, 
    4.953024, 4.954234, 4.963964, 4.96634, 4.967675, 4.96837, 4.968452, 
    4.970979, 4.972106, 4.972164, 4.969982, 4.965353, 4.957918, 4.947659, 
    4.934467, 4.919428, 4.902383, 4.887368, 4.871888, 4.856811, 4.843086, 
    4.831631, 4.823244, 4.818518, 4.817794, 4.821123, 4.82827, 4.83873, 
    4.851759, 4.866421, 4.881636, 4.896245, 4.9091, 4.919161, 4.925624, 
    4.928048,
  // momentumX(18,43, 0-49)
    4.919908, 4.918075, 4.917529, 4.918031, 4.919343, 4.921244, 4.923561, 
    4.926164, 4.928969, 4.931925, 4.934999, 4.938159, 4.941349, 4.944471, 
    4.947376, 4.948405, 4.958177, 4.959578, 4.960035, 4.959912, 4.959199, 
    4.960948, 4.961421, 4.960978, 4.958283, 4.953208, 4.945422, 4.934996, 
    4.921866, 4.907401, 4.8915, 4.878047, 4.864542, 4.851766, 4.840542, 
    4.831635, 4.82568, 4.823121, 4.824172, 4.828796, 4.8367, 4.847362, 
    4.860054, 4.873881, 4.887831, 4.900847, 4.911908, 4.920138, 4.924921, 
    4.926015,
  // momentumX(18,44, 0-49)
    4.924776, 4.921913, 4.92034, 4.91985, 4.920226, 4.921264, 4.92279, 
    4.924667, 4.926798, 4.929115, 4.931567, 4.934095, 4.936621, 4.939024, 
    4.941122, 4.941914, 4.951438, 4.951888, 4.951467, 4.95051, 4.94899, 
    4.94992, 4.94973, 4.948813, 4.945714, 4.940386, 4.932531, 4.9223, 
    4.909667, 4.896218, 4.881884, 4.870344, 4.859107, 4.848838, 4.840219, 
    4.833856, 4.830224, 4.829626, 4.832157, 4.837701, 4.845929, 4.856311, 
    4.868156, 4.880635, 4.89284, 4.903851, 4.912822, 4.91908, 4.922236, 
    4.922259,
  // momentumX(18,45, 0-49)
    4.928407, 4.924418, 4.921751, 4.920234, 4.919677, 4.919885, 4.920683, 
    4.921923, 4.923484, 4.925271, 4.927204, 4.929194, 4.931141, 4.932897, 
    4.934264, 4.934757, 4.943786, 4.943328, 4.942047, 4.94026, 4.937941, 
    4.93805, 4.937223, 4.935887, 4.932515, 4.927137, 4.9195, 4.909817, 
    4.898086, 4.886047, 4.873634, 4.864293, 4.855537, 4.847908, 4.841933, 
    4.838057, 4.836599, 4.837729, 4.841436, 4.847537, 4.855672, 4.865327, 
    4.875862, 4.886545, 4.896604, 4.9053, 4.912002, 4.916276, 4.917975, 
    4.917284,
  // momentumX(18,46, 0-49)
    4.931002, 4.925789, 4.921949, 4.919353, 4.917837, 4.917222, 4.917328, 
    4.917989, 4.919061, 4.920411, 4.921917, 4.92346, 4.924904, 4.926087, 
    4.926797, 4.926932, 4.935273, 4.933967, 4.931861, 4.929269, 4.926188, 
    4.925509, 4.924102, 4.922422, 4.918921, 4.9137, 4.906552, 4.897737, 
    4.887263, 4.876956, 4.866735, 4.859797, 4.853657, 4.848723, 4.845367, 
    4.843875, 4.844419, 4.84704, 4.851633, 4.857956, 4.865634, 4.87418, 
    4.883031, 4.891579, 4.899223, 4.905437, 4.90984, 4.912262, 4.912797, 
    4.911825,
  // momentumX(18,47, 0-49)
    4.932955, 4.926421, 4.921322, 4.91757, 4.91504, 4.913567, 4.912973, 
    4.913074, 4.91369, 4.914652, 4.915792, 4.916949, 4.917954, 4.91862, 
    4.918736, 4.91845, 4.925973, 4.923887, 4.921003, 4.917657, 4.913873, 
    4.912481, 4.910572, 4.908642, 4.905159, 4.900286, 4.893863, 4.88618, 
    4.877249, 4.868914, 4.861065, 4.856644, 4.853178, 4.850926, 4.850114, 
    4.850874, 4.853234, 4.85712, 4.862342, 4.86861, 4.875546, 4.88271, 
    4.88963, 4.895852, 4.900975, 4.904717, 4.906961, 4.907805, 4.907571, 
    4.906791,
  // momentumX(18,48, 0-49)
    4.934845, 4.9269, 4.920446, 4.915445, 4.911812, 4.909406, 4.908049, 
    4.907547, 4.907685, 4.908252, 4.909031, 4.909818, 4.910404, 4.910583, 
    4.91014, 4.909373, 4.916004, 4.9132, 4.909599, 4.905562, 4.90116, 
    4.899149, 4.896842, 4.894763, 4.891435, 4.887076, 4.881566, 4.875215, 
    4.868028, 4.861816, 4.856431, 4.854557, 4.85374, 4.854105, 4.855721, 
    4.858578, 4.862577, 4.867533, 4.873183, 4.879201, 4.885219, 4.890858, 
    4.895762, 4.899647, 4.902333, 4.903794, 4.904185, 4.903849, 4.903304, 
    4.90318,
  // momentumX(18,49, 0-49)
    4.943079, 4.933022, 4.92444, 4.917368, 4.911783, 4.907586, 4.904629, 
    4.902708, 4.901586, 4.901, 4.900681, 4.900353, 4.899747, 4.898587, 
    4.896599, 4.894702, 4.907625, 4.902482, 4.896469, 4.890329, 4.884231, 
    4.883526, 4.882961, 4.883486, 4.882074, 4.87913, 4.874318, 4.868094, 
    4.860242, 4.854196, 4.849467, 4.851037, 4.85378, 4.857646, 4.86253, 
    4.868235, 4.874485, 4.880953, 4.887276, 4.893087, 4.898046, 4.901875, 
    4.904406, 4.905601, 4.905601, 4.904716, 4.90344, 4.902396, 4.902278, 
    4.903772,
  // momentumX(19,0, 0-49)
    4.863467, 4.857262, 4.854007, 4.853439, 4.855211, 4.858918, 4.86413, 
    4.870421, 4.877393, 4.884692, 4.892019, 4.899126, 4.905809, 4.911901, 
    4.917256, 4.921696, 4.926414, 4.929109, 4.930936, 4.931877, 4.931879, 
    4.93122, 4.92947, 4.92665, 4.922586, 4.917221, 4.910484, 4.902398, 
    4.893026, 4.882643, 4.871445, 4.860118, 4.848811, 4.838039, 4.828342, 
    4.820229, 4.814119, 4.8103, 4.808887, 4.80981, 4.812818, 4.817494, 
    4.823306, 4.829645, 4.835906, 4.841548, 4.846171, 4.849586, 4.85186, 
    4.853332,
  // momentumX(19,1, 0-49)
    4.865608, 4.859947, 4.857208, 4.857111, 4.8593, 4.863361, 4.868865, 
    4.875392, 4.882556, 4.890017, 4.897492, 4.904748, 4.911586, 4.917842, 
    4.923354, 4.927824, 4.933651, 4.936447, 4.938407, 4.939521, 4.939701, 
    4.939492, 4.938069, 4.935489, 4.931462, 4.925898, 4.918675, 4.909807, 
    4.899339, 4.887649, 4.874897, 4.862156, 4.849326, 4.837008, 4.825834, 
    4.816401, 4.809213, 4.804626, 4.802801, 4.803697, 4.807059, 4.812455, 
    4.8193, 4.826921, 4.834619, 4.841738, 4.847753, 4.85234, 4.855436, 
    4.857277,
  // momentumX(19,2, 0-49)
    4.868079, 4.86294, 4.86067, 4.86098, 4.863502, 4.867823, 4.873523, 
    4.880189, 4.887453, 4.894991, 4.90254, 4.909874, 4.91681, 4.923179, 
    4.928813, 4.933246, 4.940066, 4.942986, 4.945104, 4.946426, 4.946843, 
    4.947165, 4.946175, 4.943969, 4.940157, 4.934615, 4.927167, 4.917808, 
    4.90655, 4.893838, 4.879786, 4.865834, 4.851622, 4.837819, 4.825143, 
    4.814283, 4.805833, 4.800229, 4.7977, 4.798252, 4.801656, 4.807476, 
    4.815114, 4.823852, 4.832918, 4.841565, 4.849153, 4.855217, 4.859553, 
    4.862253,
  // momentumX(19,3, 0-49)
    4.870552, 4.86591, 4.864064, 4.864718, 4.867503, 4.872014, 4.877833, 
    4.884569, 4.891868, 4.899426, 4.906993, 4.914361, 4.921353, 4.927806, 
    4.93355, 4.937875, 4.945512, 4.948591, 4.950888, 4.952444, 4.953139, 
    4.954044, 4.953572, 4.95185, 4.948418, 4.943113, 4.935712, 4.926178, 
    4.914483, 4.901093, 4.886057, 4.871165, 4.855776, 4.840611, 4.826462, 
    4.814105, 4.804229, 4.797366, 4.793829, 4.793693, 4.796775, 4.802673, 
    4.810785, 4.820376, 4.830633, 4.840738, 4.84995, 4.857678, 4.863564, 
    4.867543,
  // momentumX(19,4, 0-49)
    4.872817, 4.868643, 4.867184, 4.868135, 4.871129, 4.875768, 4.881651, 
    4.888405, 4.895691, 4.903227, 4.910775, 4.918141, 4.92516, 4.931677, 
    4.937528, 4.941673, 4.949905, 4.953179, 4.955673, 4.957477, 4.958472, 
    4.959987, 4.960082, 4.958926, 4.956011, 4.951143, 4.944056, 4.934675, 
    4.922916, 4.909231, 4.893579, 4.878071, 4.861773, 4.845433, 4.829899, 
    4.816028, 4.804605, 4.796266, 4.79143, 4.790257, 4.792642, 4.798227, 
    4.806442, 4.816557, 4.827739, 4.839124, 4.849892, 4.859341, 4.866971, 
    4.872547,
  // momentumX(19,5, 0-49)
    4.874774, 4.871048, 4.869942, 4.871148, 4.874307, 4.879029, 4.884934, 
    4.891664, 4.898901, 4.906378, 4.913873, 4.921207, 4.928225, 4.93479, 
    4.940752, 4.944649, 4.953211, 4.956712, 4.959419, 4.961472, 4.962777, 
    4.964893, 4.965576, 4.96503, 4.962738, 4.958478, 4.951951, 4.943034, 
    4.931594, 4.918012, 4.902144, 4.886379, 4.869491, 4.852226, 4.835463, 
    4.820125, 4.807089, 4.797104, 4.790708, 4.788169, 4.789482, 4.79436, 
    4.802285, 4.812552, 4.824332, 4.836738, 4.848891, 4.860003, 4.869445, 
    4.876825,
  // momentumX(19,6, 0-49)
    4.876401, 4.873109, 4.872334, 4.873767, 4.877055, 4.881827, 4.887718, 
    4.894387, 4.901539, 4.90892, 4.916327, 4.923593, 4.930583, 4.937176, 
    4.943255, 4.946844, 4.955447, 4.959205, 4.962132, 4.964428, 4.966038, 
    4.968722, 4.969982, 4.970057, 4.968456, 4.964935, 4.959171, 4.951004, 
    4.94024, 4.92715, 4.911473, 4.895832, 4.878706, 4.860817, 4.843043, 
    4.826352, 4.811706, 4.799966, 4.7918, 4.78761, 4.787505, 4.791297, 
    4.798542, 4.808578, 4.820599, 4.833713, 4.847009, 4.85963, 4.870845, 
    4.880115,
  // momentumX(19,7, 0-49)
    4.877742, 4.87488, 4.87442, 4.876059, 4.879453, 4.884243, 4.890086, 
    4.896661, 4.903688, 4.910936, 4.918213, 4.925372, 4.932297, 4.938896, 
    4.945095, 4.948344, 4.956688, 4.960714, 4.963864, 4.966398, 4.968299, 
    4.971492, 4.973291, 4.973963, 4.973082, 4.970386, 4.965547, 4.958364, 
    4.94859, 4.936349, 4.921254, 4.906102, 4.889108, 4.870925, 4.852411, 
    4.83455, 4.818367, 4.804838, 4.79476, 4.78869, 4.78687, 4.789238, 
    4.795435, 4.80487, 4.816771, 4.830261, 4.844414, 4.858326, 4.871181, 
    4.882321,
  // momentumX(19,8, 0-49)
    4.878867, 4.876438, 4.876289, 4.878121, 4.881602, 4.886387, 4.892151, 
    4.898596, 4.90546, 4.912529, 4.919632, 4.926641, 4.93346, 4.940037, 
    4.946343, 4.94926, 4.957064, 4.961346, 4.964719, 4.967476, 4.969651, 
    4.973279, 4.975556, 4.976775, 4.976603, 4.974774, 4.970967, 4.964946, 
    4.956418, 4.94533, 4.931167, 4.916834, 4.900319, 4.88219, 4.863243, 
    4.844447, 4.826875, 4.811594, 4.799544, 4.791435, 4.787673, 4.788329, 
    4.793161, 4.801657, 4.813101, 4.826638, 4.841345, 4.856289, 4.87059, 
    4.883487,
  // momentumX(19,9, 0-49)
    4.879853, 4.877869, 4.878036, 4.880059, 4.883614, 4.888375, 4.894034, 
    4.900314, 4.906975, 4.913821, 4.920701, 4.927508, 4.934181, 4.940696, 
    4.94708, 4.94973, 4.956745, 4.961252, 4.964836, 4.967809, 4.970237, 
    4.974212, 4.976891, 4.978584, 4.979081, 4.978118, 4.975397, 4.970651, 
    4.963554, 4.953855, 4.940918, 4.927673, 4.911951, 4.894206, 4.875144, 
    4.855691, 4.836935, 4.820017, 4.80601, 4.795788, 4.789926, 4.788655, 
    4.791863, 4.799135, 4.809819, 4.823099, 4.838062, 4.853761, 4.86927, 
    4.883741,
  // momentumX(19,10, 0-49)
    4.880766, 4.879248, 4.879743, 4.881961, 4.885587, 4.890312, 4.895844, 
    4.901929, 4.90835, 4.91493, 4.921543, 4.928103, 4.934577, 4.940979, 
    4.947385, 4.949909, 4.955944, 4.960614, 4.964392, 4.967567, 4.970238, 
    4.974462, 4.977457, 4.979537, 4.980639, 4.980505, 4.978874, 4.975456, 
    4.969903, 4.961752, 4.950266, 4.938305, 4.923625, 4.906556, 4.887687, 
    4.867873, 4.848182, 4.829807, 4.813938, 4.801608, 4.79357, 4.79023, 
    4.79162, 4.797441, 4.807114, 4.819869, 4.834813, 4.850992, 4.867447, 
    4.883266,
  // momentumX(19,11, 0-49)
    4.881644, 4.880621, 4.881466, 4.883892, 4.887596, 4.892278, 4.897672, 
    4.903541, 4.909692, 4.91597, 4.922273, 4.92854, 4.934764, 4.94099, 
    4.94733, 4.949949, 4.954883, 4.959633, 4.963575, 4.966947, 4.969853, 
    4.974226, 4.977445, 4.979825, 4.981448, 4.982079, 4.9815, 4.979406, 
    4.975439, 4.968922, 4.95904, 4.948476, 4.935015, 4.918853, 4.900454, 
    4.880566, 4.860214, 4.840611, 4.823038, 4.80868, 4.798471, 4.792996, 
    4.792449, 4.796651, 4.805115, 4.817122, 4.8318, 4.8482, 4.865337, 4.882246,
  // momentumX(19,12, 0-49)
    4.882496, 4.881999, 4.883224, 4.885882, 4.889676, 4.894325, 4.899577, 
    4.90522, 4.911082, 4.917034, 4.922996, 4.928931, 4.934853, 4.940827, 
    4.946981, 4.949989, 4.95378, 4.958515, 4.962585, 4.966149, 4.969291, 
    4.973717, 4.977075, 4.979658, 4.981715, 4.983027, 4.983429, 4.982606, 
    4.9802, 4.975337, 4.967144, 4.958006, 4.945863, 4.930773, 4.913065, 
    4.893366, 4.872625, 4.852049, 4.832983, 4.816743, 4.804437, 4.796834, 
    4.794295, 4.796777, 4.803885, 4.814964, 4.829169, 4.845552, 4.863111, 
    4.880845,
  // momentumX(19,13, 0-49)
    4.883292, 4.883357, 4.884997, 4.887918, 4.891829, 4.896464, 4.901587, 
    4.907006, 4.912575, 4.918189, 4.923789, 4.929358, 4.934927, 4.940565, 
    4.94639, 4.950139, 4.952823, 4.957446, 4.961614, 4.96537, 4.968758, 
    4.973145, 4.976562, 4.979265, 4.981663, 4.983564, 4.98485, 4.985204, 
    4.984283, 4.981029, 4.974552, 4.966794, 4.955986, 4.942058, 4.9252, 
    4.905908, 4.885034, 4.863748, 4.84343, 4.825501, 4.811233, 4.801569, 
    4.797047, 4.797762, 4.803423, 4.813437, 4.826993, 4.84315, 4.86089, 
    4.879182,
  // momentumX(19,14, 0-49)
    4.883975, 4.884635, 4.886726, 4.889947, 4.894012, 4.898662, 4.903681, 
    4.908897, 4.914186, 4.919464, 4.924696, 4.929881, 4.935049, 4.940267, 
    4.945613, 4.950459, 4.952142, 4.956577, 4.960824, 4.964785, 4.968439, 
    4.972709, 4.976121, 4.978877, 4.981533, 4.983922, 4.985978, 4.987384, 
    4.98782, 4.986081, 4.981294, 4.974806, 4.965281, 4.952532, 4.936615, 
    4.917893, 4.897106, 4.875359, 4.85404, 4.83465, 4.818594, 4.806993, 
    4.800546, 4.799497, 4.803661, 4.812512, 4.825278, 4.841026, 4.858731, 
    4.877334,
  // momentumX(19,15, 0-49)
    4.884464, 4.885746, 4.888322, 4.891884, 4.896142, 4.900849, 4.905801, 
    4.910846, 4.915881, 4.920848, 4.925724, 4.930517, 4.93526, 4.939989, 
    4.94473, 4.95096, 4.951797, 4.956015, 4.960347, 4.964542, 4.968503, 
    4.972597, 4.97596, 4.978716, 4.981555, 4.984333, 4.987031, 4.989339, 
    4.990971, 4.990606, 4.987436, 4.98206, 4.973706, 4.962089, 4.94714, 
    4.929091, 4.908561, 4.886575, 4.864501, 4.843886, 4.82625, 4.812865, 
    4.804594, 4.801823, 4.804478, 4.812106, 4.823973, 4.83916, 4.856639, 
    4.875334,
  // momentumX(19,16, 0-49)
    4.884663, 4.88658, 4.889668, 4.893605, 4.898099, 4.902907, 4.907837, 
    4.912756, 4.917584, 4.922279, 4.926834, 4.931263, 4.935582, 4.939795, 
    4.943863, 4.951606, 4.951766, 4.955799, 4.960267, 4.964756, 4.969089, 
    4.972967, 4.976264, 4.978997, 4.981962, 4.985034, 4.988237, 4.991272, 
    4.993902, 4.994734, 4.993072, 4.988607, 4.981264, 4.970675, 4.956662, 
    4.93933, 4.919178, 4.897139, 4.874533, 4.85293, 4.833932, 4.818943, 
    4.808976, 4.804556, 4.805722, 4.812094, 4.822984, 4.837489, 4.854583, 
    4.873177,
  // momentumX(19,17, 0-49)
    4.884471, 4.887014, 4.890623, 4.894957, 4.899719, 4.904669, 4.909626, 
    4.914478, 4.919161, 4.923654, 4.92796, 4.932091, 4.936043, 4.939777, 
    4.943196, 4.952326, 4.951941, 4.9559, 4.960605, 4.965496, 4.970294, 
    4.973958, 4.977208, 4.979924, 4.982979, 4.986258, 4.989816, 4.993383, 
    4.996779, 4.998592, 4.998283, 4.994504, 4.987976, 4.978271, 4.96511, 
    4.948489, 4.928789, 4.90684, 4.883897, 4.861527, 4.841388, 4.824988, 
    4.813472, 4.8075, 4.807219, 4.81233, 4.822189, 4.835921, 4.852504, 
    4.870842,
  // momentumX(19,18, 0-49)
    4.883793, 4.886919, 4.891025, 4.895751, 4.900793, 4.905913, 4.910947, 
    4.915798, 4.920425, 4.924825, 4.929009, 4.932978, 4.936702, 4.940094, 
    4.94299, 4.953041, 4.952164, 4.956231, 4.961337, 4.966779, 4.972184, 
    4.975669, 4.978938, 4.981686, 4.984823, 4.988232, 4.991991, 4.995869, 
    4.999767, 5.002297, 5.003136, 4.999793, 4.993859, 4.984858, 4.972429, 
    4.956472, 4.937254, 4.915499, 4.892387, 4.869453, 4.848384, 4.830771, 
    4.817868, 4.810457, 4.808792, 4.812659, 4.821465, 4.834362, 4.850341, 
    4.868311,
  // momentumX(19,19, 0-49)
    4.882538, 4.886151, 4.890681, 4.895749, 4.901048, 4.906345, 4.911496, 
    4.916429, 4.921131, 4.92561, 4.929882, 4.933926, 4.937669, 4.94096, 
    4.943571, 4.95371, 4.952253, 4.956655, 4.962374, 4.968572, 4.974777, 
    4.978183, 4.981593, 4.984472, 4.987724, 4.991202, 4.994999, 4.998935, 
    5.003021, 5.00595, 5.007671, 5.004481, 4.998894, 4.990393, 4.978553, 
    4.963183, 4.944447, 4.922963, 4.899824, 4.876513, 4.854719, 4.836087, 
    4.821965, 4.813243, 4.810278, 4.812939, 4.820692, 4.832723, 4.848042, 
    4.865566,
  // momentumX(19,20, 0-49)
    4.881588, 4.886601, 4.892593, 4.899169, 4.905969, 4.912692, 4.919097, 
    4.924998, 4.930258, 4.934787, 4.938541, 4.941516, 4.943758, 4.94535, 
    4.946416, 0, 4.960864, 4.963375, 4.966852, 4.970822, 4.975077, 4.975944, 
    4.977604, 4.979422, 4.982367, 4.986216, 4.99093, 4.996161, 5.00179, 
    5.006393, 5.010077, 5.007852, 5.003162, 4.995485, 4.98438, 4.969624, 
    4.951338, 4.930086, 4.906902, 4.883231, 4.860764, 4.841182, 4.825912, 
    4.815937, 4.811708, 4.813176, 4.819865, 4.831002, 4.845614, 4.862631,
  // momentumX(19,21, 0-49)
    4.87942, 4.884988, 4.891505, 4.898539, 4.905715, 4.912723, 4.919326, 
    4.92536, 4.930717, 4.935334, 4.939191, 4.942301, 4.944708, 4.946493, 
    4.947779, 0, 4.960035, 4.963074, 4.967126, 4.971672, 4.976431, 4.976584, 
    4.977723, 4.979072, 4.98174, 4.985524, 4.990396, 4.995993, 5.002195, 
    5.007564, 5.012428, 5.010612, 5.006535, 4.999634, 4.989399, 4.975526, 
    4.958041, 4.937399, 4.914538, 4.890834, 4.867946, 4.84758, 4.831234, 
    4.819987, 4.814397, 4.814506, 4.819916, 4.829904, 4.843533, 4.859751,
  // momentumX(19,22, 0-49)
    4.876799, 4.882879, 4.889917, 4.897455, 4.905089, 4.912499, 4.919439, 
    4.925747, 4.931327, 4.936132, 4.940154, 4.943415, 4.945968, 4.947898, 
    4.949335, 0, 4.959913, 4.963387, 4.967949, 4.973043, 4.978314, 4.977839, 
    4.978555, 4.979537, 4.982003, 4.985746, 4.990732, 4.996574, 5.003149, 
    5.009007, 5.014683, 5.012933, 5.009101, 5.002608, 4.992905, 4.97964, 
    4.962763, 4.942643, 4.920128, 4.896511, 4.873403, 4.852501, 4.835343, 
    4.823078, 4.816355, 4.815298, 4.819583, 4.828539, 4.841269, 4.856745,
  // momentumX(19,23, 0-49)
    4.873835, 4.880381, 4.887924, 4.895979, 4.904121, 4.912008, 4.91938, 
    4.926068, 4.931972, 4.937049, 4.941298, 4.944747, 4.947457, 4.949518, 
    4.951072, 0, 4.960715, 4.964478, 4.969381, 4.974841, 4.980453, 4.979389, 
    4.979692, 4.980315, 4.982558, 4.986212, 4.991232, 4.997212, 5.004019, 
    5.010185, 5.016409, 5.014583, 5.010819, 5.004539, 4.995176, 4.982343, 
    4.96594, 4.946269, 4.924097, 4.900642, 4.877457, 4.856218, 4.838474, 
    4.825424, 4.817783, 4.815747, 4.819055, 4.827091, 4.838994, 4.853765,
  // momentumX(19,24, 0-49)
    4.870672, 4.877634, 4.885653, 4.894224, 4.902894, 4.911297, 4.91916, 
    4.926295, 4.932595, 4.93801, 4.94254, 4.946218, 4.949106, 4.951304, 
    4.952971, 0, 4.962595, 4.966502, 4.971569, 4.977206, 4.982986, 4.981498, 
    4.981503, 4.981868, 4.98394, 4.987504, 4.992511, 4.998539, 5.005456, 
    5.011777, 5.018311, 5.016373, 5.012581, 5.006359, 4.997128, 4.984486, 
    4.968306, 4.948847, 4.926829, 4.903417, 4.880123, 4.858602, 4.840403, 
    4.826757, 4.818415, 4.815626, 4.818173, 4.82548, 4.836718, 4.850913,
  // momentumX(19,25, 0-49)
    4.867481, 4.874813, 4.883271, 4.892335, 4.901527, 4.91046, 4.918839, 
    4.926459, 4.933195, 4.938988, 4.943835, 4.947769, 4.950856, 4.953206, 
    4.954986, 0, 4.965112, 4.969028, 4.974089, 4.979712, 4.985476, 4.983797, 
    4.983668, 4.983923, 4.985918, 4.989429, 4.994407, 5.000427, 5.007351, 
    5.013689, 5.020282, 5.018254, 5.014394, 5.008122, 4.998861, 4.986204, 
    4.970013, 4.950536, 4.92847, 4.904962, 4.881504, 4.859735, 4.841204, 
    4.827145, 4.818328, 4.815025, 4.817045, 4.823834, 4.834585, 4.848341,
  // momentumX(19,26, 0-49)
    4.864459, 4.87211, 4.880964, 4.890482, 4.900172, 4.909622, 4.918519, 
    4.926631, 4.933817, 4.940006, 4.945184, 4.949382, 4.952669, 4.955164, 
    4.957052, 0, 4.968115, 4.971904, 4.97679, 4.98221, 4.987775, 4.986162, 
    4.986086, 4.986403, 4.988436, 4.991954, 4.996908, 5.002874, 5.009715, 
    5.015938, 5.022344, 5.020271, 5.016323, 5.009913, 5.00047, 4.98759, 
    4.971152, 4.951414, 4.929086, 4.905328, 4.881636, 4.859649, 4.840906, 
    4.826628, 4.817581, 4.814027, 4.815778, 4.822286, 4.832751, 4.846226,
  // momentumX(19,27, 0-49)
    4.861812, 4.869731, 4.878926, 4.888848, 4.898993, 4.908931, 4.918322, 
    4.926916, 4.934547, 4.941125, 4.946622, 4.951062, 4.954522, 4.957128, 
    4.959073, 0, 4.97163, 4.975142, 4.979673, 4.984694, 4.989872, 4.988544, 
    4.988675, 4.989195, 4.991359, 4.994929, 4.999852, 5.005712, 5.012372, 
    5.018343, 5.024315, 5.022226, 5.018149, 5.011499, 5.001717, 4.988418, 
    4.971513, 4.951303, 4.928545, 4.904437, 4.880499, 4.858378, 4.839594, 
    4.825338, 4.816338, 4.812825, 4.814583, 4.821054, 4.831435, 4.844779,
  // momentumX(19,28, 0-49)
    4.859741, 4.867873, 4.877347, 4.887616, 4.898163, 4.908547, 4.918406, 
    4.927459, 4.935514, 4.942453, 4.948228, 4.952856, 4.956412, 4.959038, 
    4.960937, 0, 4.975993, 4.979054, 4.983034, 4.987453, 4.992063, 4.991148, 
    4.991572, 4.99238, 4.994724, 4.998356, 5.003215, 5.008902, 5.015275, 
    5.020853, 5.026161, 5.024028, 5.019733, 5.012695, 5.002378, 4.988438, 
    4.970845, 4.949972, 4.926649, 4.90214, 4.87801, 4.8559, 4.837305, 
    4.823361, 4.814726, 4.811572, 4.813638, 4.820332, 4.830835, 4.844201,
  // momentumX(19,29, 0-49)
    4.858432, 4.866712, 4.876399, 4.88695, 4.897851, 4.908648, 4.918948, 
    4.92844, 4.936892, 4.944144, 4.950123, 4.95483, 4.958349, 4.960835, 
    4.962511, 0, 4.980938, 4.983357, 4.986584, 4.990198, 4.994048, 4.993536, 
    4.994227, 4.995311, 4.997817, 5.001482, 5.006229, 5.011665, 5.017635, 
    5.022667, 5.027061, 5.024763, 5.020088, 5.012481, 5.00145, 4.986721, 
    4.968343, 4.946784, 4.922968, 4.898229, 4.874156, 4.852381, 4.834337, 
    4.821075, 4.813166, 4.810695, 4.81334, 4.820467, 4.831241, 4.8447,
  // momentumX(19,30, 0-49)
    4.857325, 4.864811, 4.87362, 4.883223, 4.89315, 4.903017, 4.912543, 
    4.921545, 4.929926, 4.937651, 4.944711, 4.951098, 4.956753, 4.961548, 
    4.965257, 4.981699, 4.974598, 4.979191, 4.985151, 4.991585, 4.998013, 
    5.000706, 5.003804, 5.006528, 5.009774, 5.013294, 5.017124, 5.021049, 
    5.02509, 5.027961, 5.029866, 5.026049, 5.019855, 5.010766, 4.998342, 
    4.982376, 4.962988, 4.940724, 4.916574, 4.891904, 4.868294, 4.847318, 
    4.830311, 4.818207, 4.811459, 4.810057, 4.813608, 4.821434, 4.832671, 
    4.846352,
  // momentumX(19,31, 0-49)
    4.858174, 4.865802, 4.874738, 4.884463, 4.894507, 4.904485, 4.9141, 
    4.923157, 4.931543, 4.939215, 4.946176, 4.952444, 4.958014, 4.962843, 
    4.966795, 4.981744, 4.976817, 4.98103, 4.986337, 4.99197, 4.997562, 
    5.000377, 5.003357, 5.005968, 5.009114, 5.01259, 5.016417, 5.020319, 
    5.02421, 5.026711, 5.027736, 5.023791, 5.017277, 5.007711, 4.994723, 
    4.978187, 4.958328, 4.935792, 4.911653, 4.88733, 4.8644, 4.844378, 
    4.828509, 4.817608, 4.812016, 4.811631, 4.815988, 4.824363, 4.835867, 
    4.849523,
  // momentumX(19,32, 0-49)
    4.860078, 4.867659, 4.876506, 4.886116, 4.896039, 4.905897, 4.915404, 
    4.924363, 4.932662, 4.940258, 4.947163, 4.953413, 4.959052, 4.964091, 
    4.968487, 4.981169, 4.978074, 4.982155, 4.987026, 4.992065, 4.997014, 
    5.000091, 5.003103, 5.005722, 5.008819, 5.012202, 5.015869, 5.019507, 
    5.02294, 5.024753, 5.024618, 5.020299, 5.013247, 5.003031, 4.989363, 
    4.972216, 4.95193, 4.929254, 4.905345, 4.881649, 4.859718, 4.840992, 
    4.826592, 4.817206, 4.813052, 4.813928, 4.819293, 4.828377, 4.840262, 
    4.853956,
  // momentumX(19,33, 0-49)
    4.863094, 4.870475, 4.879053, 4.888352, 4.897948, 4.907487, 4.916703, 
    4.925407, 4.9335, 4.940943, 4.947758, 4.953999, 4.959738, 4.965044, 
    4.969951, 4.980079, 4.97859, 4.982728, 4.987326, 4.991925, 4.996374, 
    4.999796, 5.002942, 5.005651, 5.008716, 5.011941, 5.015303, 5.018456, 
    5.021159, 5.022017, 5.020511, 5.015593, 5.007808, 4.996795, 4.982359, 
    4.964593, 4.943953, 4.921297, 4.897847, 4.875063, 4.854445, 4.837331, 
    4.824705, 4.817112, 4.814642, 4.816987, 4.823531, 4.833456, 4.845809, 
    4.859584,
  // momentumX(19,34, 0-49)
    4.867206, 4.874252, 4.882409, 4.891233, 4.900333, 4.909385, 4.918148, 
    4.926455, 4.934219, 4.941414, 4.948065, 4.954243, 4.960041, 4.96557, 
    4.970939, 4.978593, 4.978584, 4.98288, 4.987299, 4.991557, 4.995606, 
    4.999401, 5.002732, 5.005574, 5.008594, 5.011591, 5.014505, 5.016977, 
    5.018713, 5.018397, 5.015368, 5.009659, 5.000988, 4.989071, 4.973829, 
    4.955482, 4.934607, 4.912163, 4.889425, 4.867839, 4.848833, 4.833615, 
    4.823024, 4.817452, 4.816856, 4.820828, 4.828676, 4.839528, 4.852401, 
    4.86627,
  // momentumX(19,35, 0-49)
    4.872328, 4.878919, 4.886526, 4.89474, 4.903203, 4.911632, 4.919809, 
    4.927599, 4.934926, 4.941772, 4.948174, 4.954204, 4.959976, 4.965626, 
    4.971318, 4.976828, 4.978239, 4.982703, 4.986978, 4.990948, 4.99466, 
    4.998809, 5.002337, 5.005319, 5.008259, 5.010948, 5.01328, 5.014896, 
    5.015461, 5.013795, 5.009148, 5.002493, 4.992821, 4.979948, 4.963921, 
    4.945088, 4.92415, 4.90215, 4.880391, 4.860284, 4.843158, 4.83008, 
    4.821725, 4.818338, 4.819746, 4.825438, 4.834654, 4.84647, 4.859871, 
    4.873812,
  // momentumX(19,36, 0-49)
    4.878319, 4.884347, 4.891294, 4.898786, 4.906506, 4.914204, 4.921698, 
    4.928871, 4.935667, 4.942079, 4.948146, 4.953941, 4.95958, 4.965217, 
    4.97104, 4.974863, 4.977667, 4.982239, 4.986354, 4.99006, 4.993469, 
    4.997919, 5.001616, 5.004714, 5.007523, 5.009817, 5.011443, 5.012049, 
    5.011275, 5.008129, 5.00182, 4.994109, 4.98338, 4.969563, 4.952835, 
    4.933675, 4.912894, 4.891598, 4.871095, 4.852732, 4.837718, 4.826962, 
    4.820982, 4.819872, 4.823338, 4.830776, 4.841359, 4.854115, 4.868001, 
    4.881951,
  // momentumX(19,37, 0-49)
    4.884991, 4.890361, 4.896557, 4.903244, 4.910141, 4.917033, 4.923767, 
    4.930253, 4.936448, 4.942355, 4.948011, 4.953487, 4.958893, 4.964376, 
    4.97013, 4.972736, 4.976905, 4.981477, 4.985387, 4.988821, 4.991942, 
    4.996607, 5.000417, 5.003583, 5.006192, 5.008002, 5.008813, 5.008285, 
    5.006043, 5.001339, 4.993384, 4.98456, 4.972786, 4.958107, 4.940834, 
    4.921567, 4.901206, 4.880898, 4.861922, 4.845537, 4.832814, 4.824502, 
    4.820959, 4.822139, 4.827637, 4.836768, 4.848647, 4.862257, 4.876529, 
    4.890384,
  // momentumX(19,38, 0-49)
    4.892121, 4.896754, 4.902132, 4.907953, 4.913973, 4.920011, 4.92594, 
    4.931687, 4.937231, 4.942576, 4.947761, 4.952847, 4.957928, 4.963131, 
    4.968633, 4.970451, 4.975925, 4.980362, 4.984005, 4.987148, 4.989974, 
    4.994747, 4.99859, 5.001753, 5.004083, 5.005324, 5.005226, 5.003472, 
    4.999688, 4.993407, 4.983876, 4.973956, 4.96122, 4.945838, 4.928244, 
    4.909145, 4.889503, 4.870472, 4.853275, 4.839058, 4.828744, 4.82292, 
    4.821793, 4.825191, 4.832617, 4.843311, 4.856339, 4.870652, 4.885157, 
    4.898771,
  // momentumX(19,39, 0-49)
    4.899467, 4.903297, 4.907806, 4.912726, 4.917843, 4.923001, 4.928099, 
    4.933086, 4.937946, 4.942693, 4.947358, 4.951997, 4.95668, 4.961504, 
    4.966603, 4.967971, 4.974646, 4.978811, 4.982118, 4.984936, 4.987445, 
    4.992202, 4.995981, 4.999056, 5.00102, 5.001617, 5.000542, 4.997513, 
    4.99217, 4.984358, 4.973391, 4.962465, 4.948932, 4.93308, 4.915452, 
    4.896836, 4.878227, 4.860754, 4.845551, 4.833638, 4.825777, 4.822405, 
    4.823591, 4.829056, 4.838219, 4.850267, 4.864228, 4.879025, 4.893557, 
    4.906746,
  // momentumX(19,40, 0-49)
    4.906766, 4.909746, 4.913357, 4.917359, 4.921566, 4.925843, 4.930111, 
    4.934331, 4.938495, 4.942622, 4.94674, 4.950891, 4.95512, 4.959492, 
    4.964085, 4.965239, 4.97296, 4.976724, 4.979627, 4.98208, 4.984232, 
    4.988842, 4.992447, 4.995337, 4.996855, 4.996744, 4.994654, 4.990354, 
    4.983506, 4.974283, 4.962084, 4.950325, 4.936236, 4.920212, 4.902885, 
    4.885092, 4.867829, 4.852161, 4.839121, 4.829577, 4.824143, 4.823107, 
    4.82642, 4.833713, 4.844347, 4.857467, 4.872072, 4.887079, 4.901387, 
    4.913939,
  // momentumX(19,41, 0-49)
    4.913755, 4.915848, 4.918544, 4.921631, 4.924941, 4.928359, 4.931815, 
    4.935283, 4.938761, 4.942267, 4.945827, 4.949466, 4.953209, 4.957081, 
    4.961106, 4.962186, 4.970744, 4.974006, 4.976444, 4.97848, 4.980226, 
    4.984553, 4.987868, 4.990473, 4.991469, 4.990608, 4.987513, 4.982002, 
    4.973772, 4.963334, 4.950175, 4.93783, 4.923496, 4.90765, 4.890987, 
    4.874359, 4.858728, 4.845076, 4.8343, 4.827125, 4.824011, 4.825119, 
    4.830297, 4.839108, 4.850871, 4.864708, 4.879611, 4.894502, 4.908296, 
    4.919983,
  // momentumX(19,42, 0-49)
    4.92017, 4.921348, 4.923127, 4.925314, 4.927758, 4.930353, 4.933038, 
    4.935792, 4.938614, 4.94152, 4.944527, 4.94765, 4.950894, 4.954247, 
    4.957675, 4.958741, 4.967895, 4.970575, 4.972492, 4.974058, 4.975332, 
    4.979243, 4.982157, 4.984379, 4.984793, 4.983174, 4.979122, 4.97252, 
    4.963109, 4.951718, 4.937935, 4.92532, 4.911098, 4.895811, 4.880182, 
    4.865045, 4.851295, 4.839802, 4.83133, 4.826448, 4.825478, 4.828466, 
    4.835182, 4.845138, 4.857627, 4.871772, 4.886574, 4.900981, 4.913953, 
    4.924549,
  // momentumX(19,43, 0-49)
    4.925763, 4.926003, 4.926868, 4.928182, 4.929801, 4.931626, 4.933599, 
    4.935696, 4.937914, 4.94026, 4.942748, 4.945375, 4.948125, 4.950956, 
    4.953793, 4.954841, 4.96433, 4.966375, 4.967723, 4.968758, 4.969495, 
    4.972867, 4.975272, 4.977025, 4.97682, 4.974465, 4.969556, 4.962043, 
    4.951717, 4.939699, 4.925668, 4.913147, 4.899427, 4.885087, 4.87084, 
    4.857475, 4.845798, 4.836551, 4.830351, 4.827622, 4.828561, 4.833115, 
    4.840987, 4.851663, 4.86443, 4.878427, 4.892694, 4.906231, 4.91807, 
    4.927366,
  // momentumX(19,44, 0-49)
    4.930317, 4.929597, 4.929554, 4.930022, 4.930867, 4.931989, 4.933323, 
    4.934839, 4.936524, 4.938376, 4.940395, 4.942565, 4.944849, 4.94718, 
    4.949445, 4.950438, 4.960001, 4.961379, 4.962115, 4.96256, 4.962694, 
    4.965418, 4.967226, 4.968439, 4.967605, 4.964572, 4.95895, 4.950758, 
    4.93984, 4.927562, 4.913687, 4.901648, 4.888824, 4.875793, 4.863242, 
    4.85188, 4.842403, 4.835417, 4.831395, 4.830625, 4.833188, 4.838951, 
    4.847569, 4.85851, 4.87108, 4.884458, 4.897746, 4.910027, 4.920442, 
    4.928277,
  // momentumX(19,45, 0-49)
    4.933671, 4.931966, 4.931014, 4.930665, 4.930786, 4.931273, 4.932052, 
    4.933077, 4.934319, 4.935762, 4.937385, 4.939156, 4.941019, 4.942884, 
    4.944615, 4.945492, 4.954885, 4.955587, 4.955676, 4.955476, 4.954947, 
    4.956939, 4.958081, 4.958708, 4.957262, 4.953647, 4.947495, 4.938894, 
    4.92774, 4.915594, 4.902283, 4.89111, 4.879552, 4.868159, 4.857555, 
    4.848358, 4.841139, 4.836369, 4.834379, 4.835332, 4.839209, 4.845804, 
    4.854742, 4.86549, 4.877389, 4.889682, 4.901563, 4.912237, 4.920988, 
    4.927265,
  // momentumX(19,46, 0-49)
    4.935753, 4.933025, 4.931156, 4.930007, 4.929449, 4.929368, 4.929675, 
    4.930304, 4.931202, 4.932328, 4.933641, 4.935088, 4.936592, 4.938042, 
    4.939281, 4.939974, 4.948993, 4.949016, 4.948432, 4.947545, 4.946309, 
    4.947513, 4.947949, 4.947968, 4.945961, 4.941886, 4.935413, 4.926697, 
    4.915676, 4.904049, 4.89169, 4.881741, 4.871771, 4.862283, 4.853815, 
    4.846878, 4.841915, 4.83926, 4.839114, 4.841527, 4.846392, 4.853445, 
    4.862292, 4.872415, 4.883203, 4.893989, 4.904093, 4.912873, 4.919795, 
    4.924508,
  // momentumX(19,47, 0-49)
    4.936611, 4.932811, 4.929999, 4.92805, 4.926839, 4.926242, 4.92615, 
    4.92647, 4.927119, 4.928027, 4.929121, 4.930323, 4.931534, 4.932622, 
    4.93342, 4.933862, 4.942347, 4.941703, 4.94043, 4.938825, 4.936858, 
    4.937251, 4.936972, 4.936396, 4.933905, 4.929514, 4.922946, 4.914406, 
    4.903878, 4.893131, 4.882066, 4.873648, 4.86553, 4.858142, 4.851929, 
    4.847281, 4.844512, 4.843832, 4.84532, 4.848924, 4.854459, 4.861622, 
    4.870004, 4.879118, 4.888425, 4.897368, 4.905418, 4.912122, 4.917159, 
    4.920394,
  // momentumX(19,48, 0-49)
    4.936437, 4.931505, 4.927708, 4.924939, 4.923077, 4.921989, 4.921544, 
    4.921619, 4.922096, 4.922868, 4.923826, 4.924857, 4.925838, 4.926618, 
    4.92702, 4.927145, 4.934983, 4.93369, 4.931725, 4.929393, 4.926692, 
    4.926288, 4.925319, 4.924188, 4.921313, 4.916768, 4.910326, 4.90224, 
    4.892526, 4.88297, 4.87348, 4.866836, 4.860761, 4.855598, 4.851686, 
    4.849298, 4.848623, 4.849751, 4.852652, 4.857186, 4.863106, 4.870075, 
    4.877688, 4.885501, 4.89306, 4.89994, 4.905788, 4.910366, 4.913583, 
    4.915535,
  // momentumX(19,49, 0-49)
    4.939479, 4.932686, 4.927199, 4.922946, 4.919828, 4.917706, 4.916431, 
    4.915837, 4.915757, 4.916022, 4.916465, 4.916909, 4.91717, 4.917032, 
    4.916247, 4.915366, 4.929752, 4.926197, 4.921779, 4.917198, 4.912539, 
    4.913105, 4.913378, 4.914213, 4.912521, 4.90855, 4.901885, 4.89297, 
    4.881677, 4.871408, 4.861761, 4.857852, 4.85482, 4.852896, 4.852281, 
    4.853092, 4.855345, 4.858965, 4.86378, 4.869527, 4.875886, 4.882484, 
    4.888945, 4.894903, 4.900057, 4.904189, 4.907223, 4.909227, 4.910436, 
    4.91124,
  // momentumX(20,0, 0-49)
    4.860252, 4.86001, 4.861908, 4.865577, 4.870636, 4.876714, 4.883478, 
    4.890644, 4.897981, 4.905314, 4.912512, 4.919477, 4.926129, 4.932405, 
    4.938227, 4.943402, 4.949084, 4.953224, 4.956752, 4.959602, 4.961658, 
    4.963098, 4.963417, 4.962541, 4.960215, 4.956271, 4.950531, 4.9429, 
    4.933327, 4.921966, 4.908915, 4.894793, 4.879703, 4.864185, 4.848875, 
    4.834458, 4.821619, 4.810974, 4.803027, 4.798102, 4.796328, 4.797613, 
    4.801653, 4.80796, 4.815895, 4.82473, 4.833702, 4.842091, 4.849298, 
    4.854918,
  // momentumX(20,1, 0-49)
    4.862436, 4.862621, 4.86489, 4.86887, 4.874181, 4.880456, 4.887374, 
    4.894657, 4.902087, 4.909499, 4.91677, 4.923805, 4.93053, 4.936876, 
    4.94276, 4.947818, 4.954359, 4.958505, 4.962062, 4.965001, 4.967188, 
    4.969077, 4.969801, 4.969337, 4.967341, 4.963618, 4.957946, 4.950209, 
    4.94033, 4.92852, 4.914805, 4.900119, 4.884272, 4.867824, 4.851451, 
    4.835898, 4.821912, 4.810189, 4.8013, 4.795636, 4.793375, 4.794456, 
    4.798588, 4.805271, 4.813842, 4.823527, 4.833501, 4.842969, 4.851245, 
    4.857827,
  // momentumX(20,2, 0-49)
    4.864428, 4.86499, 4.867573, 4.871808, 4.877315, 4.883739, 4.890766, 
    4.898131, 4.905627, 4.913094, 4.920412, 4.927494, 4.934264, 4.94065, 
    4.946568, 4.951439, 4.958696, 4.962821, 4.966372, 4.969354, 4.971641, 
    4.973957, 4.97509, 4.97507, 4.97349, 4.970134, 4.964743, 4.957186, 
    4.947346, 4.935463, 4.921481, 4.90663, 4.890397, 4.873343, 4.856158, 
    4.839617, 4.824526, 4.811648, 4.801634, 4.794953, 4.791851, 4.792322, 
    4.79611, 4.802735, 4.811536, 4.821715, 4.832422, 4.842813, 4.852137, 
    4.85981,
  // momentumX(20,3, 0-49)
    4.866155, 4.86705, 4.869899, 4.874338, 4.879996, 4.886528, 4.893631, 
    4.90105, 4.908585, 4.916081, 4.923425, 4.930527, 4.937315, 4.943715, 
    4.949641, 4.954255, 4.962042, 4.966132, 4.969641, 4.972626, 4.974976, 
    4.977679, 4.979204, 4.979639, 4.978534, 4.975669, 4.970754, 4.963642, 
    4.954173, 4.94259, 4.928738, 4.914125, 4.897903, 4.880599, 4.862891, 
    4.845562, 4.829454, 4.815392, 4.804106, 4.796156, 4.791875, 4.791333, 
    4.794338, 4.800455, 4.809047, 4.819333, 4.830458, 4.841559, 4.851843, 
    4.860661,
  // momentumX(20,4, 0-49)
    4.867635, 4.868824, 4.871896, 4.876496, 4.882263, 4.888866, 4.896011, 
    4.903454, 4.910999, 4.918499, 4.925837, 4.932927, 4.939702, 4.946087, 
    4.952006, 4.956291, 4.964385, 4.968431, 4.971873, 4.974825, 4.977198, 
    4.980241, 4.982126, 4.982999, 4.982406, 4.980123, 4.975844, 4.969408, 
    4.960617, 4.949678, 4.936331, 4.922343, 4.906526, 4.889344, 4.871434, 
    4.85356, 4.836578, 4.82136, 4.808711, 4.799289, 4.793529, 4.791602, 
    4.793405, 4.798576, 4.80653, 4.816529, 4.827738, 4.8393, 4.850401, 
    4.860345,
  // momentumX(20,5, 0-49)
    4.868941, 4.870391, 4.873652, 4.878376, 4.884216, 4.890854, 4.898007, 
    4.905436, 4.912956, 4.920418, 4.927711, 4.934752, 4.941473, 4.947814, 
    4.953711, 4.957606, 4.965757, 4.969759, 4.973117, 4.976005, 4.978372, 
    4.981693, 4.983891, 4.98517, 4.985097, 4.983453, 4.979932, 4.97436, 
    4.966503, 4.956503, 4.944001, 4.930983, 4.915935, 4.899241, 4.881466, 
    4.863327, 4.845665, 4.82938, 4.815343, 4.80431, 4.796834, 4.793207, 
    4.793438, 4.797264, 4.804183, 4.813521, 4.824488, 4.836249, 4.84799, 
    4.858978,
  // momentumX(20,6, 0-49)
    4.870184, 4.871867, 4.875287, 4.880104, 4.885983, 4.892617, 4.899735, 
    4.907109, 4.914557, 4.921935, 4.929136, 4.936078, 4.942703, 4.948964, 
    4.95482, 4.958287, 4.966236, 4.970192, 4.97346, 4.976264, 4.978598, 
    4.982133, 4.984593, 4.986225, 4.986656, 4.985677, 4.982993, 4.978419, 
    4.971696, 4.962874, 4.95149, 4.939726, 4.925767, 4.9099, 4.892593, 
    4.874488, 4.856383, 4.83918, 4.823804, 4.8111, 4.801749, 4.796178, 
    4.794536, 4.796683, 4.802223, 4.810569, 4.820991, 4.832695, 4.844877, 
    4.856782,
  // momentumX(20,7, 0-49)
    4.871486, 4.873385, 4.876938, 4.881816, 4.887699, 4.894289, 4.901329, 
    4.908598, 4.915922, 4.923161, 4.930209, 4.936997, 4.943477, 4.949618, 
    4.955414, 4.958443, 4.965936, 4.969844, 4.97302, 4.975732, 4.978019, 
    4.981705, 4.984363, 4.986288, 4.987187, 4.986865, 4.985055, 4.981565, 
    4.976113, 4.968638, 4.958585, 4.948279, 4.935663, 4.92091, 4.904378, 
    4.886606, 4.868324, 4.850407, 4.833809, 4.819458, 4.808159, 4.800493, 
    4.796761, 4.796972, 4.800858, 4.807934, 4.81755, 4.828959, 4.841378, 
    4.854039,
  // momentumX(20,8, 0-49)
    4.872965, 4.875064, 4.878729, 4.883643, 4.889493, 4.895999, 4.902913, 
    4.910024, 4.917163, 4.924199, 4.931038, 4.937615, 4.943896, 4.949877, 
    4.955583, 4.958203, 4.965009, 4.968857, 4.971947, 4.974571, 4.976808, 
    4.980578, 4.983373, 4.98552, 4.986834, 4.987137, 4.986202, 4.983829, 
    4.979728, 4.973704, 4.965117, 4.956395, 4.945295, 4.931881, 4.916384, 
    4.899226, 4.88104, 4.862648, 4.845007, 4.829113, 4.815887, 4.806065, 
    4.800118, 4.798223, 4.800258, 4.805854, 4.81445, 4.825356, 4.837813, 
    4.851048,
  // momentumX(20,9, 0-49)
    4.874715, 4.877008, 4.88077, 4.885693, 4.891478, 4.897859, 4.904594, 
    4.911492, 4.918387, 4.925161, 4.931726, 4.938032, 4.944063, 4.949836, 
    4.955409, 4.957707, 4.963628, 4.967393, 4.970406, 4.972955, 4.975152, 
    4.978941, 4.981811, 4.984108, 4.985774, 4.98665, 4.986557, 4.985291, 
    4.982565, 4.978032, 4.970989, 4.96389, 4.954402, 4.942473, 4.928211, 
    4.911908, 4.894079, 4.87547, 4.857014, 4.839749, 4.824699, 4.812755, 
    4.804565, 4.800483, 4.800548, 4.804519, 4.811933, 4.82216, 4.834473, 
    4.848091,
  // momentumX(20,10, 0-49)
    4.876799, 4.879285, 4.883133, 4.888045, 4.893735, 4.899947, 4.906461, 
    4.913087, 4.919682, 4.926131, 4.932365, 4.938345, 4.944074, 4.949587, 
    4.954967, 4.957089, 4.961978, 4.965627, 4.968569, 4.971067, 4.973243, 
    4.97699, 4.979874, 4.98225, 4.984199, 4.985584, 4.986276, 4.986076, 
    4.984701, 4.981645, 4.976162, 4.970654, 4.962789, 4.952418, 4.939521, 
    4.924259, 4.907021, 4.88845, 4.869433, 4.851023, 4.834328, 4.82038, 
    4.810005, 4.803736, 4.801787, 4.804056, 4.810177, 4.819589, 4.831591, 
    4.845403,
  // momentumX(20,11, 0-49)
    4.879239, 4.881923, 4.885851, 4.890735, 4.896304, 4.902315, 4.908561, 
    4.91487, 4.921111, 4.927186, 4.933039, 4.938643, 4.944018, 4.949213, 
    4.954324, 4.956469, 4.960239, 4.963728, 4.966609, 4.969083, 4.971266, 
    4.974913, 4.977757, 4.980145, 4.982306, 4.984129, 4.985535, 4.986328, 
    4.986242, 4.98461, 4.980663, 4.976647, 4.97035, 4.961532, 4.950062, 
    4.935967, 4.919504, 4.901208, 4.881889, 4.862591, 4.844482, 4.828718, 
    4.816289, 4.807916, 4.80398, 4.804524, 4.80929, 4.81778, 4.829328, 
    4.843155,
  // momentumX(20,12, 0-49)
    4.88201, 4.884904, 4.888915, 4.893763, 4.899191, 4.904974, 4.910917, 
    4.916871, 4.922716, 4.928374, 4.933802, 4.938989, 4.943964, 4.948782, 
    4.953533, 4.95595, 4.958569, 4.961857, 4.964685, 4.967168, 4.969397, 
    4.972889, 4.975645, 4.977991, 4.980297, 4.982482, 4.984518, 4.986214, 
    4.987322, 4.987028, 4.984559, 4.981891, 4.977048, 4.969718, 4.959666, 
    4.946801, 4.93125, 4.913426, 4.894051, 4.874133, 4.854875, 4.837531, 
    4.823242, 4.812902, 4.807063, 4.805912, 4.809299, 4.816798, 4.827771, 
    4.841449,
  // momentumX(20,13, 0-49)
    4.885045, 4.888165, 4.892267, 4.897079, 4.902358, 4.907895, 4.913514, 
    4.919086, 4.924509, 4.929721, 4.934696, 4.939434, 4.943967, 4.948348, 
    4.952642, 4.955595, 4.957088, 4.960145, 4.962937, 4.965468, 4.967791, 
    4.971079, 4.973709, 4.975964, 4.978357, 4.980833, 4.98341, 4.985902, 
    4.98809, 4.989025, 4.987952, 4.986454, 4.982911, 4.976952, 4.968254, 
    4.956622, 4.942061, 4.92486, 4.905646, 4.885368, 4.865235, 4.846574, 
    4.830656, 4.818532, 4.810918, 4.808143, 4.810166, 4.816629, 4.826932, 
    4.840311,
  // momentumX(20,14, 0-49)
    4.888229, 4.8916, 4.895807, 4.900593, 4.905726, 4.911015, 4.916304, 
    4.921482, 4.92647, 4.931225, 4.935732, 4.940003, 4.944067, 4.947958, 
    4.951711, 4.955437, 4.955875, 4.958696, 4.961479, 4.964108, 4.966577, 
    4.969624, 4.9721, 4.974234, 4.976667, 4.979364, 4.98239, 4.985562, 
    4.988698, 4.990733, 4.990968, 4.99044, 4.988013, 4.983267, 4.975816, 
    4.965367, 4.951819, 4.935346, 4.916467, 4.896061, 4.875321, 4.855616, 
    4.838318, 4.824619, 4.815388, 4.811089, 4.811786, 4.817195, 4.826753, 
    4.839705,
  // momentumX(20,15, 0-49)
    4.891417, 4.895063, 4.899403, 4.904181, 4.909182, 4.914233, 4.919199, 
    4.923991, 4.928551, 4.932856, 4.936903, 4.940707, 4.944289, 4.947664, 
    4.950818, 4.955467, 4.954948, 4.957564, 4.96039, 4.963179, 4.965862, 
    4.968639, 4.970955, 4.972952, 4.975391, 4.978249, 4.981628, 4.985358, 
    4.989294, 4.99229, 4.993727, 4.993963, 4.99245, 4.988739, 4.982389, 
    4.973036, 4.96048, 4.944787, 4.926372, 4.906035, 4.884928, 4.864438, 
    4.846014, 4.830963, 4.820285, 4.814578, 4.81401, 4.818363, 4.827119, 
    4.839538,
  // momentumX(20,16, 0-49)
    4.894438, 4.898385, 4.902883, 4.90768, 4.912577, 4.917415, 4.922084, 
    4.926518, 4.93068, 4.934565, 4.938181, 4.941544, 4.944665, 4.94753, 
    4.950081, 4.955651, 4.954271, 4.956758, 4.959707, 4.962741, 4.965721, 
    4.968219, 4.970386, 4.972255, 4.974681, 4.977648, 4.981289, 4.985443, 
    4.990022, 4.993821, 4.99635, 4.997137, 4.996331, 4.993463, 4.98805, 
    4.97967, 4.968042, 4.953138, 4.935272, 4.915156, 4.893888, 4.87285, 
    4.853538, 4.837351, 4.825407, 4.818417, 4.816652, 4.819967, 4.827884, 
    4.839682,
  // momentumX(20,17, 0-49)
    4.897111, 4.901378, 4.906057, 4.910903, 4.915725, 4.920388, 4.924805, 
    4.92893, 4.93275, 4.936276, 4.939528, 4.942516, 4.945239, 4.947652, 
    4.949658, 4.955938, 4.95375, 4.956237, 4.959424, 4.962814, 4.966193, 
    4.968428, 4.970485, 4.972262, 4.974679, 4.977714, 4.981524, 4.985966, 
    4.991012, 4.995444, 4.99893, 5.000061, 4.999754, 4.997528, 4.992876, 
    4.985324, 4.974533, 4.960389, 4.943113, 4.92333, 4.90207, 4.880688, 
    4.860705, 4.843585, 4.830546, 4.822402, 4.819518, 4.82182, 4.828876, 
    4.839989,
  // momentumX(20,18, 0-49)
    4.899259, 4.903844, 4.908713, 4.913628, 4.918412, 4.922945, 4.927167, 
    4.931057, 4.934627, 4.9379, 4.940901, 4.943637, 4.946083, 4.948168, 
    4.94976, 4.956294, 4.953275, 4.955921, 4.959491, 4.963376, 4.967283, 
    4.969299, 4.971318, 4.973071, 4.97551, 4.97859, 4.98248, 4.987064, 
    4.992386, 4.997256, 5.001545, 5.002809, 5.002788, 5.001004, 4.996927, 
    4.990052, 4.979986, 4.966546, 4.949867, 4.930487, 4.909364, 4.887812, 
    4.867347, 4.849483, 4.83551, 4.826337, 4.822413, 4.823737, 4.829926, 
    4.840314,
  // momentumX(20,19, 0-49)
    4.900722, 4.905582, 4.910621, 4.915603, 4.920366, 4.924819, 4.928921, 
    4.932685, 4.936142, 4.939328, 4.942264, 4.944942, 4.947306, 4.949254, 
    4.950626, 4.956723, 4.952731, 4.955709, 4.959822, 4.964365, 4.968961, 
    4.970843, 4.972939, 4.974776, 4.977301, 4.980426, 4.984317, 4.988889, 
    4.994273, 4.99935, 5.004237, 5.005415, 5.005468, 5.00392, 5.000231, 
    4.993872, 4.984408, 4.971598, 4.9555, 4.936566, 4.915679, 4.894096, 
    4.873318, 4.854876, 4.840123, 4.83004, 4.825162, 4.825555, 4.830888, 
    4.840529,
  // momentumX(20,20, 0-49)
    4.90239, 4.908547, 4.914843, 4.921025, 4.926898, 4.932327, 4.937214, 
    4.9415, 4.945158, 4.948183, 4.950596, 4.952441, 4.953793, 4.954744, 
    4.955407, 0, 4.958249, 4.960236, 4.962961, 4.965996, 4.969181, 4.968955, 
    4.969491, 4.97025, 4.972277, 4.975456, 4.979868, 4.985317, 4.991841, 
    4.998215, 5.004694, 5.006587, 5.007314, 5.006402, 5.00332, 4.997553, 
    4.988664, 4.976397, 4.960779, 4.942212, 4.921516, 4.899904, 4.878851, 
    4.859899, 4.844436, 4.83351, 4.827723, 4.827208, 4.831687, 4.840559,
  // momentumX(20,21, 0-49)
    4.902546, 4.909152, 4.915813, 4.922264, 4.928308, 4.93382, 4.938725, 
    4.942987, 4.946609, 4.949608, 4.952027, 4.953918, 4.955361, 4.956449, 
    4.957307, 0, 4.95625, 4.958742, 4.96202, 4.965616, 4.96931, 4.968532, 
    4.968688, 4.969118, 4.970976, 4.974154, 4.978734, 4.984498, 4.991485, 
    4.998459, 5.005868, 5.007966, 5.009057, 5.008655, 5.006201, 5.001147, 
    4.99302, 4.981514, 4.966591, 4.948582, 4.928237, 4.906707, 4.885434, 
    4.865964, 4.849724, 4.837832, 4.830966, 4.829334, 4.832719, 4.840568,
  // momentumX(20,22, 0-49)
    4.902033, 4.909122, 4.916215, 4.92303, 4.929366, 4.935092, 4.940144, 
    4.944501, 4.948182, 4.951223, 4.953678, 4.955619, 4.957127, 4.958311, 
    4.959311, 0, 4.955119, 4.958027, 4.96179, 4.965904, 4.970087, 4.968813, 
    4.968649, 4.968804, 4.970531, 4.973706, 4.978404, 4.984384, 4.991682, 
    4.999045, 5.007104, 5.009167, 5.010358, 5.010189, 5.00809, 5.003501, 
    4.995925, 4.985018, 4.970692, 4.953214, 4.933263, 4.911923, 4.89059, 
    4.870792, 4.853981, 4.841319, 4.833551, 4.830953, 4.833365, 4.84028,
  // momentumX(20,23, 0-49)
    4.900946, 4.908532, 4.916096, 4.92334, 4.930048, 4.936085, 4.941385, 
    4.945931, 4.949752, 4.952897, 4.955433, 4.95744, 4.959013, 4.96027, 
    4.961375, 0, 4.954969, 4.958154, 4.962238, 4.966699, 4.971208, 4.969459, 
    4.96897, 4.968847, 4.970413, 4.973536, 4.978281, 4.984387, 4.991886, 
    4.999502, 5.008006, 5.009949, 5.011131, 5.011066, 5.009185, 5.00492, 
    4.99776, 4.987338, 4.973525, 4.956533, 4.936977, 4.915878, 4.894584, 
    4.874597, 4.857371, 4.844103, 4.835588, 4.832156, 4.833704, 4.839765,
  // momentumX(20,24, 0-49)
    4.899428, 4.907504, 4.915555, 4.92326, 4.930388, 4.936795, 4.942407, 
    4.947209, 4.951232, 4.95453, 4.957183, 4.959279, 4.96092, 4.962241, 
    4.963425, 0, 4.95597, 4.959291, 4.963529, 4.968157, 4.972827, 4.970741, 
    4.970021, 4.969701, 4.971145, 4.974215, 4.978966, 4.985128, 4.992729, 
    5.000482, 5.009243, 5.011076, 5.012208, 5.012159, 5.010361, 5.006243, 
    4.999289, 4.98912, 4.975582, 4.958858, 4.939522, 4.918553, 4.897259, 
    4.877122, 4.859592, 4.845881, 4.836812, 4.832757, 4.833642, 4.839036,
  // momentumX(20,25, 0-49)
    4.897653, 4.906196, 4.91472, 4.922887, 4.93045, 4.937253, 4.943209, 
    4.948304, 4.952564, 4.956049, 4.958841, 4.961037, 4.962751, 4.964127, 
    4.965363, 0, 4.957728, 4.961046, 4.96527, 4.969884, 4.974544, 4.972311, 
    4.971497, 4.971106, 4.972506, 4.975554, 4.980302, 4.986476, 4.994102, 
    5.001885, 5.010712, 5.012488, 5.013579, 5.013506, 5.011698, 5.007585, 
    5.000655, 4.990522, 4.977032, 4.960351, 4.941041, 4.920062, 4.898702, 
    4.878432, 4.860693, 4.846697, 4.837277, 4.832819, 4.833266, 4.838201,
  // momentumX(20,26, 0-49)
    4.895818, 4.904783, 4.913742, 4.922344, 4.930325, 4.937515, 4.943821, 
    4.949216, 4.953726, 4.957407, 4.960343, 4.962636, 4.964409, 4.965817, 
    4.967063, 0, 4.960133, 4.963308, 4.967357, 4.971776, 4.976251, 4.974082, 
    4.973327, 4.973009, 4.974462, 4.977538, 4.982289, 4.98844, 4.996022, 
    5.003737, 5.012439, 5.014235, 5.015309, 5.015183, 5.013282, 5.009041, 
    5.001948, 4.99163, 4.97794, 4.961062, 4.941566, 4.920424, 4.898925, 
    4.878536, 4.860688, 4.846581, 4.837034, 4.832421, 4.832682, 4.8374,
  // momentumX(20,27, 0-49)
    4.894114, 4.903435, 4.912771, 4.921757, 4.930116, 4.937665, 4.944301, 
    4.949985, 4.954732, 4.958596, 4.961658, 4.964022, 4.965817, 4.967206, 
    4.968397, 0, 4.96324, 4.966122, 4.969824, 4.973864, 4.97798, 4.976048, 
    4.975473, 4.975338, 4.976915, 4.98005, 4.984796, 4.990885, 4.998345, 
    5.00589, 5.014274, 5.016143, 5.01721, 5.016988, 5.014902, 5.010391, 
    5.002958, 4.992247, 4.978143, 4.960862, 4.941015, 4.919603, 4.897938, 
    4.87749, 4.859674, 4.845661, 4.836235, 4.831735, 4.832074, 4.836821,
  // momentumX(20,28, 0-49)
    4.892716, 4.902316, 4.911954, 4.921258, 4.92994, 4.937809, 4.94474, 
    4.950686, 4.955645, 4.959659, 4.962801, 4.965176, 4.966919, 4.9682, 
    4.969231, 0, 4.967395, 4.969824, 4.972999, 4.976473, 4.980055, 4.978459, 
    4.97812, 4.978223, 4.979947, 4.983134, 4.987837, 4.993802, 5.001053, 
    5.008318, 5.016205, 5.018162, 5.019183, 5.018777, 5.016371, 5.011417, 
    5.00344, 4.992121, 4.977393, 4.95953, 4.939205, 4.917471, 4.895676, 
    4.875288, 4.8577, 4.844033, 4.835011, 4.830916, 4.831614, 4.836638,
  // momentumX(20,29, 0-49)
    4.891768, 4.901561, 4.91142, 4.920973, 4.929929, 4.938075, 4.945275, 
    4.951451, 4.956579, 4.960682, 4.963824, 4.966108, 4.967679, 4.968717, 
    4.969442, 0, 4.972353, 4.974166, 4.976633, 4.979355, 4.982222, 4.980926, 
    4.980772, 4.981068, 4.982892, 4.986081, 4.990681, 4.996451, 5.003397, 
    5.010265, 5.017463, 5.019434, 5.020311, 5.019595, 5.016734, 5.011202, 
    5.002559, 4.990538, 4.975133, 4.956691, 4.935954, 4.914032, 4.892297, 
    4.872213, 4.855128, 4.842093, 4.833755, 4.830319, 4.831594, 4.837072,
  // momentumX(20,30, 0-49)
    4.890552, 4.899473, 4.908428, 4.917069, 4.925149, 4.932522, 4.939125, 
    4.94497, 4.950115, 4.954631, 4.958583, 4.961999, 4.964857, 4.967066, 
    4.968472, 4.979602, 4.96907, 4.971892, 4.976008, 4.980648, 4.98542, 
    4.986781, 4.988743, 4.990612, 4.993301, 4.996634, 5.000715, 5.005429, 
    5.010921, 5.01609, 5.021275, 5.022079, 5.021772, 5.019878, 5.015864, 
    5.009229, 4.99956, 4.986626, 4.970476, 4.951515, 4.930534, 4.90868, 
    4.887331, 4.867914, 4.851709, 4.839678, 4.832371, 4.829907, 4.832027, 
    4.838179,
  // momentumX(20,31, 0-49)
    4.890921, 4.899925, 4.908952, 4.91766, 4.925797, 4.93321, 4.939828, 
    4.945653, 4.950732, 4.95514, 4.958956, 4.962236, 4.965003, 4.967213, 
    4.968752, 4.979363, 4.971177, 4.97361, 4.977141, 4.98109, 4.985148, 
    4.986675, 4.988585, 4.990395, 4.993023, 4.996342, 5.00046, 5.005226, 
    5.010689, 5.015679, 5.020274, 5.021196, 5.02085, 5.01876, 5.014407, 
    5.007318, 4.997122, 4.983652, 4.967027, 4.947731, 4.926632, 4.904924, 
    4.883998, 4.865252, 4.849897, 4.83881, 4.832448, 4.830843, 4.833675, 
    4.840341,
  // momentumX(20,32, 0-49)
    4.891858, 4.900726, 4.909607, 4.918174, 4.926184, 4.933486, 4.940012, 
    4.945757, 4.950766, 4.955113, 4.958885, 4.962158, 4.964985, 4.967364, 
    4.969228, 4.978518, 4.972463, 4.974708, 4.977826, 4.98125, 4.984755, 
    4.986572, 4.988569, 4.990442, 4.993085, 4.996394, 5.000472, 5.005139, 
    5.010365, 5.014951, 5.01875, 5.019603, 5.019039, 5.016583, 5.011744, 
    5.004078, 4.993276, 4.979236, 4.962163, 4.942626, 4.921564, 4.900208, 
    4.879947, 4.86213, 4.847888, 4.837993, 4.832799, 4.832254, 4.835965, 
    4.843286,
  // momentumX(20,33, 0-49)
    4.893402, 4.901961, 4.910522, 4.918782, 4.926514, 4.933579, 4.93991, 
    4.945505, 4.950407, 4.954688, 4.958445, 4.961763, 4.964719, 4.96735, 
    4.96964, 4.977197, 4.973083, 4.975312, 4.978167, 4.981205, 4.984287, 
    4.986477, 4.98866, 4.990693, 4.993394, 4.996678, 5.000629, 5.005051, 
    5.009844, 5.013827, 5.016671, 5.017282, 5.016326, 5.013347, 5.00788, 
    4.999536, 4.988063, 4.973445, 4.955978, 4.936319, 4.915467, 4.894683, 
    4.87533, 4.858694, 4.845803, 4.83732, 4.833489, 4.834168, 4.838899, 
    4.846986,
  // momentumX(20,34, 0-49)
    4.89555, 4.903658, 4.911766, 4.919588, 4.926923, 4.933646, 4.939695, 
    4.945072, 4.949821, 4.954011, 4.957741, 4.961105, 4.964197, 4.967091, 
    4.969819, 4.975549, 4.97322, 4.975553, 4.978248, 4.981001, 4.983756, 
    4.986354, 4.988786, 4.991036, 4.993814, 4.997042, 5.000778, 5.004812, 
    5.008993, 5.012204, 5.01397, 5.014173, 5.01267, 5.009023, 5.002813, 
    4.993709, 4.981535, 4.966369, 4.9486, 4.928967, 4.908524, 4.88854, 
    4.870338, 4.855117, 4.843793, 4.836905, 4.834589, 4.836618, 4.842463, 
    4.851387,
  // momentumX(20,35, 0-49)
    4.898267, 4.905814, 4.913355, 4.920641, 4.92749, 4.933788, 4.939488, 
    4.944591, 4.949139, 4.953203, 4.956876, 4.960257, 4.963455, 4.966567, 
    4.969674, 4.973719, 4.973058, 4.975548, 4.978137, 4.98067, 4.983167, 
    4.986171, 4.988875, 4.991373, 4.994223, 4.997348, 5.000774, 5.004288, 
    5.007689, 5.009979, 5.010575, 5.010211, 5.008013, 5.003575, 4.996533, 
    4.986623, 4.973759, 4.958113, 4.940172, 4.920749, 4.900939, 4.881996, 
    4.865181, 4.851587, 4.842009, 4.83686, 4.836168, 4.83962, 4.846628, 
    4.856417,
  // momentumX(20,36, 0-49)
    4.901495, 4.908389, 4.915284, 4.921958, 4.92825, 4.934066, 4.939364, 
    4.944149, 4.948456, 4.952359, 4.955939, 4.959299, 4.962548, 4.965801, 
    4.969179, 4.971826, 4.972733, 4.975375, 4.977877, 4.980225, 4.982509, 
    4.985884, 4.988856, 4.991599, 4.994495, 4.99746, 5.00048, 5.003342, 
    5.005812, 5.007051, 5.006406, 5.005326, 5.002304, 4.996975, 4.989042, 
    4.97832, 4.964816, 4.948807, 4.930867, 4.911874, 4.892938, 4.87528, 
    4.860076, 4.848299, 4.84061, 4.837299, 4.838289, 4.843188, 4.85136, 
    4.861993,
  // momentumX(20,37, 0-49)
    4.905167, 4.911334, 4.917521, 4.923526, 4.929215, 4.934506, 4.939363, 
    4.943795, 4.947833, 4.95154, 4.954994, 4.958288, 4.961529, 4.964836, 
    4.968349, 4.969948, 4.972336, 4.975077, 4.977478, 4.979656, 4.981754, 
    4.985441, 4.988646, 4.991607, 4.994504, 4.99724, 4.999755, 5.001844, 
    5.003247, 5.003323, 5.001387, 4.999458, 4.995503, 4.989217, 4.980371, 
    4.968874, 4.954834, 4.938624, 4.9209, 4.902584, 4.884777, 4.868644, 
    4.855253, 4.845448, 4.839749, 4.838326, 4.841006, 4.847328, 4.856611, 
    4.868018,
  // momentumX(20,38, 0-49)
    4.909193, 4.914583, 4.920015, 4.925317, 4.930371, 4.935106, 4.939497, 
    4.943548, 4.947289, 4.950776, 4.954073, 4.957259, 4.960435, 4.96371, 
    4.967225, 4.968122, 4.971893, 4.974655, 4.976923, 4.97893, 4.980852, 
    4.984771, 4.988155, 4.991285, 4.994119, 4.996551, 4.998464, 4.999669, 
    4.999884, 4.99871, 4.995449, 4.992558, 4.987595, 4.98032, 4.970589, 
    4.958406, 4.943982, 4.927779, 4.910518, 4.893145, 4.876726, 4.862342, 
    4.85094, 4.84322, 4.839568, 4.840035, 4.844362, 4.852028, 4.862319, 
    4.874377,
  // momentumX(20,39, 0-49)
    4.913477, 4.918053, 4.922704, 4.927279, 4.931678, 4.93584, 4.939745, 
    4.943396, 4.946823, 4.950062, 4.953173, 4.956218, 4.959277, 4.962446, 
    4.965847, 4.966341, 4.971383, 4.974071, 4.976166, 4.977993, 4.979737, 
    4.983795, 4.987283, 4.990516, 4.993211, 4.995252, 4.99647, 4.996691, 
    4.995628, 4.99314, 4.988544, 4.984612, 4.978605, 4.970356, 4.959818, 
    4.94709, 4.932482, 4.916533, 4.900011, 4.883851, 4.869068, 4.856631, 
    4.847351, 4.841784, 4.840184, 4.842492, 4.848373, 4.857256, 4.868401, 
    4.880943,
  // momentumX(20,40, 0-49)
    4.917906, 4.921646, 4.925501, 4.929339, 4.933074, 4.936653, 4.940061, 
    4.9433, 4.946392, 4.949367, 4.952266, 4.955137, 4.958039, 4.961041, 
    4.964238, 4.964564, 4.970736, 4.97326, 4.975143, 4.976772, 4.978323, 
    4.982419, 4.985922, 4.989172, 4.991644, 4.993212, 4.993649, 4.99281, 
    4.990404, 4.98657, 4.980658, 4.975645, 4.968606, 4.959457, 4.948241, 
    4.93516, 4.920611, 4.905192, 4.889691, 4.87501, 4.86208, 4.851747, 
    4.844676, 4.84128, 4.841683, 4.845729, 4.853019, 4.862945, 4.874746, 
    4.887564,
  // momentumX(20,41, 0-49)
    4.922345, 4.925241, 4.928298, 4.9314, 4.934471, 4.937466, 4.940372, 
    4.943191, 4.945935, 4.948627, 4.951293, 4.953965, 4.956676, 4.95947, 
    4.9624, 4.962718, 4.969854, 4.972135, 4.973769, 4.975179, 4.976512, 
    4.980538, 4.983962, 4.987133, 4.989291, 4.9903, 4.98989, 4.987938, 
    4.984165, 4.978992, 4.971818, 4.965739, 4.957735, 4.94781, 4.936104, 
    4.92291, 4.908694, 4.894094, 4.879889, 4.866925, 4.856025, 4.847902, 
    4.84307, 4.841802, 4.844105, 4.849738, 4.858246, 4.868992, 4.881212, 
    4.894058,
  // momentumX(20,42, 0-49)
    4.926642, 4.928699, 4.930964, 4.93334, 4.935758, 4.938178, 4.940584, 
    4.942979, 4.945368, 4.947763, 4.950179, 4.95263, 4.955127, 4.957681, 
    4.960309, 4.96071, 4.96862, 4.970598, 4.971952, 4.973114, 4.974197, 
    4.978046, 4.981288, 4.98428, 4.986035, 4.986415, 4.985108, 4.982025, 
    4.976905, 4.970449, 4.962109, 4.955034, 4.946192, 4.935675, 4.923714, 
    4.910677, 4.897085, 4.88359, 4.870934, 4.859879, 4.851132, 4.845262, 
    4.842635, 4.843394, 4.847439, 4.854456, 4.863945, 4.875252, 4.887619, 
    4.900222,
  // momentumX(20,43, 0-49)
    4.930626, 4.931849, 4.933344, 4.935014, 4.936798, 4.938658, 4.940579, 
    4.942554, 4.944587, 4.94668, 4.948834, 4.951047, 4.953313, 4.955612, 
    4.957922, 4.958442, 4.966921, 4.968552, 4.9696, 4.970482, 4.971275, 
    4.974844, 4.977806, 4.980515, 4.981785, 4.981482, 4.979256, 4.975064, 
    4.968668, 4.961029, 4.951668, 4.943729, 4.934234, 4.923361, 4.911418, 
    4.898832, 4.886153, 4.874021, 4.86312, 4.854114, 4.847578, 4.843935, 
    4.843416, 4.846041, 4.851618, 4.85977, 4.869962, 4.881538, 4.893755, 
    4.905829,
  // momentumX(20,44, 0-49)
    4.93411, 4.934515, 4.935261, 4.936253, 4.937433, 4.938762, 4.940217, 
    4.941791, 4.943477, 4.94527, 4.94716, 4.949131, 4.951157, 4.953195, 
    4.955183, 4.955816, 4.964656, 4.965913, 4.966628, 4.967195, 4.967651, 
    4.970848, 4.973435, 4.975765, 4.976482, 4.975461, 4.972332, 4.967094, 
    4.959548, 4.950883, 4.940692, 4.93208, 4.922171, 4.911213, 4.89958, 
    4.887739, 4.876243, 4.865695, 4.856701, 4.849814, 4.845474, 4.843967, 
    4.845396, 4.84967, 4.856519, 4.865516, 4.876104, 4.887634, 4.899394, 
    4.910653,
  // momentumX(20,45, 0-49)
    4.936903, 4.936502, 4.936521, 4.936871, 4.937485, 4.938321, 4.939349, 
    4.940551, 4.941915, 4.943424, 4.945058, 4.946791, 4.948578, 4.950358, 
    4.952039, 4.952745, 4.961742, 4.962612, 4.962971, 4.963184, 4.963254, 
    4.965993, 4.968124, 4.96999, 4.970107, 4.968362, 4.964381, 4.958209, 
    4.949688, 4.940206, 4.929422, 4.920379, 4.910328, 4.899585, 4.888559, 
    4.877738, 4.867655, 4.858856, 4.851855, 4.847086, 4.844861, 4.845332, 
    4.848487, 4.854145, 4.861969, 4.87149, 4.882148, 4.893308, 4.904304, 
    4.914479,
  // momentumX(20,46, 0-49)
    4.938819, 4.937624, 4.936943, 4.936685, 4.936779, 4.93717, 4.937817, 
    4.938693, 4.939772, 4.94103, 4.942434, 4.943947, 4.945509, 4.947042, 
    4.948433, 4.949158, 4.958127, 4.958603, 4.958583, 4.958401, 4.958039, 
    4.960252, 4.961856, 4.963193, 4.962687, 4.960245, 4.955501, 4.948549, 
    4.939279, 4.929226, 4.918125, 4.908927, 4.899035, 4.888804, 4.878668, 
    4.869109, 4.860616, 4.853668, 4.848677, 4.845958, 4.845698, 4.847935, 
    4.852553, 4.859291, 4.86776, 4.877473, 4.887864, 4.898334, 4.908283, 
    4.91715,
  // momentumX(20,47, 0-49)
    4.93972, 4.937729, 4.936366, 4.935534, 4.935153, 4.935151, 4.935477, 
    4.936083, 4.936932, 4.937986, 4.939202, 4.940526, 4.941891, 4.9432, 
    4.944324, 4.945001, 4.953781, 4.953864, 4.95344, 4.952825, 4.951988, 
    4.953621, 4.954652, 4.955418, 4.954295, 4.951216, 4.945836, 4.938297, 
    4.928536, 4.918194, 4.907071, 4.898016, 4.888585, 4.879151, 4.870152, 
    4.862043, 4.85526, 4.850199, 4.847168, 4.84637, 4.847877, 4.851622, 
    4.857403, 4.864896, 4.873673, 4.883236, 4.893039, 4.902533, 4.911198, 
    4.918588,
  // momentumX(20,48, 0-49)
    4.939519, 4.93672, 4.934682, 4.933303, 4.932487, 4.932148, 4.932213, 
    4.932616, 4.933301, 4.934213, 4.935294, 4.936477, 4.937681, 4.938794, 
    4.939677, 4.940239, 4.948703, 4.94839, 4.94754, 4.946457, 4.945107, 
    4.946132, 4.946567, 4.946746, 4.945043, 4.94142, 4.935561, 4.927656, 
    4.917686, 4.907351, 4.896503, 4.88789, 4.879201, 4.870818, 4.863158, 
    4.856635, 4.85162, 4.848419, 4.847244, 4.848188, 4.851223, 4.856192, 
    4.862821, 4.870739, 4.879495, 4.888591, 4.89752, 4.905799, 4.913006, 
    4.918834,
  // momentumX(20,49, 0-49)
    4.940613, 4.936409, 4.933164, 4.930776, 4.929138, 4.928135, 4.927667, 
    4.927631, 4.927937, 4.928491, 4.9292, 4.92996, 4.930647, 4.931097, 
    4.931102, 4.930818, 4.946164, 4.943949, 4.940964, 4.937904, 4.934816, 
    4.936986, 4.938692, 4.94071, 4.939893, 4.93633, 4.929495, 4.919771, 
    4.907046, 4.894641, 4.882136, 4.8747, 4.867539, 4.861034, 4.855579, 
    4.851521, 4.849131, 4.84859, 4.849968, 4.853214, 4.858169, 4.864559, 
    4.872037, 4.88018, 4.888537, 4.896647, 4.90409, 4.910515, 4.915682, 
    4.919499,
  // momentumX(21,0, 0-49)
    4.867756, 4.87136, 4.876185, 4.881904, 4.888227, 4.894917, 4.901782, 
    4.908686, 4.915534, 4.922264, 4.928842, 4.935246, 4.941461, 4.947464, 
    4.953222, 4.958513, 4.964422, 4.96916, 4.973463, 4.977247, 4.98037, 
    4.982961, 4.984521, 4.984962, 4.984047, 4.981614, 4.977492, 4.971577, 
    4.963781, 4.95417, 4.942726, 4.929893, 4.915575, 4.900093, 4.883879, 
    4.867457, 4.851445, 4.836494, 4.823259, 4.812335, 4.804196, 4.799148, 
    4.797297, 4.798529, 4.802532, 4.808812, 4.816741, 4.82561, 4.834689, 
    4.843285,
  // momentumX(21,1, 0-49)
    4.869227, 4.873135, 4.878213, 4.88414, 4.890633, 4.897455, 4.904428, 
    4.911416, 4.918332, 4.925114, 4.931731, 4.938162, 4.944387, 4.950385, 
    4.956112, 4.961147, 4.967659, 4.972268, 4.976444, 4.980152, 4.983257, 
    4.986171, 4.988067, 4.988924, 4.988447, 4.98646, 4.982759, 4.977232, 
    4.969764, 4.960455, 4.949201, 4.93672, 4.922586, 4.907089, 4.890637, 
    4.87375, 4.857055, 4.841236, 4.827, 4.815002, 4.805791, 4.799745, 
    4.797029, 4.797587, 4.801143, 4.807224, 4.815208, 4.824379, 4.833981, 
    4.843285,
  // momentumX(21,2, 0-49)
    4.87042, 4.874584, 4.879874, 4.885972, 4.892601, 4.899534, 4.906593, 
    4.913648, 4.920613, 4.927431, 4.934066, 4.940497, 4.946706, 4.952666, 
    4.958333, 4.963048, 4.970029, 4.974471, 4.978471, 4.982044, 4.985077, 
    4.988253, 4.990441, 4.991687, 4.991656, 4.99017, 4.987002, 4.982033, 
    4.97512, 4.966384, 4.955632, 4.943846, 4.930265, 4.915128, 4.898799, 
    4.881767, 4.864641, 4.848114, 4.832927, 4.819794, 4.809337, 4.802019, 
    4.798089, 4.79757, 4.800246, 4.805697, 4.813336, 4.822461, 4.832316, 
    4.842153,
  // momentumX(21,3, 0-49)
    4.871417, 4.875794, 4.881257, 4.88749, 4.894225, 4.90124, 4.90836, 
    4.91546, 4.922452, 4.92928, 4.935906, 4.942309, 4.948469, 4.954359, 
    4.959938, 4.964278, 4.971559, 4.975809, 4.979591, 4.982981, 4.985889, 
    4.989264, 4.991691, 4.993279, 4.993685, 4.992729, 4.990175, 4.985899, 
    4.979735, 4.971802, 4.96182, 4.951028, 4.938334, 4.923909, 4.908056, 
    4.891205, 4.873922, 4.856891, 4.840857, 4.826586, 4.81477, 4.805964, 
    4.800524, 4.798568, 4.799973, 4.804396, 4.811304, 4.820037, 4.829866, 
    4.840038,
  // momentumX(21,4, 0-49)
    4.872332, 4.876885, 4.882481, 4.888814, 4.895623, 4.902688, 4.909839, 
    4.916954, 4.923941, 4.930746, 4.937329, 4.943668, 4.949744, 4.955535, 
    4.961005, 4.964917, 4.972301, 4.976346, 4.979885, 4.983051, 4.985792, 
    4.989301, 4.991906, 4.993781, 4.994592, 4.994171, 4.992283, 4.9888, 
    4.983535, 4.976586, 4.967588, 4.958031, 4.946498, 4.933095, 4.91804, 
    4.90169, 4.884544, 4.867239, 4.850518, 4.835167, 4.821952, 4.811521, 
    4.804342, 4.800659, 4.800459, 4.8035, 4.809333, 4.817359, 4.826887, 
    4.837183,
  // momentumX(21,5, 0-49)
    4.873298, 4.87799, 4.883683, 4.890078, 4.896924, 4.904002, 4.91115, 
    4.91824, 4.925184, 4.931925, 4.938425, 4.94466, 4.950615, 4.956275, 
    4.961616, 4.965065, 4.972339, 4.976171, 4.979454, 4.982371, 4.984913, 
    4.988491, 4.99121, 4.993308, 4.994482, 4.994578, 4.993377, 4.990749, 
    4.986489, 4.980652, 4.972798, 4.964639, 4.954481, 4.942347, 4.928371, 
    4.912815, 4.896089, 4.878769, 4.861557, 4.845256, 4.830675, 4.818562, 
    4.809506, 4.803884, 4.801821, 4.803196, 4.807662, 4.8147, 4.823673, 
    4.833878,
  // momentumX(21,6, 0-49)
    4.874443, 4.879241, 4.884993, 4.891414, 4.898254, 4.905306, 4.912405, 
    4.919427, 4.926284, 4.932917, 4.939289, 4.945377, 4.951174, 4.956671, 
    4.961865, 4.964837, 4.971784, 4.975398, 4.97842, 4.981078, 4.983403, 
    4.986985, 4.989758, 4.992006, 4.993488, 4.994068, 4.99355, 4.991801, 
    4.988611, 4.983963, 4.977353, 4.970687, 4.962039, 4.951355, 4.938675, 
    4.924161, 4.908125, 4.891047, 4.87358, 4.856506, 4.840674, 4.826908, 
    4.815924, 4.808243, 4.804142, 4.803638, 4.806506, 4.812325, 4.820523, 
    4.830435,
  // momentumX(21,7, 0-49)
    4.87588, 4.880752, 4.88653, 4.892937, 4.899731, 4.90671, 4.913714, 
    4.920619, 4.927339, 4.933815, 4.940012, 4.945911, 4.951509, 4.956812, 
    4.961838, 4.964347, 4.970757, 4.97415, 4.976916, 4.979318, 4.981421, 
    4.98495, 4.987716, 4.990044, 4.991772, 4.992788, 4.992926, 4.992055, 
    4.989957, 4.986527, 4.981206, 4.976059, 4.968983, 4.959855, 4.948626, 
    4.93535, 4.92023, 4.903647, 4.886172, 4.868548, 4.851635, 4.836328, 
    4.823456, 4.813686, 4.807459, 4.804945, 4.806056, 4.810474, 4.81771, 
    4.82715,
  // momentumX(21,8, 0-49)
    4.8777, 4.882618, 4.888388, 4.894741, 4.901444, 4.908303, 4.915162, 
    4.9219, 4.928433, 4.934703, 4.940678, 4.946343, 4.951704, 4.95678, 
    4.961609, 4.963711, 4.969393, 4.972557, 4.975082, 4.977241, 4.979133, 
    4.982553, 4.985257, 4.987593, 4.989506, 4.990901, 4.99165, 4.991627, 
    4.990613, 4.988391, 4.984363, 4.980696, 4.975188, 4.967651, 4.957954, 
    4.946052, 4.932031, 4.916164, 4.898924, 4.880996, 4.863228, 4.846558, 
    4.831919, 4.82012, 4.811763, 4.807185, 4.806442, 4.80934, 4.81547, 
    4.824277,
  // momentumX(21,9, 0-49)
    4.879959, 4.884899, 4.890628, 4.89689, 4.903462, 4.910154, 4.916817, 
    4.923337, 4.929632, 4.935648, 4.941355, 4.946746, 4.951833, 4.956645, 
    4.961241, 4.963027, 4.967825, 4.970748, 4.97305, 4.974993, 4.976692, 
    4.979956, 4.982547, 4.98483, 4.986863, 4.988575, 4.989882, 4.990657, 
    4.99069, 4.989635, 4.986869, 4.984592, 4.98059, 4.974617, 4.966471, 
    4.956012, 4.943221, 4.928251, 4.911475, 4.893493, 4.87512, 4.857318, 
    4.8411, 4.827405, 4.816993, 4.810369, 4.807745, 4.80905, 4.813972, 
    4.822018,
  // momentumX(21,10, 0-49)
    4.882683, 4.887622, 4.893283, 4.899419, 4.905817, 4.912298, 4.918719, 
    4.924973, 4.930984, 4.936702, 4.942099, 4.947176, 4.951952, 4.956465, 
    4.960778, 4.962388, 4.966177, 4.968843, 4.970945, 4.972705, 4.974249, 
    4.977313, 4.979748, 4.98192, 4.984013, 4.985978, 4.98778, 4.989291, 
    4.99031, 4.990362, 4.988803, 4.987789, 4.985182, 4.980694, 4.97406, 
    4.965057, 4.953567, 4.939633, 4.923513, 4.905717, 4.887003, 4.868331, 
    4.85077, 4.835371, 4.823044, 4.814457, 4.809978, 4.809673, 4.813326, 
    4.820508,
  // momentumX(21,11, 0-49)
    4.885859, 4.890782, 4.896351, 4.902331, 4.90852, 4.914749, 4.920887, 
    4.926834, 4.932517, 4.937896, 4.942946, 4.947676, 4.952104, 4.956275, 
    4.960248, 4.961854, 4.964558, 4.966954, 4.968882, 4.970501, 4.971934, 
    4.974759, 4.977002, 4.979015, 4.981116, 4.983275, 4.985504, 4.987677, 
    4.989609, 4.990688, 4.990268, 4.990361, 4.989007, 4.985883, 4.980674, 
    4.973091, 4.962924, 4.950112, 4.934801, 4.917403, 4.898602, 4.879333, 
    4.860695, 4.843828, 4.829777, 4.819361, 4.813109, 4.811215, 4.813574, 
    4.819819,
  // momentumX(21,12, 0-49)
    4.88944, 4.894337, 4.899799, 4.905598, 4.911548, 4.917494, 4.923313, 
    4.928915, 4.934238, 4.939242, 4.943916, 4.948267, 4.952316, 4.956103, 
    4.959673, 4.961469, 4.963051, 4.965169, 4.966954, 4.968485, 4.96986, 
    4.972414, 4.974438, 4.976257, 4.978319, 4.980617, 4.983204, 4.985958, 
    4.988717, 4.990734, 4.99138, 4.99241, 4.992143, 4.990234, 4.986331, 
    4.980086, 4.971216, 4.959564, 4.945173, 4.928348, 4.909691, 4.890091, 
    4.870652, 4.852578, 4.837027, 4.824958, 4.81705, 4.813632, 4.814701, 
    4.819964,
  // momentumX(21,13, 0-49)
    4.893345, 4.898217, 4.90356, 4.909164, 4.914856, 4.920492, 4.925966, 
    4.931196, 4.936131, 4.94074, 4.945012, 4.948959, 4.952602, 4.955966, 
    4.959073, 4.961245, 4.961709, 4.963559, 4.96524, 4.96674, 4.96812, 
    4.970376, 4.972166, 4.973768, 4.975757, 4.978142, 4.981021, 4.984272, 
    4.987758, 4.990619, 4.99226, 4.994047, 4.99469, 4.993832, 4.991089, 
    4.98607, 4.978432, 4.967936, 4.954527, 4.93841, 4.920095, 4.900408, 
    4.880437, 4.861424, 4.844614, 4.831095, 4.821679, 4.816827, 4.816639, 
    4.820898,
  // momentumX(21,14, 0-49)
    4.897468, 4.902321, 4.907547, 4.912951, 4.918373, 4.923688, 4.928799, 
    4.93364, 4.93817, 4.942365, 4.946223, 4.949754, 4.95297, 4.95588, 
    4.958479, 4.961169, 4.960548, 4.962161, 4.963795, 4.965333, 4.966787, 
    4.968728, 4.97028, 4.971656, 4.973548, 4.975982, 4.979085, 4.982744, 
    4.986854, 4.990458, 4.993018, 4.995389, 4.996763, 4.99678, 4.995036, 
    4.991111, 4.98461, 4.975227, 4.962822, 4.947505, 4.929689, 4.910128, 
    4.889874, 4.870183, 4.852361, 4.837605, 4.826849, 4.820671, 4.819281, 
    4.822535,
  // momentumX(21,15, 0-49)
    4.901683, 4.906533, 4.911652, 4.916859, 4.922011, 4.927, 4.931743, 
    4.936191, 4.94031, 4.944088, 4.94753, 4.950641, 4.953424, 4.955871, 
    4.957943, 4.96121, 4.959546, 4.960984, 4.962644, 4.9643, 4.965909, 
    4.967529, 4.968853, 4.970014, 4.971802, 4.974249, 4.977513, 4.981489, 
    4.986113, 4.990354, 4.993762, 4.996544, 4.998473, 4.999189, 4.998278, 
    4.995298, 4.989818, 4.981478, 4.970063, 4.955593, 4.938392, 4.919131, 
    4.898813, 4.878683, 4.860091, 4.844313, 4.832389, 4.825014, 4.822492, 
    4.824755,
  // momentumX(21,16, 0-49)
    4.905852, 4.910719, 4.915746, 4.92077, 4.925663, 4.930331, 4.934713, 
    4.938773, 4.942492, 4.945868, 4.948905, 4.951612, 4.953979, 4.955981, 
    4.95755, 4.961321, 4.958642, 4.960001, 4.961782, 4.963653, 4.965511, 
    4.966817, 4.967943, 4.968918, 4.970611, 4.973051, 4.976418, 4.980618, 
    4.985636, 4.9904, 4.994579, 4.99761, 4.999923, 5.001165, 5.00092, 
    4.99873, 4.994142, 4.986749, 4.976277, 4.962667, 4.946156, 4.927331, 
    4.907132, 4.886779, 4.86764, 4.851046, 4.838132, 4.82969, 4.826118, 
    4.82742,
  // momentumX(21,17, 0-49)
    4.909837, 4.914738, 4.919692, 4.924548, 4.929195, 4.93356, 4.9376, 
    4.941293, 4.944641, 4.947648, 4.950324, 4.95267, 4.954671, 4.956281, 
    4.957415, 4.961463, 4.957752, 4.959157, 4.961174, 4.963372, 4.965584, 
    4.966605, 4.967587, 4.968428, 4.970053, 4.97248, 4.975895, 4.980227, 
    4.985517, 4.99068, 4.995541, 4.998661, 5.001194, 5.002797, 5.003052, 
    5.001498, 4.997662, 4.991107, 4.98151, 4.968741, 4.95296, 4.934667, 
    4.914736, 4.894343, 4.874856, 4.857644, 4.843911, 4.834536, 4.83, 4.830382,
  // momentumX(21,18, 0-49)
    4.913497, 4.918441, 4.923331, 4.928032, 4.932451, 4.936535, 4.940263, 
    4.943635, 4.946665, 4.949371, 4.951762, 4.953833, 4.955557, 4.956873, 
    4.957686, 4.961622, 4.956789, 4.958377, 4.96076, 4.963412, 4.9661, 
    4.966885, 4.967799, 4.968584, 4.970194, 4.972615, 4.97604, 4.980412, 
    4.985839, 4.991264, 4.996696, 4.999753, 5.002348, 5.004149, 5.004743, 
    5.003669, 5.000443, 4.994608, 4.985798, 4.973829, 4.958785, 4.94109, 
    4.921543, 4.901266, 4.881607, 4.863956, 4.849568, 4.839391, 4.833985, 
    4.833497,
  // momentumX(21,19, 0-49)
    4.9167, 4.921665, 4.926477, 4.931019, 4.93522, 4.939054, 4.942522, 
    4.945646, 4.948455, 4.950972, 4.953205, 4.955136, 4.956722, 4.957885, 
    4.958528, 4.961836, 4.95568, 4.957586, 4.960464, 4.963702, 4.967002, 
    4.967633, 4.968585, 4.96942, 4.971097, 4.973547, 4.976954, 4.981276, 
    4.986701, 4.992226, 4.998084, 5.00092, 5.003414, 5.00525, 5.006023, 
    5.005275, 5.00252, 4.997281, 4.989166, 4.977938, 4.963619, 4.94656, 
    4.927482, 4.90745, 4.887774, 4.869849, 4.854956, 4.84411, 4.837931, 
    4.836633,
  // momentumX(21,20, 0-49)
    4.920373, 4.926408, 4.932198, 4.937615, 4.942574, 4.947017, 4.95092, 
    4.954266, 4.957061, 4.959322, 4.961086, 4.962402, 4.963344, 4.963996, 
    4.96446, 0, 4.958336, 4.959911, 4.962055, 4.964373, 4.966731, 4.965669, 
    4.965298, 4.965133, 4.966242, 4.968559, 4.972223, 4.977122, 4.983384, 
    4.989923, 4.997092, 5.000469, 5.003476, 5.005798, 5.007044, 5.006776, 
    5.004527, 4.999839, 4.992319, 4.981717, 4.96802, 4.951524, 4.932887, 
    4.913119, 4.893489, 4.875374, 4.860076, 4.848648, 4.841766, 4.839701,
  // momentumX(21,21, 0-49)
    4.922716, 4.928973, 4.934875, 4.9403, 4.945176, 4.949471, 4.95318, 
    4.956317, 4.958914, 4.96101, 4.962654, 4.963908, 4.964848, 4.965567, 
    4.966182, 0, 4.955145, 4.957202, 4.959885, 4.962759, 4.965636, 4.964164, 
    4.963536, 4.963161, 4.964198, 4.966575, 4.970424, 4.975614, 4.982278, 
    4.989311, 4.997245, 5.000715, 5.003937, 5.006592, 5.008276, 5.008539, 
    5.006902, 5.002893, 4.996096, 4.986228, 4.97323, 4.957343, 4.939162, 
    4.919639, 4.900001, 4.881614, 4.865797, 4.85364, 4.845881, 4.842846,
  // momentumX(21,22, 0-49)
    4.924577, 4.931123, 4.937216, 4.942735, 4.947618, 4.951845, 4.955435, 
    4.958422, 4.960857, 4.962803, 4.964324, 4.965492, 4.966395, 4.967139, 
    4.967857, 0, 4.952854, 4.955309, 4.958461, 4.96184, 4.965202, 4.963355, 
    4.962503, 4.961944, 4.962914, 4.96533, 4.96931, 4.974701, 4.981636, 
    4.988995, 4.997468, 5.000855, 5.004099, 5.006884, 5.008801, 5.009401, 
    5.008202, 5.004722, 4.998529, 4.989316, 4.976982, 4.961714, 4.944051, 
    4.92488, 4.905382, 4.886895, 4.870741, 4.858034, 4.849556, 4.845685,
  // momentumX(21,23, 0-49)
    4.925975, 4.932854, 4.939191, 4.944864, 4.949818, 4.954044, 4.957575, 
    4.960462, 4.962778, 4.964598, 4.966004, 4.967083, 4.967932, 4.968668, 
    4.969452, 0, 4.951511, 4.954235, 4.957705, 4.961428, 4.965119, 4.962908, 
    4.961822, 4.961064, 4.961936, 4.964339, 4.968385, 4.973899, 4.98101, 
    4.988581, 4.997424, 5.000678, 5.003872, 5.006702, 5.008762, 5.009603, 
    5.008744, 5.0057, 5.000029, 4.9914, 4.97968, 4.96501, 4.947873, 4.929098, 
    4.909818, 4.891339, 4.874972, 4.861847, 4.852779, 4.848183,
  // momentumX(21,24, 0-49)
    4.926955, 4.934186, 4.940796, 4.946662, 4.951729, 4.956, 4.959518, 
    4.962349, 4.964579, 4.966302, 4.96761, 4.968601, 4.969385, 4.970094, 
    4.970906, 0, 4.951337, 4.954191, 4.957818, 4.961719, 4.965586, 4.963124, 
    4.961879, 4.96099, 4.961792, 4.964177, 4.968248, 4.973822, 4.981027, 
    4.988714, 4.997774, 5.000921, 5.004061, 5.006891, 5.009009, 5.009973, 
    5.009304, 5.006517, 5.001168, 4.992916, 4.981607, 4.967354, 4.950599, 
    4.932136, 4.913054, 4.894632, 4.878164, 4.864782, 4.855316, 4.850201,
  // momentumX(21,25, 0-49)
    4.927581, 4.93516, 4.94205, 4.948121, 4.953326, 4.957671, 4.961206, 
    4.964014, 4.96619, 4.967835, 4.969058, 4.969966, 4.970678, 4.971337, 
    4.972132, 0, 4.951993, 4.954841, 4.958466, 4.962369, 4.966248, 4.963695, 
    4.962402, 4.961487, 4.962284, 4.964675, 4.968763, 4.974359, 4.981592, 
    4.989312, 4.998431, 5.001542, 5.004662, 5.007491, 5.009628, 5.010636, 
    5.010038, 5.007354, 5.002141, 4.994059, 4.982945, 4.968903, 4.952358, 
    4.934081, 4.915137, 4.896785, 4.880301, 4.866809, 4.857136, 4.851721,
  // momentumX(21,26, 0-49)
    4.927925, 4.935825, 4.942978, 4.949254, 4.954605, 4.959037, 4.962613, 
    4.965418, 4.967557, 4.969142, 4.970285, 4.971105, 4.971728, 4.972306, 
    4.973034, 0, 4.953425, 4.95613, 4.959591, 4.963326, 4.96705, 4.964577, 
    4.963362, 4.962536, 4.963402, 4.965837, 4.969944, 4.975535, 4.982742, 
    4.990416, 4.999442, 5.002605, 5.005761, 5.008602, 5.010732, 5.011711, 
    5.011069, 5.008329, 5.003057, 4.994917, 4.983764, 4.969701, 4.953165, 
    4.934923, 4.91604, 4.89776, 4.881342, 4.867894, 4.858222, 4.852753,
  // momentumX(21,27, 0-49)
    4.92806, 4.936237, 4.943624, 4.950087, 4.955577, 4.960105, 4.963733, 
    4.96655, 4.968665, 4.970191, 4.971249, 4.971961, 4.972464, 4.972912, 
    4.973501, 0, 4.955719, 4.958138, 4.961273, 4.964661, 4.968061, 4.965804, 
    4.964757, 4.964105, 4.965088, 4.967585, 4.971696, 4.977244, 4.98436, 
    4.99191, 5.000689, 5.003982, 5.007212, 5.01007, 5.012156, 5.013031, 
    5.01223, 5.009284, 5.00377, 4.995371, 4.983961, 4.969677, 4.952976, 
    4.93465, 4.915774, 4.897588, 4.881337, 4.868097, 4.85864, 4.853362,
  // momentumX(21,28, 0-49)
    4.928054, 4.936454, 4.944035, 4.950661, 4.956285, 4.960913, 4.964603, 
    4.967442, 4.969531, 4.970989, 4.971935, 4.972499, 4.972823, 4.973068, 
    4.973427, 0, 4.959241, 4.961226, 4.963868, 4.966732, 4.969642, 4.967668, 
    4.96682, 4.966366, 4.967466, 4.969997, 4.974066, 4.979512, 4.986459, 
    4.993795, 5.002191, 5.005653, 5.008963, 5.011804, 5.013775, 5.014439, 
    5.013337, 5.010012, 5.004061, 4.995199, 4.983335, 4.968651, 4.951647, 
    4.933157, 4.914279, 4.896254, 4.880302, 4.867464, 4.858457, 4.853627,
  // momentumX(21,29, 0-49)
    4.92797, 4.936532, 4.944271, 4.951048, 4.956806, 4.961545, 4.965309, 
    4.968172, 4.970227, 4.971584, 4.972364, 4.972703, 4.972755, 4.972694, 
    4.972711, 0, 4.963769, 4.965175, 4.967158, 4.969325, 4.971568, 4.96982, 
    4.969094, 4.968768, 4.969911, 4.972406, 4.976363, 4.981632, 4.988328, 
    4.995357, 5.003223, 5.006826, 5.010169, 5.01293, 5.014711, 5.015079, 
    5.013591, 5.0098, 5.003335, 4.99394, 4.981572, 4.966462, 4.949168, 
    4.930563, 4.911772, 4.894035, 4.878546, 4.866288, 4.85792, 4.853728,
  // momentumX(21,30, 0-49)
    4.926956, 4.934618, 4.941468, 4.947391, 4.952364, 4.956439, 4.959708, 
    4.962296, 4.964333, 4.965935, 4.967184, 4.968123, 4.968738, 4.968968, 
    4.968709, 4.975595, 4.962874, 4.964472, 4.967275, 4.970613, 4.974156, 
    4.97453, 4.975579, 4.976661, 4.978667, 4.98145, 4.985137, 4.989669, 
    4.995262, 5.000958, 5.007199, 5.009936, 5.012409, 5.014312, 5.015257, 
    5.014821, 5.012557, 5.008026, 5.000863, 4.990838, 4.977942, 4.962452, 
    4.944969, 4.926406, 4.9079, 4.890683, 4.875904, 4.864484, 4.857009, 
    4.853695,
  // momentumX(21,31, 0-49)
    4.926929, 4.934672, 4.941601, 4.947601, 4.95264, 4.956754, 4.960025, 
    4.962573, 4.964523, 4.965997, 4.967094, 4.96788, 4.968374, 4.968542, 
    4.968293, 4.975252, 4.964764, 4.96593, 4.968161, 4.970851, 4.97374, 
    4.974269, 4.975286, 4.976324, 4.978278, 4.981052, 4.98479, 4.98941, 
    4.995051, 5.0007, 5.006574, 5.009628, 5.012319, 5.014328, 5.015259, 
    5.014685, 5.012158, 5.007254, 4.999632, 4.989102, 4.975713, 4.959807, 
    4.942053, 4.923415, 4.905064, 4.888221, 4.874006, 4.863276, 4.856546, 
    4.853962,
  // momentumX(21,32, 0-49)
    4.926838, 4.934477, 4.941327, 4.947276, 4.952287, 4.956389, 4.959658, 
    4.962198, 4.964133, 4.965584, 4.966657, 4.967435, 4.967957, 4.968214, 
    4.968139, 4.974419, 4.966065, 4.966943, 4.968725, 4.970888, 4.973237, 
    4.974019, 4.975111, 4.976216, 4.978195, 4.980991, 4.984751, 4.989377, 
    4.994931, 5.000389, 5.005764, 5.009021, 5.011818, 5.013818, 5.014621, 
    5.013795, 5.0109, 5.005525, 4.997361, 4.986272, 4.972367, 4.956063, 
    4.938097, 4.919488, 4.901426, 4.885119, 4.871639, 4.861775, 4.855964, 
    4.854273,
  // momentumX(21,33, 0-49)
    4.926754, 4.934147, 4.940796, 4.946594, 4.951506, 4.955551, 4.958797, 
    4.961343, 4.963299, 4.964785, 4.96591, 4.966764, 4.967407, 4.967854, 
    4.968068, 4.973201, 4.966861, 4.967598, 4.969047, 4.970792, 4.972705, 
    4.973806, 4.97506, 4.976316, 4.978374, 4.981203, 4.984944, 4.989483, 
    4.994825, 4.999962, 5.004738, 5.008092, 5.010881, 5.012757, 5.013318, 
    5.012129, 5.00876, 5.002823, 4.994051, 4.982362, 4.967942, 4.951282, 
    4.93319, 4.914731, 4.897108, 4.881502, 4.868926, 4.86009, 4.855348, 
    4.854691,
  // momentumX(21,34, 0-49)
    4.926736, 4.933774, 4.940129, 4.945702, 4.950455, 4.954404, 4.95761, 
    4.960158, 4.962151, 4.9637, 4.964916, 4.96589, 4.966699, 4.967385, 
    4.967942, 4.971733, 4.967276, 4.967985, 4.969195, 4.970612, 4.972173, 
    4.973621, 4.975093, 4.976563, 4.978733, 4.98159, 4.98526, 4.989622, 
    4.994627, 4.999331, 5.003438, 5.006778, 5.009446, 5.011085, 5.011292, 
    5.009635, 5.005699, 4.999127, 4.989699, 4.977401, 4.962496, 4.945557, 
    4.927455, 4.909292, 4.892269, 4.877531, 4.866017, 4.858353, 4.854806, 
    4.855289,
  // momentumX(21,35, 0-49)
    4.926836, 4.933433, 4.939422, 4.944709, 4.949258, 4.953081, 4.956228, 
    4.95877, 4.960804, 4.96243, 4.96375, 4.964861, 4.965849, 4.966776, 
    4.967676, 4.970145, 4.967444, 4.968202, 4.969242, 4.970393, 4.971665, 
    4.973465, 4.975183, 4.976903, 4.979197, 4.982062, 4.985603, 4.989695, 
    4.994246, 4.998414, 5.001794, 5.005006, 5.007436, 5.008721, 5.008463, 
    5.00624, 5.001657, 4.994396, 4.984295, 4.971416, 4.9561, 4.938995, 
    4.921033, 4.903339, 4.887095, 4.873391, 4.863085, 4.856715, 4.854457, 
    4.856152,
  // momentumX(21,36, 0-49)
    4.927101, 4.933189, 4.938755, 4.943709, 4.948019, 4.951687, 4.954755, 
    4.957284, 4.959356, 4.961058, 4.962487, 4.963735, 4.964891, 4.966037, 
    4.967238, 4.96855, 4.967488, 4.968328, 4.969235, 4.970166, 4.9712, 
    4.973329, 4.975299, 4.977283, 4.979695, 4.982537, 4.985882, 4.989611, 
    4.993591, 4.997127, 4.999732, 5.00269, 5.004757, 5.005571, 5.00474, 
    5.00186, 4.996566, 4.988592, 4.977838, 4.964443, 4.948833, 4.931724, 
    4.91409, 4.897061, 4.881786, 4.869282, 4.860319, 4.855337, 4.85443, 
    4.857368,
  // momentumX(21,37, 0-49)
    4.927572, 4.933101, 4.938197, 4.942782, 4.946818, 4.950309, 4.95328, 
    4.955783, 4.957885, 4.959661, 4.961193, 4.962566, 4.963869, 4.965193, 
    4.966624, 4.967034, 4.967501, 4.96842, 4.969209, 4.969953, 4.970782, 
    4.9732, 4.975408, 4.97765, 4.980156, 4.982931, 4.986008, 4.989279, 
    4.992575, 4.995385, 4.997163, 4.999734, 5.00131, 5.001532, 5.000024, 
    4.996412, 4.990367, 4.981685, 4.970336, 4.956542, 4.940803, 4.923894, 
    4.906811, 4.890669, 4.876559, 4.865418, 4.857912, 4.854388, 4.854856, 
    4.859026,
  // momentumX(21,38, 0-49)
    4.928286, 4.933214, 4.937806, 4.941989, 4.945725, 4.949013, 4.951869, 
    4.954332, 4.956453, 4.95829, 4.959915, 4.9614, 4.962823, 4.964279, 
    4.965862, 4.965644, 4.967535, 4.968503, 4.969175, 4.969752, 4.970407, 
    4.97306, 4.975472, 4.977946, 4.980508, 4.983161, 4.985892, 4.988606, 
    4.991111, 4.993099, 4.993998, 4.996039, 4.99699, 4.996502, 4.994226, 
    4.989821, 4.983016, 4.97367, 4.961834, 4.947803, 4.932146, 4.915679, 
    4.899399, 4.884381, 4.87164, 4.86201, 4.856055, 4.854027, 4.85586, 
    4.861211,
  // momentumX(21,39, 0-49)
    4.929265, 4.933565, 4.937625, 4.941379, 4.944791, 4.947852, 4.950571, 
    4.952974, 4.955095, 4.95698, 4.958681, 4.960257, 4.961775, 4.963317, 
    4.964976, 4.964395, 4.967595, 4.96857, 4.969121, 4.969549, 4.97005, 
    4.972878, 4.975447, 4.978108, 4.980676, 4.983141, 4.985444, 4.987503, 
    4.989108, 4.990186, 4.990143, 4.991511, 4.991702, 4.990395, 4.987274, 
    4.982047, 4.974504, 4.964581, 4.952405, 4.938348, 4.923028, 4.907279, 
    4.892075, 4.878423, 4.867244, 4.859259, 4.854925, 4.8544, 4.857553, 
    4.863996,
  // momentumX(21,40, 0-49)
    4.930509, 4.934163, 4.937672, 4.940976, 4.944041, 4.946851, 4.949409, 
    4.951728, 4.953829, 4.95574, 4.957498, 4.959143, 4.96073, 4.962318, 
    4.963991, 4.96327, 4.967656, 4.968591, 4.969017, 4.969309, 4.969671, 
    4.972606, 4.975278, 4.97807, 4.980577, 4.982781, 4.984569, 4.985875, 
    4.986485, 4.986562, 4.985514, 4.986065, 4.985376, 4.983157, 4.979137, 
    4.973087, 4.964869, 4.954496, 4.942178, 4.928343, 4.913644, 4.898909, 
    4.885057, 4.873009, 4.86357, 4.857339, 4.854666, 4.855622, 4.860014, 
    4.867422,
  // momentumX(21,41, 0-49)
    4.931998, 4.934996, 4.937942, 4.94078, 4.943478, 4.946014, 4.948385, 
    4.950592, 4.952645, 4.954556, 4.956345, 4.958038, 4.959667, 4.961271, 
    4.962908, 4.962221, 4.967657, 4.968509, 4.968806, 4.968975, 4.969211, 
    4.972187, 4.974899, 4.977754, 4.980126, 4.981987, 4.983173, 4.983639, 
    4.983162, 4.982157, 4.980039, 4.979643, 4.977969, 4.974769, 4.969831, 
    4.962996, 4.954207, 4.943558, 4.931327, 4.917993, 4.904217, 4.890792, 
    4.878562, 4.868335, 4.860787, 4.856392, 4.855388, 4.857768, 4.863286, 
    4.8715,
  // momentumX(21,42, 0-49)
    4.933681, 4.93602, 4.938399, 4.940762, 4.943074, 4.945315, 4.947473, 
    4.949539, 4.951512, 4.953393, 4.955186, 4.9569, 4.958545, 4.960138, 
    4.961708, 4.961169, 4.967508, 4.968248, 4.968419, 4.968473, 4.968589, 
    4.971543, 4.97423, 4.977072, 4.979232, 4.980669, 4.981169, 4.980713, 
    4.979079, 4.976922, 4.973677, 4.972228, 4.969491, 4.965276, 4.95944, 
    4.951901, 4.942686, 4.931967, 4.920083, 4.907539, 4.894986, 4.883152, 
    4.872786, 4.864562, 4.859018, 4.856503, 4.857143, 4.860859, 4.867363, 
    4.876194,
  // momentumX(21,43, 0-49)
    4.935478, 4.937166, 4.938977, 4.940857, 4.942774, 4.9447, 4.946618, 
    4.948514, 4.950376, 4.952195, 4.953959, 4.955664, 4.957301, 4.958864, 
    4.960346, 4.960024, 4.967107, 4.967718, 4.967767, 4.967717, 4.967713, 
    4.970584, 4.973182, 4.975931, 4.977798, 4.978734, 4.978477, 4.977031, 
    4.974191, 4.970835, 4.966425, 4.963848, 4.960012, 4.95479, 4.948117, 
    4.939998, 4.930539, 4.919984, 4.908716, 4.897247, 4.886191, 4.876195, 
    4.867887, 4.861801, 4.858331, 4.857696, 4.859924, 4.86486, 4.87218, 
    4.88142,
  // momentumX(21,44, 0-49)
    4.937275, 4.938323, 4.939574, 4.940974, 4.942487, 4.944084, 4.945742, 
    4.947441, 4.949162, 4.950884, 4.95259, 4.954257, 4.955863, 4.957377, 
    4.958764, 4.958681, 4.966344, 4.966816, 4.966756, 4.966607, 4.966479, 
    4.969213, 4.971659, 4.974236, 4.975735, 4.976098, 4.975027, 4.972552, 
    4.968484, 4.96391, 4.958328, 4.954591, 4.949665, 4.943493, 4.936093, 
    4.927554, 4.91806, 4.907915, 4.897525, 4.887393, 4.878069, 4.8701, 
    4.863985, 4.860114, 4.858732, 4.859934, 4.863651, 4.869663, 4.877614, 
    4.887039,
  // momentumX(21,45, 0-49)
    4.938926, 4.939353, 4.940056, 4.940982, 4.942094, 4.943354, 4.944736, 
    4.946219, 4.947771, 4.949369, 4.950988, 4.952592, 4.954145, 4.955598, 
    4.956888, 4.957033, 4.965114, 4.965453, 4.965286, 4.965036, 4.964778, 
    4.967328, 4.969562, 4.97189, 4.972956, 4.972693, 4.970773, 4.967258, 
    4.961981, 4.956205, 4.949481, 4.944608, 4.938652, 4.931637, 4.923662, 
    4.914896, 4.905593, 4.896097, 4.886826, 4.878241, 4.870824, 4.865007, 
    4.861149, 4.859497, 4.860159, 4.863107, 4.868181, 4.875099, 4.883481, 
    4.892863,
  // momentumX(21,46, 0-49)
    4.940262, 4.940084, 4.940259, 4.940728, 4.941444, 4.942371, 4.943476, 
    4.944729, 4.946098, 4.947554, 4.949063, 4.950583, 4.952066, 4.953447, 
    4.954642, 4.95498, 4.963323, 4.963535, 4.963268, 4.96291, 4.962506, 
    4.964828, 4.9668, 4.968812, 4.969393, 4.968471, 4.965699, 4.961167, 
    4.954741, 4.947829, 4.940039, 4.934107, 4.927235, 4.919528, 4.911165, 
    4.902386, 4.893498, 4.884871, 4.876911, 4.870032, 4.864622, 4.861, 
    4.859388, 4.859892, 4.862491, 4.867044, 4.873307, 4.880941, 4.889546, 
    4.898666,
  // momentumX(21,47, 0-49)
    4.941096, 4.940332, 4.939998, 4.940029, 4.940372, 4.940979, 4.941815, 
    4.942842, 4.944026, 4.945332, 4.94672, 4.948144, 4.949549, 4.950854, 
    4.951961, 4.952435, 4.960899, 4.960996, 4.960621, 4.960141, 4.959572, 
    4.961631, 4.963296, 4.964937, 4.965001, 4.963412, 4.959817, 4.954334, 
    4.946867, 4.938931, 4.930195, 4.923338, 4.915718, 4.907512, 4.898972, 
    4.890397, 4.882132, 4.874554, 4.868045, 4.862955, 4.859578, 4.858113, 
    4.858655, 4.861183, 4.865554, 4.871528, 4.878778, 4.886925, 4.895541, 
    4.904192,
  // momentumX(21,48, 0-49)
    4.941243, 4.939906, 4.939085, 4.938703, 4.938699, 4.939013, 4.939602, 
    4.940422, 4.941435, 4.942599, 4.943874, 4.945204, 4.946529, 4.947761, 
    4.948786, 4.949333, 4.957789, 4.957774, 4.957283, 4.956659, 4.955901, 
    4.95767, 4.958993, 4.960226, 4.959764, 4.95753, 4.953178, 4.946849, 
    4.938492, 4.929691, 4.920184, 4.91259, 4.904428, 4.895942, 4.887444, 
    4.879278, 4.871814, 4.865419, 4.860435, 4.857142, 4.855741, 4.856319, 
    4.858856, 4.863209, 4.869135, 4.876301, 4.884318, 4.892757, 4.901187, 
    4.909195,
  // momentumX(21,49, 0-49)
    4.941844, 4.93949, 4.937799, 4.936679, 4.936049, 4.935833, 4.935967, 
    4.936391, 4.937048, 4.937884, 4.938838, 4.939832, 4.94078, 4.941552, 
    4.941981, 4.941836, 4.957452, 4.955976, 4.953788, 4.951624, 4.94955, 
    4.952877, 4.955788, 4.959049, 4.959525, 4.957204, 4.951482, 4.942688, 
    4.930685, 4.918662, 4.906098, 4.898111, 4.889776, 4.881432, 4.873471, 
    4.866293, 4.860284, 4.855782, 4.853061, 4.852297, 4.853556, 4.856781, 
    4.861804, 4.868344, 4.876037, 4.88445, 4.893135, 4.901632, 4.909525, 
    4.916467,
  // momentumX(22,0, 0-49)
    4.880537, 4.886049, 4.892055, 4.89834, 4.90474, 4.911143, 4.917471, 
    4.923685, 4.92976, 4.935697, 4.941501, 4.947173, 4.952713, 4.958113, 
    4.963342, 4.968148, 4.973527, 4.977929, 4.981947, 4.985516, 4.988526, 
    4.991129, 4.992905, 4.993828, 4.99375, 4.992583, 4.990228, 4.986621, 
    4.981689, 4.975449, 4.967793, 4.959002, 4.948776, 4.937156, 4.924249, 
    4.910238, 4.895406, 4.880136, 4.864914, 4.850298, 4.836879, 4.825234, 
    4.815861, 4.809134, 4.805259, 4.804258, 4.805966, 4.810053, 4.816054, 
    4.823408,
  // momentumX(22,1, 0-49)
    4.881404, 4.887128, 4.893311, 4.899741, 4.906262, 4.912758, 4.919157, 
    4.925417, 4.93152, 4.937462, 4.943248, 4.948881, 4.954358, 4.959669, 
    4.964782, 4.969224, 4.975, 4.979175, 4.982958, 4.986339, 4.989226, 
    4.992044, 4.994077, 4.995368, 4.995728, 4.995061, 4.993247, 4.99022, 
    4.985889, 4.980306, 4.973286, 4.96537, 4.95594, 4.94499, 4.932577, 
    4.918843, 4.904028, 4.888497, 4.872729, 4.857299, 4.842846, 4.830007, 
    4.819363, 4.81137, 4.806323, 4.804312, 4.805237, 4.808805, 4.814574, 
    4.821985,
  // momentumX(22,2, 0-49)
    4.882138, 4.888039, 4.894367, 4.900916, 4.907531, 4.914097, 4.920544, 
    4.926829, 4.932936, 4.938857, 4.944596, 4.950159, 4.955542, 4.960733, 
    4.965704, 4.969741, 4.975807, 4.979735, 4.983255, 4.986413, 4.989146, 
    4.992136, 4.994386, 4.996001, 4.99677, 4.996595, 4.995338, 4.992937, 
    4.989284, 4.984453, 4.978187, 4.971295, 4.962846, 4.952787, 4.941124, 
    4.927945, 4.913436, 4.897918, 4.881842, 4.865784, 4.850403, 4.836392, 
    4.824409, 4.815003, 4.808563, 4.805276, 4.805117, 4.807853, 4.813084, 
    4.820271,
  // momentumX(22,3, 0-49)
    4.88286, 4.888899, 4.895341, 4.901977, 4.908658, 4.915267, 4.921736, 
    4.92802, 4.9341, 4.93997, 4.945633, 4.951095, 4.956351, 4.961398, 
    4.966206, 4.969803, 4.976026, 4.979697, 4.982938, 4.98585, 4.988398, 
    4.991513, 4.99393, 4.995817, 4.996953, 4.997241, 4.996539, 4.994784, 
    4.991858, 4.987838, 4.982406, 4.976634, 4.969298, 4.960302, 4.949604, 
    4.937222, 4.923286, 4.908053, 4.891929, 4.875461, 4.859316, 4.844221, 
    4.830904, 4.820007, 4.812023, 4.807248, 4.80575, 4.807377, 4.811787, 
    4.818478,
  // momentumX(22,4, 0-49)
    4.883684, 4.889828, 4.896346, 4.903038, 4.90975, 4.916372, 4.922831, 
    4.929082, 4.935105, 4.940893, 4.946448, 4.951777, 4.956883, 4.96176, 
    4.966392, 4.969527, 4.975749, 4.97916, 4.982116, 4.984766, 4.987107, 
    4.990293, 4.992825, 4.99492, 4.996367, 4.997078, 4.996912, 4.995807, 
    4.993631, 4.990452, 4.985897, 4.981287, 4.975144, 4.96733, 4.957751, 
    4.94637, 4.93324, 4.918549, 4.902637, 4.886006, 4.869302, 4.853272, 
    4.838696, 4.826305, 4.8167, 4.810288, 4.807254, 4.807538, 4.810874, 
    4.816814,
  // momentumX(22,5, 0-49)
    4.884719, 4.890928, 4.897486, 4.904196, 4.910906, 4.917505, 4.92392, 
    4.930103, 4.936036, 4.941709, 4.947129, 4.952298, 4.957226, 4.961914, 
    4.96636, 4.969028, 4.97508, 4.978233, 4.980904, 4.983284, 4.985404, 
    4.98861, 4.991196, 4.993429, 4.995127, 4.99621, 4.996547, 4.996074, 
    4.994657, 4.992321, 4.988653, 4.985206, 4.980282, 4.973714, 4.96536, 
    4.955123, 4.942988, 4.929064, 4.913613, 4.897071, 4.880046, 4.86328, 
    4.847586, 4.833769, 4.822536, 4.814412, 4.809701, 4.80846, 4.81051, 
    4.815478,
  // momentumX(22,6, 0-49)
    4.886049, 4.892287, 4.898846, 4.905535, 4.912204, 4.918742, 4.925076, 
    4.931158, 4.936968, 4.942498, 4.947752, 4.952737, 4.957466, 4.961949, 
    4.9662, 4.968412, 4.974121, 4.97702, 4.979414, 4.981527, 4.983417, 
    4.986587, 4.98917, 4.991468, 4.99335, 4.994747, 4.995544, 4.99568, 
    4.995009, 4.993502, 4.990707, 4.988382, 4.984662, 4.979352, 4.972273, 
    4.963274, 4.952274, 4.9393, 4.924531, 4.908326, 4.89123, 4.873957, 
    4.857336, 4.842224, 4.829421, 4.819574, 4.813116, 4.810222, 4.810823, 
    4.814631,
  // momentumX(22,7, 0-49)
    4.887733, 4.893962, 4.900485, 4.907114, 4.913703, 4.920143, 4.92636, 
    4.932308, 4.937963, 4.94332, 4.948382, 4.953161, 4.957674, 4.961939, 
    4.965983, 4.967781, 4.972977, 4.975623, 4.977752, 4.979605, 4.981266, 
    4.984348, 4.986871, 4.989161, 4.991158, 4.992808, 4.994019, 4.994727, 
    4.994781, 4.994075, 4.992127, 4.990852, 4.98828, 4.984199, 4.978396, 
    4.970678, 4.960901, 4.949014, 4.935112, 4.919465, 4.902544, 4.885012, 
    4.867685, 4.851458, 4.837206, 4.825689, 4.817468, 4.812854, 4.811893, 
    4.814398,
  // momentumX(22,8, 0-49)
    4.88981, 4.895993, 4.902441, 4.908971, 4.915441, 4.921747, 4.927812, 
    4.933593, 4.939067, 4.944226, 4.949075, 4.953628, 4.957908, 4.96194, 
    4.965762, 4.967212, 4.971738, 4.974128, 4.976008, 4.977619, 4.979063, 
    4.982004, 4.98441, 4.986624, 4.988671, 4.990512, 4.992086, 4.993325, 
    4.994076, 4.994135, 4.992996, 4.992678, 4.991173, 4.988257, 4.983695, 
    4.977253, 4.968738, 4.958027, 4.945134, 4.930234, 4.913712, 4.896164, 
    4.878372, 4.86124, 4.845705, 4.832624, 4.822687, 4.816338, 4.813755, 
    4.814858,
  // momentumX(22,9, 0-49)
    4.892284, 4.898389, 4.904727, 4.911123, 4.917439, 4.923574, 4.929457, 
    4.935043, 4.94031, 4.945249, 4.949864, 4.954177, 4.958208, 4.96199, 
    4.965567, 4.966765, 4.970487, 4.972616, 4.974267, 4.975658, 4.976905, 
    4.979655, 4.981893, 4.983966, 4.986002, 4.987977, 4.989863, 4.991588, 
    4.993001, 4.993782, 4.993412, 4.993945, 4.993408, 4.991569, 4.988178, 
    4.982973, 4.975715, 4.966225, 4.954433, 4.940427, 4.924498, 4.90716, 
    4.889142, 4.871335, 4.854712, 4.84022, 4.828661, 4.820616, 4.8164, 
    4.816047,
  // momentumX(22,10, 0-49)
    4.895145, 4.901142, 4.907338, 4.913567, 4.919698, 4.925632, 4.931304, 
    4.93667, 4.941706, 4.946405, 4.950773, 4.95483, 4.958596, 4.96211, 
    4.965409, 4.96648, 4.969285, 4.971148, 4.972591, 4.973794, 4.974871, 
    4.977384, 4.979412, 4.981291, 4.983261, 4.985313, 4.987463, 4.989625, 
    4.991659, 4.993119, 4.993484, 4.99475, 4.995069, 4.994203, 4.991892, 
    4.987855, 4.981818, 4.973549, 4.96291, 4.949902, 4.93472, 4.917789, 
    4.899768, 4.881516, 4.864025, 4.8483, 4.835255, 4.825601, 4.819786, 
    4.817967,
  // momentumX(22,11, 0-49)
    4.898359, 4.904222, 4.910252, 4.916286, 4.922204, 4.927913, 4.93335, 
    4.938472, 4.943258, 4.947702, 4.951809, 4.955594, 4.959082, 4.962301, 
    4.965283, 4.966367, 4.968176, 4.969769, 4.971031, 4.972083, 4.973031, 
    4.975266, 4.977045, 4.978685, 4.980544, 4.98263, 4.984991, 4.987542, 
    4.990149, 4.992247, 4.993314, 4.995196, 4.996253, 4.996246, 4.994911, 
    4.991952, 4.987071, 4.979993, 4.970516, 4.958566, 4.944244, 4.927882, 
    4.910058, 4.891582, 4.873441, 4.856687, 4.842321, 4.831179, 4.823837, 
    4.82058,
  // momentumX(22,12, 0-49)
    4.901878, 4.907592, 4.913434, 4.919252, 4.924936, 4.930398, 4.935579, 
    4.940441, 4.944962, 4.949134, 4.952963, 4.956466, 4.959656, 4.962557, 
    4.965181, 4.966418, 4.967177, 4.968506, 4.96962, 4.970567, 4.97143, 
    4.973352, 4.974858, 4.976231, 4.977943, 4.980022, 4.98255, 4.985436, 
    4.988568, 4.991255, 4.992997, 4.995377, 4.997054, 4.99779, 4.997318, 
    4.995336, 4.991525, 4.98558, 4.977245, 4.966374, 4.952986, 4.937315, 
    4.919857, 4.901359, 4.882782, 4.865209, 4.849709, 4.837227, 4.828466, 
    4.823829,
  // momentumX(22,13, 0-49)
    4.90565, 4.911202, 4.916841, 4.922431, 4.927863, 4.933063, 4.937972, 
    4.942556, 4.946795, 4.950685, 4.954226, 4.957429, 4.960305, 4.962861, 
    4.96509, 4.966601, 4.96628, 4.967366, 4.968375, 4.969272, 4.970106, 
    4.971691, 4.97291, 4.973999, 4.975545, 4.977583, 4.980232, 4.9834, 
    4.986999, 4.990225, 4.992621, 4.995386, 4.997564, 4.998925, 4.999202, 
    4.998087, 4.99525, 4.990359, 4.983118, 4.973319, 4.960899, 4.946009, 
    4.92905, 4.910706, 4.891897, 4.873711, 4.857275, 4.843622, 4.83357, 
    4.827637,
  // momentumX(22,14, 0-49)
    4.909611, 4.915001, 4.920432, 4.925782, 4.930954, 4.935875, 4.940499, 
    4.944792, 4.948737, 4.952328, 4.955569, 4.958461, 4.961009, 4.963201, 
    4.965012, 4.966866, 4.965448, 4.966335, 4.967295, 4.968207, 4.969079, 
    4.970313, 4.971245, 4.97205, 4.973421, 4.975398, 4.978127, 4.981521, 
    4.985519, 4.989235, 4.992261, 4.995299, 4.997867, 4.999737, 5.000646, 
    5.000288, 4.998318, 4.994392, 4.988178, 4.979414, 4.96797, 4.953912, 
    4.937561, 4.919518, 4.900659, 4.882061, 4.864886, 4.850241, 4.839045, 
    4.831921,
  // momentumX(22,15, 0-49)
    4.913706, 4.918937, 4.924161, 4.929266, 4.934164, 4.938797, 4.943122, 
    4.947111, 4.950749, 4.954034, 4.956963, 4.959537, 4.961747, 4.96357, 
    4.964959, 4.967154, 4.964622, 4.965373, 4.966358, 4.967362, 4.968349, 
    4.96923, 4.969894, 4.970437, 4.971638, 4.973541, 4.976313, 4.979875, 
    4.984203, 4.988347, 4.99198, 4.995186, 4.998031, 5.000298, 5.001725, 
    5.002008, 5.000802, 4.997742, 4.992472, 4.984691, 4.974206, 4.96101, 
    4.945339, 4.927721, 4.908974, 4.89015, 4.87243, 4.856977, 4.844789, 
    4.836594,
  // momentumX(22,16, 0-49)
    4.917878, 4.922956, 4.927972, 4.932827, 4.937447, 4.94178, 4.945793, 
    4.949466, 4.952789, 4.95576, 4.958376, 4.960632, 4.962512, 4.963979, 
    4.964971, 4.967404, 4.963717, 4.964427, 4.965526, 4.966713, 4.967906, 
    4.968447, 4.96888, 4.969199, 4.970256, 4.972084, 4.974867, 4.978536, 
    4.983116, 4.987617, 4.991826, 4.995096, 4.998113, 5.000667, 5.002501, 
    5.003314, 5.00276, 5.000465, 4.996054, 4.989187, 4.979626, 4.967295, 
    4.952357, 4.935261, 4.916767, 4.897888, 4.879806, 4.863722, 4.850706, 
    4.841565,
  // momentumX(22,17, 0-49)
    4.92207, 4.926999, 4.931807, 4.936404, 4.940733, 4.944755, 4.948444, 
    4.951794, 4.9548, 4.957461, 4.959776, 4.961733, 4.963308, 4.964456, 
    4.965109, 4.967572, 4.962652, 4.963425, 4.964743, 4.966219, 4.967717, 
    4.967952, 4.96821, 4.968366, 4.96932, 4.971087, 4.973859, 4.977577, 
    4.982324, 4.9871, 4.991838, 4.99507, 4.998154, 5.000888, 5.00302, 
    5.004251, 5.00424, 5.002608, 4.998962, 4.992938, 4.984252, 4.972774, 
    4.9586, 4.942105, 4.923982, 4.905201, 4.886931, 4.870391, 4.856705, 
    4.846749,
  // momentumX(22,18, 0-49)
    4.926219, 4.930993, 4.935577, 4.939902, 4.943923, 4.94762, 4.950982, 
    4.954012, 4.956714, 4.95909, 4.961139, 4.96284, 4.964164, 4.96506, 
    4.965462, 4.967654, 4.961352, 4.962304, 4.963949, 4.965824, 4.967738, 
    4.967719, 4.967881, 4.967954, 4.96887, 4.970606, 4.973351, 4.977064, 
    4.981887, 4.986845, 4.99204, 4.995138, 4.998181, 5.000986, 5.003305, 
    5.004848, 5.005273, 5.004199, 5.001225, 4.995965, 4.988102, 4.977455, 
    4.964059, 4.948224, 4.930574, 4.912029, 4.893728, 4.876899, 4.862697, 
    4.852058,
  // momentumX(22,19, 0-49)
    4.930254, 4.934838, 4.939164, 4.943184, 4.946876, 4.950236, 4.953277, 
    4.95601, 4.958449, 4.960598, 4.962448, 4.963972, 4.965132, 4.96587, 
    4.966131, 4.967701, 4.959782, 4.961017, 4.963089, 4.965472, 4.967917, 
    4.967721, 4.967884, 4.967977, 4.968936, 4.970692, 4.973415, 4.977076, 
    4.981885, 4.986914, 4.992465, 4.995318, 4.998209, 5.000971, 5.003365, 
    5.005108, 5.005862, 5.005246, 5.002851, 4.998276, 4.991178, 4.981333, 
    4.968722, 4.953592, 4.936501, 4.918311, 4.900126, 4.883163, 4.868595, 
    4.857404,
  // momentumX(22,20, 0-49)
    4.935121, 4.940522, 4.945562, 4.95019, 4.954374, 4.958099, 4.961357, 
    4.964148, 4.966482, 4.968373, 4.969851, 4.970959, 4.971753, 4.972302, 
    4.972693, 0, 4.959976, 4.961293, 4.963098, 4.965001, 4.966878, 4.965349, 
    4.964415, 4.963618, 4.964009, 4.965533, 4.968349, 4.972388, 4.97783, 
    4.983681, 4.990357, 4.993667, 4.997002, 5.000195, 5.003012, 5.00518, 
    5.006382, 5.006256, 5.004407, 5.000442, 4.994011, 4.984875, 4.972975, 
    4.958509, 4.941978, 4.924188, 4.906198, 4.8892, 4.874375, 4.862727,
  // momentumX(22,21, 0-49)
    4.939007, 4.944368, 4.949268, 4.953667, 4.957558, 4.960947, 4.963851, 
    4.966298, 4.968316, 4.969938, 4.971203, 4.972163, 4.972878, 4.973427, 
    4.973916, 0, 4.955731, 4.957488, 4.959795, 4.962227, 4.964609, 4.962763, 
    4.96166, 4.960739, 4.961128, 4.962759, 4.965786, 4.970114, 4.975934, 
    4.982237, 4.989596, 4.992975, 4.996485, 4.999949, 5.003128, 5.00574, 
    5.007459, 5.007914, 5.006705, 5.003426, 4.997713, 4.989299, 4.978093, 
    4.964244, 4.948203, 4.930723, 4.912822, 4.895671, 4.880454, 4.868197,
  // momentumX(22,22, 0-49)
    4.942727, 4.948107, 4.952914, 4.957129, 4.960762, 4.96384, 4.966405, 
    4.968505, 4.970191, 4.971513, 4.972527, 4.973292, 4.973882, 4.974389, 
    4.974936, 0, 4.952352, 4.954473, 4.957218, 4.960129, 4.962974, 4.960836, 
    4.959574, 4.958531, 4.958904, 4.960607, 4.963778, 4.968307, 4.974384, 
    4.980988, 4.988835, 4.992147, 4.995678, 4.999262, 5.002652, 5.005566, 
    5.007674, 5.008605, 5.007951, 5.005296, 5.000262, 4.99256, 4.982064, 
    4.968881, 4.953407, 4.936348, 4.918674, 4.901524, 4.886073, 4.873363,
  // momentumX(22,23, 0-49)
    4.946211, 4.951646, 4.956401, 4.960465, 4.963868, 4.966659, 4.968901, 
    4.970664, 4.972017, 4.973031, 4.973774, 4.974321, 4.974754, 4.975182, 
    4.975747, 0, 4.949856, 4.952229, 4.955276, 4.958517, 4.961682, 4.959258, 
    4.957822, 4.956636, 4.956953, 4.958671, 4.961921, 4.966574, 4.97282, 
    4.979625, 4.98781, 4.991016, 4.994521, 4.998165, 5.001703, 5.004858, 
    5.007296, 5.008648, 5.0085, 5.006428, 5.002038, 4.995022, 4.98522, 
    4.972703, 4.957818, 4.94122, 4.923836, 4.906774, 4.891189, 4.878129,
  // momentumX(22,24, 0-49)
    4.949394, 4.954908, 4.959633, 4.963575, 4.966775, 4.969305, 4.971246, 
    4.972689, 4.973722, 4.97443, 4.9749, 4.975216, 4.975473, 4.975791, 
    4.976331, 0, 4.948518, 4.951012, 4.954212, 4.957628, 4.960968, 4.958356, 
    4.95681, 4.955535, 4.955814, 4.957535, 4.960822, 4.965538, 4.971878, 
    4.978793, 4.987182, 4.990316, 4.993803, 4.997482, 5.001118, 5.004433, 
    5.007102, 5.008749, 5.008963, 5.007317, 5.003409, 4.996915, 4.987658, 
    4.975676, 4.961286, 4.945103, 4.928017, 4.911108, 4.895511, 4.882263,
  // momentumX(22,25, 0-49)
    4.952204, 4.957809, 4.962523, 4.966364, 4.969392, 4.971691, 4.973362, 
    4.97451, 4.975244, 4.975662, 4.975863, 4.975944, 4.97601, 4.976191, 
    4.976657, 0, 4.948055, 4.950538, 4.953739, 4.957167, 4.960527, 4.957858, 
    4.956294, 4.955017, 4.955307, 4.957049, 4.960361, 4.965107, 4.971481, 
    4.978438, 4.986895, 4.990032, 4.993546, 4.99728, 5.001002, 5.004436, 
    5.00726, 5.0091, 5.009548, 5.008173, 5.004572, 4.998418, 4.989519, 
    4.977905, 4.96387, 4.948008, 4.931185, 4.914455, 4.898934, 4.885649,
  // momentumX(22,26, 0-49)
    4.95458, 4.960278, 4.964995, 4.96876, 4.971643, 4.973747, 4.975185, 
    4.976077, 4.97654, 4.97669, 4.976631, 4.976472, 4.976333, 4.976344, 
    4.976682, 0, 4.948453, 4.950796, 4.953845, 4.957116, 4.960338, 4.957754, 
    4.956271, 4.955087, 4.95545, 4.95724, 4.960577, 4.965328, 4.97169, 
    4.978623, 4.98702, 4.990255, 4.993862, 4.997688, 5.001496, 5.005016, 
    5.007926, 5.009855, 5.010394, 5.00912, 5.00563, 4.999599, 4.990843, 
    4.979391, 4.965537, 4.949868, 4.933245, 4.916705, 4.901348, 4.888179,
  // momentumX(22,27, 0-49)
    4.95647, 4.962255, 4.966988, 4.970704, 4.973483, 4.975435, 4.976684, 
    4.977357, 4.977584, 4.977483, 4.977173, 4.976769, 4.976398, 4.976196, 
    4.976342, 0, 4.94983, 4.951895, 4.954633, 4.957582, 4.960505, 4.958111, 
    4.956778, 4.955749, 4.956214, 4.95806, 4.961405, 4.966125, 4.972418, 
    4.979264, 4.98748, 4.990894, 4.994651, 4.998594, 5.002487, 5.006057, 
    5.008984, 5.010896, 5.011392, 5.010053, 5.006485, 5.000376, 4.991556, 
    4.98007, 4.96623, 4.950636, 4.934154, 4.917815, 4.902705, 4.889807,
  // momentumX(22,28, 0-49)
    4.957836, 4.963705, 4.968472, 4.972172, 4.974893, 4.976745, 4.977857, 
    4.978356, 4.978376, 4.978041, 4.977476, 4.976804, 4.976159, 4.975689, 
    4.975567, 0, 4.952566, 4.954219, 4.956491, 4.958948, 4.961411, 4.95925, 
    4.958077, 4.957208, 4.95776, 4.959622, 4.962923, 4.967553, 4.973707, 
    4.980392, 4.988312, 4.991958, 4.995893, 4.999952, 5.003895, 5.00745, 
    5.010296, 5.012068, 5.012367, 5.010787, 5.006949, 5.000559, 4.991478, 
    4.979781, 4.965812, 4.950198, 4.933821, 4.917719, 4.90296, 4.890495,
  // momentumX(22,29, 0-49)
    4.95867, 4.964626, 4.969453, 4.973186, 4.975905, 4.977718, 4.978745, 
    4.979113, 4.978947, 4.978374, 4.97753, 4.976545, 4.975567, 4.974751, 
    4.974271, 0, 4.95646, 4.95757, 4.959221, 4.961021, 4.962852, 4.960859, 
    4.959756, 4.958962, 4.95951, 4.961305, 4.96448, 4.968947, 4.974889, 
    4.981332, 4.988841, 4.992712, 4.996807, 5.000953, 5.004909, 5.008403, 
    5.011117, 5.012687, 5.012722, 5.010827, 5.006638, 4.999887, 4.990465, 
    4.978487, 4.964337, 4.94868, 4.932421, 4.916602, 4.902275, 4.890357,
  // momentumX(22,30, 0-49)
    4.958047, 4.963116, 4.967086, 4.970015, 4.972012, 4.973216, 4.973781, 
    4.973852, 4.973566, 4.973029, 4.972315, 4.97146, 4.970461, 4.969284, 
    4.96787, 4.971422, 4.957416, 4.958146, 4.959991, 4.962359, 4.964968, 
    4.964603, 4.964927, 4.965328, 4.966667, 4.968801, 4.971864, 4.975824, 
    4.980929, 4.98633, 4.992523, 4.995769, 4.999239, 5.002778, 5.006158, 
    5.009108, 5.011305, 5.01238, 5.011932, 5.009561, 5.00491, 4.997726, 
    4.987928, 4.975666, 4.961368, 4.945735, 4.929695, 4.914293, 4.900559, 
    4.889373,
  // momentumX(22,31, 0-49)
    4.95789, 4.963067, 4.967144, 4.970172, 4.972244, 4.973488, 4.974046, 
    4.974065, 4.973676, 4.972998, 4.972118, 4.97109, 4.969933, 4.968622, 
    4.967101, 4.971066, 4.959039, 4.959276, 4.960526, 4.96225, 4.964221, 
    4.963971, 4.964255, 4.964615, 4.965906, 4.968037, 4.971161, 4.975234, 
    4.980437, 4.98588, 4.991862, 4.995546, 4.999402, 5.003253, 5.00686, 
    5.009934, 5.012142, 5.013105, 5.012422, 5.009698, 5.004597, 4.9969, 
    4.986571, 4.973823, 4.959142, 4.94329, 4.927226, 4.912013, 4.898664, 
    4.888015,
  // momentumX(22,32, 0-49)
    4.957166, 4.962335, 4.966437, 4.969514, 4.971652, 4.972965, 4.973582, 
    4.97364, 4.973271, 4.972588, 4.971687, 4.970632, 4.969455, 4.968151, 
    4.96666, 4.970359, 4.96031, 4.960156, 4.960892, 4.962051, 4.963462, 
    4.963401, 4.963728, 4.964138, 4.96545, 4.967617, 4.970803, 4.974948, 
    4.980169, 4.985564, 4.991252, 4.995315, 4.999488, 5.003579, 5.007331, 
    5.010444, 5.012566, 5.013313, 5.012284, 5.009094, 5.003433, 4.995127, 
    4.984194, 4.970913, 4.955841, 4.939794, 4.923772, 4.908843, 4.895998, 
    4.886026,
  // momentumX(22,33, 0-49)
    4.955983, 4.961055, 4.965122, 4.968218, 4.970413, 4.971811, 4.972531, 
    4.972694, 4.972424, 4.971832, 4.971011, 4.970033, 4.968942, 4.967745, 
    4.966402, 4.969375, 4.961257, 4.960827, 4.96114, 4.961818, 4.962752, 
    4.962927, 4.963367, 4.963902, 4.965289, 4.967519, 4.970751, 4.974916, 
    4.980073, 4.985337, 4.990673, 4.995048, 4.999469, 5.003721, 5.007534, 
    5.010592, 5.01253, 5.012957, 5.011473, 5.007711, 5.001394, 4.992397, 
    4.980807, 4.966975, 4.951529, 4.935343, 4.919448, 4.904913, 4.892695, 
    4.883534,
  // momentumX(22,34, 0-49)
    4.954448, 4.95936, 4.963346, 4.966434, 4.968682, 4.970178, 4.971027, 
    4.971339, 4.971222, 4.970782, 4.970108, 4.969277, 4.968343, 4.967324, 
    4.966204, 4.968204, 4.961935, 4.961338, 4.961315, 4.96159, 4.962114, 
    4.962554, 4.963157, 4.963874, 4.965377, 4.967681, 4.970933, 4.975061, 
    4.980067, 4.985126, 4.99007, 4.994689, 4.999281, 5.003613, 5.007399, 
    5.010306, 5.01196, 5.011963, 5.009924, 5.005498, 4.998452, 4.988713, 
    4.976445, 4.962076, 4.946308, 4.930067, 4.914408, 4.900389, 4.888928, 
    4.880701,
  // momentumX(22,35, 0-49)
    4.952672, 4.957375, 4.961246, 4.964301, 4.966592, 4.968191, 4.969186, 
    4.969673, 4.969746, 4.969497, 4.969015, 4.968374, 4.967635, 4.966836, 
    4.965979, 4.966949, 4.962429, 4.961751, 4.961463, 4.961401, 4.961579, 
    4.962293, 4.96309, 4.964033, 4.965674, 4.968048, 4.971286, 4.975313, 
    4.980082, 4.984866, 4.989388, 4.994173, 4.99885, 5.00317, 5.006832, 
    5.00949, 5.010759, 5.010242, 5.00756, 5.002398, 4.994569, 4.984073, 
    4.971148, 4.9563, 4.940302, 4.924123, 4.908833, 4.895466, 4.88489, 
    4.877709,
  // momentumX(22,36, 0-49)
    4.950771, 4.955221, 4.958945, 4.961947, 4.96427, 4.965969, 4.967115, 
    4.96779, 4.968071, 4.968041, 4.967778, 4.967352, 4.96683, 4.966259, 
    4.965673, 4.965696, 4.962821, 4.962123, 4.961627, 4.961285, 4.961173, 
    4.96215, 4.963158, 4.96435, 4.96614, 4.968571, 4.97175, 4.975606, 
    4.980051, 4.984489, 4.988561, 4.993416, 4.99808, 5.002285, 5.005719, 
    5.008024, 5.008811, 5.007683, 5.004285, 4.998341, 4.98972, 4.978488, 
    4.96497, 4.949749, 4.933655, 4.917694, 4.902929, 4.890361, 4.880794, 
    4.874759,
  // momentumX(22,37, 0-49)
    4.948856, 4.953017, 4.956562, 4.959488, 4.961827, 4.963615, 4.964911, 
    4.965777, 4.966276, 4.966475, 4.966443, 4.966245, 4.965945, 4.9656, 
    4.965266, 4.964514, 4.963181, 4.962499, 4.961835, 4.961262, 4.960908, 
    4.962128, 4.963348, 4.964801, 4.966734, 4.969196, 4.972267, 4.975879, 
    4.979912, 4.983932, 4.987516, 4.992332, 4.996866, 5.000842, 5.003934, 
    5.005777, 5.005983, 5.004169, 5.000006, 4.993264, 4.983874, 4.971982, 
    4.957987, 4.942545, 4.926535, 4.910977, 4.896918, 4.885301, 4.876864, 
    4.872054,
  // momentumX(22,38, 0-49)
    4.947029, 4.95087, 4.954208, 4.957035, 4.959365, 4.961228, 4.962661, 
    4.96371, 4.964424, 4.964855, 4.965057, 4.965089, 4.965008, 4.964876, 
    4.964758, 4.963451, 4.963553, 4.962902, 4.962105, 4.961343, 4.960793, 
    4.962229, 4.963652, 4.965358, 4.967416, 4.969876, 4.972776, 4.976065, 
    4.979594, 4.983118, 4.98617, 4.990817, 4.995093, 4.99871, 5.00134, 
    5.002613, 5.00215, 4.999588, 4.994634, 4.987115, 4.977029, 4.964597, 
    4.950294, 4.934833, 4.919126, 4.904189, 4.891028, 4.880522, 4.873323, 
    4.869796,
  // momentumX(22,39, 0-49)
    4.945388, 4.948878, 4.95198, 4.954679, 4.956977, 4.958889, 4.960439, 
    4.961655, 4.962572, 4.963227, 4.96366, 4.963917, 4.964046, 4.964107, 
    4.964168, 4.96253, 4.963966, 4.963343, 4.962438, 4.96153, 4.960828, 
    4.962446, 4.964049, 4.965991, 4.968144, 4.970555, 4.973221, 4.976102, 
    4.979031, 4.981975, 4.984433, 4.988768, 4.992643, 4.995764, 4.997804, 
    4.9984, 4.997189, 4.993839, 4.988104, 4.979869, 4.969203, 4.956405, 
    4.94201, 4.926777, 4.911627, 4.89755, 4.885493, 4.876248, 4.870383, 
    4.868177,
  // momentumX(22,40, 0-49)
    4.944005, 4.947119, 4.949958, 4.952499, 4.954735, 4.956668, 4.958309, 
    4.959668, 4.960769, 4.96163, 4.962281, 4.962752, 4.96308, 4.963314, 
    4.963518, 4.961757, 4.964414, 4.963816, 4.962826, 4.961812, 4.960998, 
    4.962762, 4.964519, 4.966666, 4.968871, 4.971179, 4.973535, 4.975921, 
    4.978155, 4.980425, 4.982213, 4.986079, 4.989399, 4.99188, 4.993204, 
    4.993023, 4.991001, 4.986851, 4.980374, 4.971526, 4.960449, 4.947505, 
    4.933281, 4.918559, 4.904246, 4.891278, 4.880527, 4.87269, 4.868237, 
    4.867364,
  // momentumX(22,41, 0-49)
    4.942934, 4.945651, 4.948199, 4.950552, 4.952695, 4.954617, 4.956311, 
    4.957786, 4.959041, 4.960086, 4.960935, 4.961604, 4.962116, 4.962505, 
    4.962822, 4.961109, 4.964873, 4.964289, 4.963243, 4.96216, 4.961271, 
    4.963148, 4.965024, 4.967335, 4.969543, 4.971682, 4.973652, 4.975451, 
    4.976894, 4.978395, 4.979421, 4.98265, 4.985257, 4.986954, 4.987439, 
    4.986394, 4.983522, 4.978585, 4.971448, 4.962138, 4.950858, 4.938031, 
    4.924275, 4.910371, 4.897185, 4.885581, 4.876331, 4.870027, 4.86704, 
    4.867486,
  // momentumX(22,42, 0-49)
    4.942198, 4.944501, 4.946737, 4.948874, 4.950887, 4.952759, 4.954475, 
    4.956024, 4.957401, 4.9586, 4.959621, 4.960468, 4.961146, 4.961676, 
    4.962083, 4.960546, 4.965296, 4.964724, 4.963648, 4.962533, 4.961604, 
    4.963559, 4.96552, 4.967943, 4.970094, 4.971998, 4.973501, 4.974625, 
    4.975183, 4.975811, 4.975973, 4.978401, 4.980134, 4.980906, 4.980445, 
    4.978471, 4.974735, 4.969062, 4.961384, 4.951796, 4.940564, 4.928149, 
    4.91518, 4.90241, 4.890639, 4.880638, 4.873065, 4.868399, 4.866908, 
    4.868633,
  // momentumX(22,43, 0-49)
    4.941798, 4.943673, 4.945574, 4.947466, 4.949317, 4.951102, 4.952796, 
    4.954382, 4.95584, 4.957156, 4.958319, 4.959318, 4.960145, 4.9608, 
    4.961287, 4.960012, 4.965619, 4.965061, 4.963984, 4.962872, 4.961929, 
    4.963934, 4.965942, 4.968421, 4.970454, 4.972047, 4.973005, 4.973367, 
    4.972955, 4.97261, 4.971803, 4.973268, 4.973981, 4.973707, 4.972209, 
    4.969264, 4.964683, 4.958358, 4.950296, 4.940651, 4.929743, 4.918052, 
    4.906193, 4.894865, 4.884781, 4.876598, 4.870849, 4.867894, 4.867904, 
    4.870842,
  // momentumX(22,44, 0-49)
    4.941687, 4.943127, 4.944678, 4.9463, 4.947957, 4.949617, 4.95125, 
    4.952827, 4.954327, 4.955722, 4.956991, 4.958113, 4.959068, 4.959835, 
    4.960393, 4.959428, 4.965758, 4.965227, 4.96418, 4.963101, 4.962169, 
    4.964197, 4.966213, 4.968689, 4.970536, 4.971749, 4.972087, 4.97161, 
    4.970154, 4.968743, 4.966866, 4.967227, 4.966793, 4.965372, 4.962781, 
    4.958857, 4.953483, 4.946626, 4.938364, 4.928908, 4.918612, 4.907955, 
    4.897513, 4.88791, 4.87975, 4.87356, 4.869744, 4.868541, 4.870022, 
    4.874084,
  // momentumX(22,45, 0-49)
    4.941793, 4.942795, 4.943985, 4.945317, 4.946753, 4.948253, 4.949785, 
    4.951314, 4.952811, 4.954244, 4.955584, 4.9568, 4.957859, 4.958724, 
    4.959352, 4.958708, 4.965632, 4.96514, 4.964149, 4.963128, 4.962224, 
    4.964252, 4.966239, 4.96865, 4.97025, 4.971015, 4.97067, 4.969294, 
    4.966736, 4.964185, 4.961152, 4.960292, 4.958618, 4.955986, 4.952279, 
    4.947404, 4.941326, 4.934086, 4.92583, 4.916817, 4.907412, 4.898078, 
    4.889328, 4.881688, 4.875639, 4.87157, 4.869749, 4.870298, 4.873192, 
    4.878266,
  // momentumX(22,46, 0-49)
    4.942007, 4.942574, 4.943394, 4.944422, 4.945613, 4.946927, 4.948323, 
    4.949766, 4.951222, 4.952654, 4.954029, 4.955307, 4.956448, 4.957397, 
    4.958094, 4.957758, 4.965144, 4.964711, 4.963798, 4.962851, 4.961987, 
    4.963995, 4.965917, 4.968205, 4.969499, 4.96976, 4.968681, 4.966363, 
    4.962676, 4.958935, 4.954689, 4.952533, 4.949564, 4.9457, 4.940897, 
    4.935141, 4.928477, 4.921025, 4.91299, 4.904661, 4.896404, 4.888639, 
    4.881803, 4.876304, 4.87249, 4.870608, 4.870795, 4.873055, 4.877275, 
    4.88323,
  // momentumX(22,47, 0-49)
    4.942184, 4.942324, 4.942777, 4.943493, 4.944427, 4.94553, 4.946764, 
    4.948091, 4.949472, 4.950871, 4.952249, 4.95356, 4.954759, 4.955781, 
    4.956546, 4.956481, 4.964205, 4.963849, 4.963029, 4.962167, 4.961345, 
    4.963313, 4.965137, 4.967248, 4.968189, 4.967905, 4.966066, 4.96279, 
    4.957972, 4.953028, 4.947546, 4.944068, 4.939801, 4.934735, 4.928899, 
    4.922368, 4.915265, 4.907782, 4.900171, 4.892743, 4.885846, 4.879838, 
    4.875064, 4.87181, 4.870286, 4.870596, 4.872749, 4.876638, 4.882066, 
    4.888757,
  // momentumX(22,48, 0-49)
    4.942157, 4.941879, 4.941971, 4.942379, 4.943048, 4.943933, 4.94499, 
    4.94618, 4.947465, 4.948805, 4.95016, 4.951481, 4.952719, 4.953801, 
    4.954633, 4.95479, 4.962732, 4.962471, 4.961751, 4.960971, 4.960187, 
    4.962099, 4.963796, 4.965682, 4.966233, 4.965381, 4.962782, 4.958564, 
    4.952653, 4.946531, 4.939835, 4.935065, 4.929556, 4.923367, 4.916611, 
    4.909441, 4.902061, 4.894722, 4.887719, 4.881363, 4.875974, 4.871838, 
    4.869196, 4.86821, 4.868954, 4.871396, 4.875418, 4.880815, 4.887309, 
    4.894578,
  // momentumX(22,49, 0-49)
    4.942302, 4.941273, 4.940712, 4.94055, 4.940726, 4.94118, 4.941866, 
    4.942734, 4.943739, 4.944835, 4.945973, 4.947086, 4.948108, 4.94893, 
    4.949424, 4.949001, 4.964243, 4.962885, 4.960816, 4.958843, 4.957083, 
    4.960893, 4.964464, 4.968607, 4.970275, 4.969415, 4.9654, 4.958524, 
    4.948629, 4.938767, 4.928291, 4.922237, 4.915466, 4.908151, 4.900531, 
    4.892879, 4.885505, 4.878732, 4.872895, 4.868293, 4.865188, 4.863756, 
    4.864096, 4.866197, 4.869948, 4.875145, 4.881518, 4.888731, 4.896425, 
    4.904231,
  // momentumX(23,0, 0-49)
    4.895426, 4.901486, 4.90759, 4.913628, 4.919533, 4.92527, 4.930825, 
    4.936199, 4.941404, 4.946454, 4.951359, 4.956124, 4.960742, 4.965197, 
    4.969453, 4.973246, 4.977482, 4.980842, 4.983828, 4.986425, 4.988595, 
    4.990544, 4.991959, 4.992893, 4.993297, 4.993151, 4.992422, 4.991085, 
    4.989092, 4.986431, 4.982956, 4.978846, 4.973688, 4.967337, 4.959653, 
    4.950525, 4.939891, 4.927777, 4.914315, 4.899775, 4.884562, 4.869212, 
    4.85435, 4.840641, 4.828725, 4.819151, 4.812321, 4.808452, 4.807563, 
    4.809484,
  // momentumX(23,1, 0-49)
    4.896116, 4.90232, 4.908538, 4.914664, 4.920634, 4.92641, 4.931978, 
    4.937342, 4.942514, 4.947505, 4.952327, 4.956984, 4.961471, 4.965774, 
    4.969862, 4.97324, 4.977746, 4.980855, 4.983581, 4.985966, 4.987989, 
    4.990112, 4.991745, 4.993001, 4.993792, 4.994096, 4.993859, 4.993059, 
    4.991638, 4.989619, 4.986797, 4.983615, 4.979371, 4.973888, 4.966999, 
    4.958545, 4.948429, 4.936629, 4.923249, 4.908527, 4.892865, 4.876808, 
    4.861016, 4.846209, 4.8331, 4.822316, 4.814339, 4.809461, 4.807758, 
    4.809104,
  // momentumX(23,2, 0-49)
    4.896848, 4.903163, 4.909467, 4.915654, 4.921661, 4.927448, 4.933006, 
    4.938334, 4.943444, 4.948349, 4.953061, 4.957585, 4.961919, 4.966052, 
    4.96996, 4.972911, 4.977615, 4.980476, 4.982946, 4.985118, 4.986993, 
    4.989272, 4.991097, 4.992633, 4.993772, 4.994483, 4.9947, 4.994403, 
    4.993524, 4.99211, 4.989905, 4.987619, 4.98428, 4.979692, 4.973659, 
    4.965992, 4.956553, 4.945277, 4.932223, 4.917595, 4.901763, 4.885261, 
    4.868759, 4.853016, 4.838797, 4.826807, 4.81761, 4.81158, 4.808866, 
    4.809398,
  // momentumX(23,3, 0-49)
    4.897707, 4.904102, 4.910461, 4.91668, 4.922695, 4.928468, 4.933987, 
    4.939251, 4.944274, 4.949068, 4.953646, 4.958017, 4.962181, 4.966132, 
    4.969855, 4.972373, 4.977182, 4.979805, 4.98203, 4.983992, 4.985715, 
    4.988125, 4.990106, 4.991872, 4.993307, 4.994374, 4.994997, 4.99516, 
    4.994784, 4.993926, 4.992285, 4.990835, 4.988363, 4.984661, 4.979513, 
    4.972706, 4.964067, 4.953493, 4.940991, 4.926718, 4.910996, 4.894328, 
    4.877372, 4.860893, 4.845701, 4.832562, 4.822122, 4.814842, 4.810956, 
    4.810467,
  // momentumX(23,4, 0-49)
    4.898767, 4.905207, 4.911588, 4.917809, 4.923801, 4.929531, 4.934984, 
    4.940162, 4.945074, 4.949735, 4.954161, 4.958361, 4.962342, 4.966105, 
    4.969644, 4.971735, 4.976532, 4.978934, 4.980926, 4.982686, 4.984258, 
    4.986763, 4.988861, 4.990802, 4.992469, 4.993831, 4.994809, 4.995383, 
    4.99547, 4.995112, 4.993973, 4.993282, 4.991616, 4.988761, 4.984494, 
    4.978585, 4.970834, 4.9611, 4.949344, 4.935659, 4.920317, 4.903763, 
    4.886617, 4.869635, 4.853644, 4.839461, 4.827805, 4.819223, 4.814049, 
    4.812364,
  // momentumX(23,5, 0-49)
    4.900073, 4.906525, 4.912896, 4.919085, 4.925028, 4.930689, 4.93605, 
    4.941118, 4.945899, 4.950413, 4.95467, 4.958691, 4.962481, 4.966052, 
    4.969409, 4.971094, 4.975749, 4.977942, 4.979719, 4.981287, 4.982709, 
    4.985273, 4.987438, 4.989486, 4.991323, 4.992917, 4.994195, 4.995135, 
    4.995642, 4.995732, 4.995035, 4.995014, 4.994076, 4.992012, 4.988597, 
    4.983593, 4.976781, 4.967987, 4.957124, 4.94423, 4.929503, 4.913324, 
    4.896254, 4.879013, 4.862425, 4.847337, 4.834532, 4.824646, 4.818106, 
    4.815096,
  // momentumX(23,6, 0-49)
    4.901654, 4.908082, 4.914409, 4.920537, 4.926403, 4.931969, 4.937221, 
    4.94216, 4.946796, 4.951147, 4.95523, 4.959061, 4.962658, 4.966038, 
    4.969217, 4.970532, 4.974907, 4.976904, 4.978485, 4.979873, 4.981148, 
    4.983724, 4.985905, 4.987993, 4.989932, 4.991693, 4.993219, 4.994479, 
    4.995372, 4.995861, 4.995553, 4.996108, 4.995815, 4.994474, 4.991864, 
    4.987747, 4.98189, 4.974093, 4.964232, 4.952282, 4.938368, 4.922791, 
    4.906042, 4.888782, 4.87181, 4.855984, 4.842136, 4.830983, 4.823049, 
    4.818624,
  // momentumX(23,7, 0-49)
    4.903516, 4.909886, 4.916139, 4.922179, 4.927942, 4.933392, 4.938515, 
    4.943311, 4.947791, 4.951973, 4.955874, 4.959517, 4.96292, 4.966109, 
    4.96911, 4.97011, 4.974067, 4.975875, 4.977278, 4.9785, 4.979634, 
    4.982173, 4.984315, 4.986372, 4.988348, 4.990219, 4.991941, 4.99348, 
    4.994731, 4.995581, 4.995622, 4.996662, 4.996929, 4.996234, 4.994371, 
    4.991102, 4.986189, 4.979417, 4.970619, 4.959719, 4.946767, 4.931982, 
    4.915766, 4.898709, 4.881564, 4.86518, 4.85042, 4.838073, 4.82876, 4.82288,
  // momentumX(23,8, 0-49)
    4.905653, 4.911932, 4.918082, 4.924006, 4.929646, 4.934963, 4.939943, 
    4.944586, 4.948904, 4.952912, 4.956631, 4.960085, 4.963297, 4.966295, 
    4.969112, 4.969871, 4.973276, 4.974898, 4.97614, 4.977212, 4.978214, 
    4.980665, 4.982713, 4.984673, 4.986623, 4.988544, 4.990419, 4.992204, 
    4.99379, 4.994974, 4.995334, 4.996774, 4.997522, 4.997402, 4.996218, 
    4.993746, 4.989747, 4.98399, 4.976279, 4.966488, 4.954601, 4.940746, 
    4.925236, 4.908576, 4.891455, 4.874695, 4.859173, 4.845736, 4.835096, 
    4.827761,
  // momentumX(23,9, 0-49)
    4.908045, 4.914205, 4.920225, 4.926012, 4.931508, 4.936678, 4.941504, 
    4.945988, 4.95014, 4.953975, 4.957514, 4.960781, 4.963801, 4.966605, 
    4.969224, 4.969835, 4.972563, 4.973999, 4.975098, 4.976038, 4.976922, 
    4.979229, 4.981129, 4.982932, 4.984797, 4.986721, 4.988709, 4.99071, 
    4.992615, 4.994116, 4.994787, 4.996551, 4.997704, 4.998085, 4.997517, 
    4.995781, 4.992645, 4.987872, 4.981241, 4.972581, 4.961812, 4.948979, 
    4.934303, 4.918199, 4.901276, 4.884313, 4.868188, 4.853786, 4.841904, 
    4.833155,
  // momentumX(23,10, 0-49)
    4.910669, 4.916684, 4.922551, 4.928182, 4.93352, 4.938529, 4.943195, 
    4.947515, 4.951498, 4.955161, 4.958521, 4.961602, 4.96443, 4.967033, 
    4.969435, 4.969999, 4.971944, 4.973189, 4.97416, 4.974993, 4.975775, 
    4.977887, 4.979592, 4.981181, 4.982915, 4.984797, 4.986864, 4.989058, 
    4.991269, 4.993081, 4.994066, 4.996086, 4.997576, 4.998394, 4.998374, 
    4.997312, 4.994981, 4.991141, 4.985553, 4.978009, 4.968371, 4.956611, 
    4.942855, 4.927424, 4.910847, 4.893844, 4.877275, 4.862051, 4.849038, 
    4.838949,
  // momentumX(23,11, 0-49)
    4.9135, 4.919349, 4.925044, 4.930502, 4.935669, 4.94051, 4.945008, 
    4.94916, 4.952974, 4.956462, 4.959645, 4.96254, 4.965172, 4.967559, 
    4.969719, 4.970341, 4.971409, 4.972464, 4.973328, 4.974075, 4.974782, 
    4.976649, 4.978117, 4.979452, 4.981015, 4.982821, 4.984939, 4.9873, 
    4.989808, 4.991928, 4.993247, 4.995461, 4.997231, 4.998425, 4.998889, 
    4.998437, 4.996847, 4.993878, 4.989277, 4.98281, 4.974285, 4.963607, 
    4.950817, 4.936144, 4.92003, 4.903127, 4.886267, 4.870369, 4.856357, 
    4.845033,
  // momentumX(23,12, 0-49)
    4.916521, 4.922186, 4.927694, 4.932967, 4.937951, 4.942612, 4.946934, 
    4.950913, 4.954554, 4.957866, 4.960867, 4.963572, 4.965996, 4.968154, 
    4.970044, 4.970819, 4.970935, 4.971805, 4.972583, 4.973278, 4.97394, 
    4.975521, 4.976722, 4.97777, 4.979136, 4.98084, 4.982984, 4.985491, 
    4.988282, 4.990713, 4.99239, 4.994746, 4.996741, 4.998255, 4.999147, 
    4.999241, 4.998323, 4.996156, 4.992476, 4.987025, 4.97957, 4.969954, 
    4.958146, 4.944283, 4.928721, 4.912042, 4.895033, 4.878615, 4.863748, 
    4.851315,
  // momentumX(23,13, 0-49)
    4.919718, 4.925189, 4.930497, 4.935571, 4.940359, 4.944829, 4.948966, 
    4.952762, 4.956221, 4.95935, 4.962162, 4.964666, 4.966873, 4.968783, 
    4.970378, 4.971375, 4.97047, 4.971176, 4.971901, 4.972583, 4.97324, 
    4.9745, 4.975414, 4.976161, 4.977314, 4.978903, 4.981051, 4.983681, 
    4.98674, 4.989478, 4.991546, 4.993996, 4.996167, 4.997951, 4.999214, 
    4.999793, 4.999481, 4.998042, 4.995209, 4.990702, 4.984257, 4.975666, 
    4.964827, 4.951798, 4.936854, 4.920501, 4.903476, 4.886686, 4.871117, 
    4.857717,
  // momentumX(23,14, 0-49)
    4.92309, 4.928356, 4.933453, 4.938313, 4.942891, 4.947155, 4.95109, 
    4.954689, 4.957953, 4.960886, 4.963496, 4.96579, 4.967766, 4.969412, 
    4.970696, 4.97194, 4.96995, 4.970529, 4.971247, 4.971963, 4.972665, 
    4.973577, 4.974202, 4.97465, 4.975592, 4.977057, 4.979191, 4.981923, 
    4.985222, 4.988264, 4.990751, 4.99325, 4.995551, 4.997555, 4.999138, 
    5.000143, 5.000372, 4.999589, 4.997525, 4.993887, 4.988383, 4.980763, 
    4.970865, 4.958676, 4.944394, 4.928452, 4.91153, 4.894514, 4.878398, 
    4.864184,
  // momentumX(23,15, 0-49)
    4.926639, 4.931692, 4.936564, 4.941194, 4.945542, 4.949579, 4.95329, 
    4.956672, 4.959722, 4.962442, 4.964838, 4.966904, 4.968638, 4.970015, 
    4.970989, 4.972441, 4.969296, 4.969801, 4.970569, 4.97138, 4.972188, 
    4.972746, 4.973093, 4.973263, 4.974007, 4.975351, 4.977458, 4.980263, 
    4.983772, 4.9871, 4.99003, 4.992534, 4.99492, 4.997099, 4.99895, 
    5.000324, 5.001028, 5.000831, 4.999461, 4.996616, 4.99198, 4.985271, 
    4.976275, 4.96492, 4.95133, 4.93587, 4.919161, 4.902054, 4.885547, 
    4.870674,
  // momentumX(23,16, 0-49)
    4.93037, 4.935199, 4.939828, 4.944206, 4.948298, 4.952079, 4.95554, 
    4.958678, 4.961491, 4.96398, 4.966144, 4.967977, 4.969463, 4.970573, 
    4.971258, 4.972813, 4.968417, 4.968924, 4.969812, 4.970793, 4.971777, 
    4.971989, 4.972089, 4.97202, 4.972597, 4.973833, 4.975907, 4.978754, 
    4.982432, 4.986019, 4.989403, 4.991866, 4.994292, 4.996596, 4.998665, 
    5.000351, 5.00147, 5.001792, 5.001044, 4.998916, 4.995078, 4.989218, 
    4.981081, 4.970545, 4.957668, 4.942747, 4.926349, 4.909281, 4.892532, 
    4.877156,
  // momentumX(23,17, 0-49)
    4.934283, 4.938868, 4.943231, 4.947325, 4.951125, 4.954617, 4.957797, 
    4.960662, 4.963215, 4.965456, 4.967381, 4.968978, 4.970225, 4.971089, 
    4.971526, 4.973015, 4.967241, 4.967832, 4.968923, 4.970154, 4.971397, 
    4.971285, 4.971189, 4.970938, 4.971395, 4.972552, 4.974586, 4.97745, 
    4.981249, 4.985054, 4.988883, 4.991256, 4.99367, 4.99605, 4.998283, 
    5.000228, 5.001703, 5.002481, 5.002286, 5.000806, 4.997698, 4.992626, 
    4.985308, 4.975571, 4.96342, 4.94909, 4.933088, 4.91618, 4.89933, 4.883603,
  // momentumX(23,18, 0-49)
    4.938361, 4.942673, 4.946726, 4.950492, 4.953959, 4.957124, 4.95999, 
    4.962561, 4.964844, 4.966834, 4.968524, 4.969899, 4.970932, 4.971589, 
    4.971833, 4.973045, 4.96572, 4.966478, 4.967849, 4.969416, 4.971005, 
    4.970614, 4.970387, 4.970029, 4.97043, 4.971549, 4.973553, 4.976407, 
    4.980273, 4.98424, 4.988482, 4.990712, 4.993061, 4.995459, 4.9978, 
    4.999946, 5.001716, 5.002888, 5.003185, 5.00229, 4.99985, 4.995514, 
    4.988973, 4.980016, 4.968597, 4.9549, 4.939373, 4.922735, 4.905919, 
    4.889985,
  // momentumX(23,19, 0-49)
    4.942561, 4.94654, 4.950226, 4.953609, 4.956694, 4.959494, 4.962023, 
    4.964293, 4.96631, 4.96807, 4.969558, 4.970748, 4.971611, 4.972114, 
    4.972234, 4.972956, 4.963853, 4.964847, 4.966568, 4.968548, 4.970571, 
    4.969965, 4.969689, 4.969313, 4.969736, 4.970868, 4.972862, 4.97569, 
    4.979569, 4.98363, 4.988221, 4.990247, 4.992464, 4.994816, 4.9972, 
    4.999482, 5.001488, 5.002994, 5.003723, 5.003355, 5.001528, 4.99788, 
    4.992079, 4.983882, 4.973204, 4.960176, 4.945191, 4.928922, 4.912266, 
    4.896266,
  // momentumX(23,20, 0-49)
    4.947812, 4.952392, 4.956592, 4.960402, 4.963821, 4.966853, 4.969504, 
    4.971782, 4.973697, 4.975266, 4.976511, 4.977463, 4.978164, 4.978666, 
    4.97904, 0, 4.962282, 4.963513, 4.965213, 4.966989, 4.9687, 4.967034, 
    4.965853, 4.964697, 4.964581, 4.965442, 4.967443, 4.970533, 4.974926, 
    4.979701, 4.98531, 4.987769, 4.990425, 4.993213, 4.996024, 4.998729, 
    5.001162, 5.003111, 5.004313, 5.004456, 5.003191, 5.000156, 4.995014, 
    4.987504, 4.977509, 4.965121, 4.950686, 4.934827, 4.918398, 4.902422,
  // momentumX(23,21, 0-49)
    4.952321, 4.956649, 4.960524, 4.963956, 4.966967, 4.969578, 4.971817, 
    4.973706, 4.975272, 4.97654, 4.977539, 4.978305, 4.978885, 4.979341, 
    4.979759, 0, 4.957336, 4.958926, 4.96105, 4.963284, 4.965437, 4.96349, 
    4.962173, 4.960936, 4.960859, 4.961868, 4.964108, 4.967514, 4.972302, 
    4.977538, 4.983817, 4.986392, 4.989252, 4.992331, 4.995506, 4.998638, 
    5.001549, 5.004018, 5.005775, 5.006501, 5.005841, 5.003427, 4.99891, 
    4.992016, 4.982603, 4.970729, 4.956704, 4.941106, 4.924758, 4.90866,
  // momentumX(23,22, 0-49)
    4.956862, 4.960968, 4.964542, 4.967612, 4.970216, 4.972399, 4.974205, 
    4.975675, 4.97685, 4.977767, 4.978467, 4.978996, 4.979407, 4.979776, 
    4.98021, 0, 4.953183, 4.955079, 4.957577, 4.960221, 4.962775, 4.960561, 
    4.959106, 4.957771, 4.957701, 4.958802, 4.961205, 4.96483, 4.969896, 
    4.975457, 4.982234, 4.984813, 4.987763, 4.991016, 4.994449, 4.997913, 
    5.001224, 5.004153, 5.00642, 5.0077, 5.007632, 5.005837, 5.001956, 
    4.995699, 4.986902, 4.975594, 4.962046, 4.946799, 4.930641, 4.914544,
  // momentumX(23,23, 0-49)
    4.961319, 4.96523, 4.968522, 4.971242, 4.973449, 4.975204, 4.976571, 
    4.977608, 4.978371, 4.97891, 4.979281, 4.979536, 4.979744, 4.979992, 
    4.980406, 0, 4.949828, 4.951932, 4.954688, 4.957613, 4.960438, 4.957965, 
    4.956351, 4.954892, 4.954782, 4.955913, 4.958411, 4.962177, 4.967437, 
    4.973226, 4.980362, 4.982919, 4.985924, 4.989314, 4.992963, 4.996723, 
    5.000404, 5.00377, 5.006535, 5.008361, 5.008878, 5.007699, 5.004451, 
    4.998827, 4.990645, 4.979904, 4.966846, 4.951975, 4.936047, 4.920007,
  // momentumX(23,24, 0-49)
    4.965569, 4.969304, 4.972334, 4.974724, 4.976551, 4.977893, 4.978831, 
    4.979438, 4.979786, 4.97994, 4.979965, 4.979927, 4.979905, 4.98, 4.98035, 
    0, 4.947584, 4.949786, 4.952665, 4.955732, 4.958699, 4.956051, 4.954333, 
    4.952793, 4.952653, 4.953795, 4.956342, 4.960189, 4.965566, 4.971498, 
    4.97887, 4.981437, 4.984508, 4.988023, 4.991858, 4.995862, 4.999844, 
    5.003561, 5.006723, 5.008988, 5.009978, 5.009296, 5.006564, 5.001464, 
    4.993795, 4.983542, 4.970922, 4.956411, 4.940742, 4.924834,
  // momentumX(23,25, 0-49)
    4.969476, 4.973059, 4.975853, 4.977944, 4.97942, 4.980377, 4.980908, 
    4.981107, 4.981056, 4.98083, 4.980508, 4.980166, 4.979897, 4.979808, 
    4.980052, 0, 4.946215, 4.948393, 4.951257, 4.954316, 4.95728, 4.954575, 
    4.95283, 4.951283, 4.951154, 4.952318, 4.9549, 4.958794, 4.96423, 
    4.970243, 4.97773, 4.980377, 4.983562, 4.987227, 4.991247, 4.995472, 
    4.999707, 5.003707, 5.007178, 5.009773, 5.011113, 5.010795, 5.008437, 
    5.003716, 4.996426, 4.986541, 4.974265, 4.960062, 4.944643, 4.928911,
  // momentumX(23,26, 0-49)
    4.972922, 4.976376, 4.97897, 4.980797, 4.981965, 4.982578, 4.982746, 
    4.982569, 4.982144, 4.981558, 4.980897, 4.980248, 4.979712, 4.979408, 
    4.979493, 0, 4.945743, 4.947777, 4.950482, 4.953379, 4.956195, 4.95355, 
    4.951866, 4.950394, 4.950324, 4.951531, 4.954144, 4.95806, 4.963513, 
    4.969546, 4.977036, 4.979848, 4.983212, 4.987065, 4.991282, 4.995709, 
    5.000151, 5.00436, 5.008039, 5.010841, 5.012385, 5.012269, 5.010112, 
    5.005596, 4.998515, 4.988846, 4.976793, 4.962817, 4.947624, 4.932106,
  // momentumX(23,27, 0-49)
    4.975794, 4.979151, 4.981586, 4.983203, 4.984118, 4.984444, 4.9843, 
    4.983793, 4.983029, 4.982104, 4.981112, 4.980152, 4.979331, 4.978775, 
    4.978641, 0, 4.946302, 4.948066, 4.950467, 4.953045, 4.955564, 4.953069, 
    4.9515, 4.950153, 4.950165, 4.951417, 4.954041, 4.957945, 4.963362, 
    4.969354, 4.976735, 4.979789, 4.983385, 4.987454, 4.991872, 4.996479, 
    5.001076, 5.005418, 5.009205, 5.012092, 5.013698, 5.013628, 5.011506, 
    5.007021, 4.999983, 4.990378, 4.978427, 4.964598, 4.9496, 4.934321,
  // momentumX(23,28, 0-49)
    4.978009, 4.981311, 4.983644, 4.985114, 4.985842, 4.985948, 4.985551, 
    4.984766, 4.983699, 4.982455, 4.981137, 4.979851, 4.978716, 4.977863, 
    4.977447, 0, 4.948286, 4.949656, 4.951609, 4.953715, 4.955791, 4.953478, 
    4.952028, 4.950802, 4.950869, 4.952122, 4.9547, 4.958529, 4.963839, 
    4.969721, 4.97689, 4.98023, 4.984081, 4.988367, 4.992958, 4.997692, 
    5.002371, 5.006748, 5.010526, 5.01336, 5.014878, 5.014691, 5.012437, 
    5.007819, 5.000664, 4.990985, 4.979025, 4.965273, 4.950454, 4.935455,
  // momentumX(23,29, 0-49)
    4.979519, 4.98282, 4.985117, 4.98652, 4.987142, 4.987102, 4.986516, 
    4.985497, 4.984156, 4.982601, 4.980945, 4.979306, 4.977814, 4.976609, 
    4.975844, 0, 4.951502, 4.952365, 4.95373, 4.955213, 4.956685, 4.954491, 
    4.953069, 4.951875, 4.951902, 4.953065, 4.955513, 4.959191, 4.964319, 
    4.970014, 4.976858, 4.980478, 4.984567, 4.989044, 4.993778, 4.998605, 
    5.003326, 5.007692, 5.011411, 5.01414, 5.015511, 5.015141, 5.012679, 
    5.007847, 5.000496, 4.990666, 4.978632, 4.964911, 4.95025, 4.93554,
  // momentumX(23,30, 0-49)
    4.979384, 4.981814, 4.983278, 4.983901, 4.98382, 4.983175, 4.9821, 
    4.980711, 4.979107, 4.977366, 4.975537, 4.973642, 4.971686, 4.969653, 
    4.967526, 4.968501, 4.95388, 4.953983, 4.955086, 4.956669, 4.958492, 
    4.957497, 4.95718, 4.956963, 4.957675, 4.959179, 4.961603, 4.964932, 
    4.969421, 4.974288, 4.980054, 4.983217, 4.986848, 4.990884, 4.995209, 
    4.999662, 5.004045, 5.008105, 5.011535, 5.013987, 5.015082, 5.014435, 
    5.011695, 5.006598, 4.999016, 4.98902, 4.976917, 4.96326, 4.948817, 
    4.934488,
  // momentumX(23,31, 0-49)
    4.979453, 4.981999, 4.983564, 4.984265, 4.984229, 4.983586, 4.982464, 
    4.980983, 4.979244, 4.977332, 4.97531, 4.973215, 4.971061, 4.968839, 
    4.966521, 4.968116, 4.955175, 4.954739, 4.955228, 4.956167, 4.957366, 
    4.956451, 4.956088, 4.955835, 4.956506, 4.958014, 4.960509, 4.963962, 
    4.96857, 4.97352, 4.979156, 4.9828, 4.986884, 4.991324, 4.995992, 
    5.000715, 5.005282, 5.009428, 5.012842, 5.01517, 5.016033, 5.015054, 
    5.011901, 5.006335, 4.99827, 4.987822, 4.975352, 4.961461, 4.94695, 
    4.932743,
  // momentumX(23,32, 0-49)
    4.978727, 4.981336, 4.98298, 4.983766, 4.983811, 4.983236, 4.982162, 
    4.980702, 4.978957, 4.977013, 4.974936, 4.972773, 4.970546, 4.968249, 
    4.965855, 4.967472, 4.956299, 4.9554, 4.955333, 4.955686, 4.956318, 
    4.955542, 4.955204, 4.95499, 4.955684, 4.95724, 4.959817, 4.963375, 
    4.968049, 4.97302, 4.978463, 4.982544, 4.987028, 4.991814, 4.996756, 
    5.001674, 5.006341, 5.010485, 5.013781, 5.015877, 5.016394, 5.014968, 
    5.011288, 5.00515, 4.996514, 4.985552, 4.97268, 4.958555, 4.944016, 
    4.929998,
  // momentumX(23,33, 0-49)
    4.977302, 4.979942, 4.981656, 4.982538, 4.982697, 4.982244, 4.981289, 
    4.979935, 4.97828, 4.976404, 4.974379, 4.972252, 4.970052, 4.967782, 
    4.965415, 4.966619, 4.957237, 4.955972, 4.955427, 4.955264, 4.955398, 
    4.954807, 4.954551, 4.954451, 4.955221, 4.956857, 4.959517, 4.963147, 
    4.967824, 4.972751, 4.977959, 4.982429, 4.987256, 4.992321, 4.997468, 
    5.002501, 5.007183, 5.011227, 5.014306, 5.01606, 5.016119, 5.014136, 
    5.009826, 5.003026, 4.99375, 4.982231, 4.968952, 4.954619, 4.940107, 
    4.926363,
  // momentumX(23,34, 0-49)
    4.975289, 4.977936, 4.979716, 4.98071, 4.981011, 4.98072, 4.979937, 
    4.978752, 4.977258, 4.975528, 4.97363, 4.971616, 4.969521, 4.967354, 
    4.965097, 4.965625, 4.958004, 4.956473, 4.955529, 4.954925, 4.954628, 
    4.954253, 4.954134, 4.954203, 4.955094, 4.956829, 4.959558, 4.963218, 
    4.967833, 4.972657, 4.977599, 4.982405, 4.987512, 4.992789, 4.998067, 
    5.003136, 5.007743, 5.011593, 5.01435, 5.015658, 5.015156, 5.012516, 
    5.007489, 4.99996, 4.990002, 4.977917, 4.964249, 4.94976, 4.935356, 
    4.921988,
  // momentumX(23,35, 0-49)
    4.972805, 4.975446, 4.977287, 4.978399, 4.978864, 4.978765, 4.978192, 
    4.977223, 4.97594, 4.97441, 4.972696, 4.970852, 4.968914, 4.966905, 
    4.964818, 4.964561, 4.958642, 4.956938, 4.955672, 4.954696, 4.954036, 
    4.953892, 4.953948, 4.954236, 4.955279, 4.957119, 4.959894, 4.963537, 
    4.96802, 4.972685, 4.977338, 4.982416, 4.987737, 4.993151, 4.998478, 
    5.003494, 5.007935, 5.011493, 5.013832, 5.014596, 5.013438, 5.010059, 
    5.004251, 4.995952, 4.985302, 4.972674, 4.958676, 4.944117, 4.929926, 
    4.917049,
  // momentumX(23,36, 0-49)
    4.969972, 4.972589, 4.974487, 4.975722, 4.97636, 4.976475, 4.976136, 
    4.975414, 4.974378, 4.973086, 4.971597, 4.969959, 4.968216, 4.966397, 
    4.964516, 4.963494, 4.959198, 4.957397, 4.955878, 4.954597, 4.953636, 
    4.953732, 4.95399, 4.954529, 4.955745, 4.957692, 4.960482, 4.964052, 
    4.968329, 4.972781, 4.977126, 4.9824, 4.987854, 4.993322, 4.99861, 
    5.00348, 5.007657, 5.010827, 5.01265, 5.01278, 5.01089, 5.006711, 
    5.000083, 4.991011, 4.979698, 4.966591, 4.952356, 4.937846, 4.924, 
    4.911744,
  // momentumX(23,37, 0-49)
    4.966919, 4.969494, 4.971436, 4.972788, 4.973604, 4.973938, 4.973849, 
    4.973393, 4.972626, 4.971597, 4.970358, 4.968953, 4.967428, 4.965818, 
    4.964155, 4.96248, 4.959714, 4.957877, 4.956165, 4.954644, 4.953441, 
    4.953775, 4.954249, 4.955064, 4.95646, 4.9585, 4.961268, 4.964707, 
    4.968708, 4.972888, 4.976903, 4.982288, 4.987783, 4.99321, 4.998359, 
    5.002985, 5.006799, 5.009483, 5.010701, 5.010118, 5.007432, 5.002418, 
    4.994967, 4.985151, 4.973249, 4.959768, 4.945435, 4.931123, 4.917774, 
    4.906282,
  // momentumX(23,38, 0-49)
    4.963768, 4.966279, 4.968248, 4.969707, 4.970693, 4.971244, 4.971407, 
    4.971223, 4.970736, 4.969985, 4.969013, 4.967857, 4.966562, 4.96517, 
    4.963725, 4.96156, 4.96023, 4.958398, 4.956545, 4.954842, 4.953458, 
    4.95402, 4.954714, 4.955815, 4.95739, 4.959505, 4.962207, 4.965453, 
    4.969102, 4.972951, 4.976608, 4.982003, 4.987434, 4.992712, 4.997617, 
    5.001892, 5.005239, 5.007343, 5.007872, 5.006511, 5.002993, 4.997136, 
    4.988894, 4.978408, 4.96603, 4.952328, 4.938067, 4.924137, 4.911459, 
    4.90088,
  // momentumX(23,39, 0-49)
    4.960637, 4.963058, 4.965035, 4.96658, 4.967719, 4.968476, 4.968884, 
    4.968968, 4.968763, 4.968296, 4.967598, 4.966702, 4.965645, 4.964471, 
    4.963233, 4.960762, 4.96077, 4.958971, 4.957023, 4.955193, 4.953681, 
    4.954453, 4.955369, 4.956755, 4.958495, 4.960657, 4.963246, 4.966229, 
    4.969455, 4.972909, 4.976169, 4.981458, 4.986709, 4.99172, 4.996265, 
    5.000077, 5.002857, 5.00429, 5.004058, 5.001873, 4.997508, 4.990834, 
    4.981874, 4.970839, 4.958142, 4.944409, 4.930429, 4.917086, 4.905265, 
    4.895751,
  // momentumX(23,40, 0-49)
    4.95763, 4.959937, 4.961891, 4.963499, 4.964767, 4.965711, 4.966346, 
    4.966689, 4.966758, 4.96657, 4.966147, 4.965512, 4.964697, 4.963742, 
    4.962697, 4.960098, 4.961344, 4.959596, 4.957597, 4.95569, 4.954103, 
    4.95507, 4.956193, 4.957851, 4.959733, 4.961905, 4.964325, 4.966981, 
    4.969707, 4.972701, 4.975508, 4.980567, 4.98551, 4.990129, 4.99419, 
    4.997423, 4.999531, 5.000209, 4.99916, 4.996129, 4.990932, 4.983507, 
    4.973942, 4.962516, 4.949704, 4.936168, 4.922704, 4.910172, 4.8994, 
    4.891098,
  // momentumX(23,41, 0-49)
    4.95484, 4.957002, 4.958905, 4.960543, 4.961915, 4.963018, 4.963856, 
    4.964436, 4.964763, 4.964844, 4.96469, 4.964315, 4.963742, 4.963002, 
    4.962139, 4.959574, 4.961953, 4.96027, 4.958256, 4.956322, 4.954705, 
    4.955848, 4.957162, 4.959065, 4.961057, 4.963192, 4.965388, 4.967646, 
    4.9698, 4.972257, 4.974547, 4.979238, 4.983736, 4.987826, 4.991275, 
    4.993814, 4.995153, 4.995003, 4.993098, 4.989223, 4.983247, 4.975173, 
    4.965159, 4.953546, 4.940858, 4.927775, 4.915082, 4.903592, 4.89406, 
    4.887104,
  // momentumX(23,42, 0-49)
    4.952335, 4.954322, 4.956143, 4.957779, 4.959219, 4.960448, 4.961461, 
    4.962251, 4.962814, 4.963148, 4.963252, 4.963131, 4.962798, 4.962269, 
    4.961581, 4.959179, 4.962581, 4.960975, 4.958985, 4.95707, 4.955463, 
    4.956761, 4.958241, 4.960354, 4.962413, 4.964461, 4.966369, 4.96816, 
    4.96967, 4.971512, 4.973205, 4.977383, 4.981291, 4.984713, 4.987421, 
    4.989151, 4.989631, 4.988597, 4.985819, 4.981133, 4.974466, 4.965889, 
    4.955624, 4.944065, 4.931768, 4.919414, 4.907753, 4.897533, 4.889417, 
    4.883925,
  // momentumX(23,43, 0-49)
    4.950162, 4.951948, 4.953654, 4.955253, 4.956722, 4.958042, 4.959195, 
    4.960165, 4.960937, 4.9615, 4.961845, 4.961969, 4.961868, 4.961549, 
    4.961031, 4.958889, 4.963201, 4.961686, 4.959754, 4.957897, 4.956337, 
    4.957767, 4.959386, 4.961664, 4.963741, 4.965644, 4.967198, 4.968454, 
    4.96925, 4.970394, 4.971401, 4.97492, 4.97809, 4.980704, 4.982542, 
    4.983356, 4.982902, 4.980946, 4.977309, 4.971876, 4.964646, 4.955748, 
    4.945463, 4.934228, 4.922611, 4.91127, 4.900899, 4.892162, 4.885618, 
    4.881681,
  // momentumX(23,44, 0-49)
    4.948341, 4.9499, 4.951458, 4.952984, 4.954449, 4.955821, 4.957075, 
    4.958187, 4.959137, 4.959904, 4.96047, 4.960821, 4.960945, 4.960835, 
    4.960487, 4.958665, 4.963771, 4.962362, 4.960526, 4.958759, 4.957273, 
    4.958815, 4.960539, 4.962932, 4.96497, 4.966668, 4.967808, 4.968459, 
    4.968475, 4.968838, 4.96906, 4.971774, 4.974064, 4.975734, 4.976582, 
    4.976389, 4.974941, 4.972054, 4.967598, 4.961523, 4.953889, 4.944887, 
    4.934844, 4.92422, 4.913573, 4.903521, 4.894681, 4.887616, 4.882772, 
    4.88045,
  // momentumX(23,45, 0-49)
    4.946861, 4.948171, 4.949554, 4.950976, 4.952395, 4.95378, 4.955097, 
    4.956316, 4.957407, 4.958346, 4.959108, 4.95967, 4.960007, 4.960099, 
    4.959925, 4.958453, 4.964239, 4.962955, 4.961242, 4.959595, 4.958201, 
    4.959833, 4.961634, 4.964084, 4.966026, 4.967455, 4.968119, 4.968105, 
    4.967281, 4.966781, 4.966122, 4.967893, 4.969166, 4.96977, 4.969526, 
    4.968252, 4.96578, 4.961977, 4.956776, 4.950191, 4.942346, 4.933481, 
    4.923957, 4.914234, 4.904842, 4.896333, 4.889235, 4.883993, 4.880938, 
    4.880261,
  // momentumX(23,46, 0-49)
    4.945683, 4.946728, 4.947913, 4.949197, 4.950539, 4.951898, 4.953238, 
    4.954524, 4.955721, 4.9568, 4.957727, 4.958476, 4.959012, 4.959301, 
    4.959304, 4.958188, 4.964537, 4.963399, 4.961836, 4.96033, 4.959041, 
    4.960747, 4.962584, 4.965035, 4.966822, 4.967922, 4.968055, 4.967322, 
    4.965609, 4.964171, 4.962538, 4.963241, 4.963384, 4.962819, 4.961406, 
    4.959006, 4.955505, 4.950835, 4.944994, 4.938061, 4.930218, 4.921744, 
    4.913013, 4.904469, 4.896591, 4.889844, 4.884655, 4.881347, 4.88013, 
    4.881088,
  // momentumX(23,47, 0-49)
    4.944736, 4.945503, 4.946472, 4.947594, 4.948827, 4.950127, 4.951453, 
    4.952766, 4.954033, 4.955215, 4.956281, 4.957191, 4.957909, 4.958385, 
    4.958569, 4.957788, 4.964588, 4.96362, 4.962227, 4.960876, 4.959701, 
    4.961462, 4.963302, 4.965695, 4.96727, 4.967989, 4.967543, 4.96605, 
    4.96341, 4.960971, 4.958283, 4.957822, 4.956746, 4.954939, 4.952308, 
    4.948769, 4.944271, 4.938815, 4.932464, 4.925364, 4.917743, 4.909908, 
    4.902228, 4.895111, 4.888963, 4.884154, 4.880991, 4.879674, 4.8803, 
    4.882845,
  // momentumX(23,48, 0-49)
    4.943918, 4.9444, 4.945139, 4.946082, 4.947184, 4.948393, 4.949674, 
    4.950984, 4.952284, 4.953536, 4.954707, 4.955752, 4.956629, 4.957283, 
    4.957647, 4.957171, 4.964309, 4.96353, 4.962326, 4.961139, 4.960081, 
    4.961879, 4.963689, 4.965969, 4.967283, 4.967573, 4.966515, 4.964235, 
    4.960649, 4.957168, 4.953364, 4.951672, 4.949322, 4.946239, 4.942382, 
    4.93773, 4.932302, 4.926166, 4.919459, 4.91238, 4.905197, 4.898226, 
    4.891818, 4.886326, 4.882068, 4.87931, 4.878233, 4.878918, 4.881347, 
    4.885399,
  // momentumX(23,49, 0-49)
    4.943139, 4.943075, 4.943346, 4.94389, 4.944658, 4.945593, 4.946653, 
    4.94779, 4.948959, 4.950121, 4.951228, 4.952226, 4.953055, 4.953636, 
    4.953867, 4.95286, 4.96727, 4.965607, 4.963223, 4.960995, 4.959105, 
    4.962934, 4.966742, 4.971398, 4.97398, 4.974425, 4.972114, 4.967323, 
    4.959898, 4.952757, 4.94517, 4.942115, 4.938286, 4.93369, 4.928385, 
    4.922455, 4.916029, 4.909282, 4.902445, 4.895787, 4.889615, 4.884236, 
    4.879951, 4.877014, 4.875607, 4.87583, 4.877696, 4.881118, 4.885932, 
    4.8919,
  // momentumX(24,0, 0-49)
    4.910848, 4.916671, 4.922301, 4.927701, 4.932858, 4.937772, 4.942453, 
    4.946915, 4.951171, 4.955228, 4.959091, 4.962752, 4.9662, 4.969418, 
    4.972382, 4.974842, 4.97764, 4.97967, 4.981387, 4.98284, 4.984052, 
    4.985279, 4.986291, 4.987188, 4.987974, 4.988667, 4.989259, 4.989744, 
    4.990077, 4.99023, 4.990046, 4.989658, 4.988633, 4.986763, 4.983824, 
    4.979576, 4.973786, 4.966261, 4.95687, 4.945582, 4.932493, 4.917852, 
    4.902067, 4.8857, 4.869432, 4.854009, 4.840175, 4.8286, 4.81981, 4.81415,
  // momentumX(24,1, 0-49)
    4.911695, 4.917596, 4.923278, 4.928706, 4.933865, 4.938758, 4.943394, 
    4.94779, 4.951956, 4.955903, 4.959635, 4.963151, 4.96644, 4.969491, 
    4.972285, 4.974345, 4.977362, 4.979176, 4.980673, 4.981947, 4.983039, 
    4.984436, 4.985643, 4.986808, 4.987906, 4.988943, 4.989892, 4.990752, 
    4.991471, 4.992055, 4.9923, 4.992604, 4.992283, 4.991125, 4.988891, 
    4.985327, 4.980186, 4.973246, 4.964348, 4.95343, 4.940554, 4.92594, 
    4.909973, 4.89321, 4.876342, 4.860144, 4.845407, 4.832861, 4.823102, 
    4.816533,
  // momentumX(24,2, 0-49)
    4.912669, 4.91862, 4.924327, 4.929756, 4.934893, 4.93974, 4.944309, 
    4.948617, 4.952674, 4.956494, 4.960084, 4.963445, 4.966572, 4.969456, 
    4.972089, 4.973764, 4.97696, 4.978581, 4.979879, 4.980993, 4.981977, 
    4.983537, 4.984918, 4.986313, 4.987674, 4.988997, 4.990244, 4.99141, 
    4.992443, 4.993364, 4.993931, 4.994814, 4.995092, 4.994552, 4.992957, 
    4.990049, 4.985571, 4.979286, 4.97101, 4.96065, 4.948229, 4.933926, 
    4.918087, 4.901238, 4.884052, 4.867312, 4.851837, 4.8384, 4.827665, 
    4.820106,
  // momentumX(24,3, 0-49)
    4.91381, 4.919782, 4.925487, 4.93089, 4.935981, 4.940762, 4.945244, 
    4.949446, 4.953381, 4.957063, 4.960503, 4.963704, 4.966669, 4.969393, 
    4.971877, 4.973185, 4.976495, 4.977949, 4.979077, 4.98005, 4.980939, 
    4.982646, 4.984173, 4.98575, 4.987319, 4.988866, 4.990348, 4.991757, 
    4.993032, 4.994204, 4.994997, 4.996337, 4.997099, 4.997078, 4.996046, 
    4.993749, 4.98993, 4.984341, 4.976785, 4.967137, 4.955381, 4.941644, 
    4.92622, 4.909581, 4.892362, 4.875326, 4.859296, 4.845084, 4.833405, 
    4.824807,
  // momentumX(24,4, 0-49)
    4.915136, 4.921102, 4.926778, 4.932133, 4.937155, 4.941853, 4.946233, 
    4.950315, 4.954117, 4.957655, 4.960942, 4.963984, 4.966791, 4.969364, 
    4.971712, 4.972683, 4.976027, 4.977337, 4.978322, 4.979175, 4.979979, 
    4.981809, 4.983449, 4.985155, 4.986871, 4.988581, 4.990238, 4.991829, 
    4.993289, 4.994633, 4.995562, 4.997245, 4.998381, 4.99878, 4.998229, 
    4.996487, 4.993301, 4.988431, 4.98166, 4.972841, 4.961918, 4.948961, 
    4.934201, 4.918041, 4.901056, 4.883966, 4.867583, 4.852731, 4.840173, 
    4.830526,
  // momentumX(24,5, 0-49)
    4.916652, 4.922581, 4.928205, 4.933492, 4.938432, 4.943027, 4.947294, 
    4.951252, 4.954916, 4.958307, 4.961441, 4.964331, 4.966985, 4.969419, 
    4.971646, 4.972317, 4.975591, 4.976784, 4.977652, 4.978406, 4.979137, 
    4.981061, 4.982773, 4.984549, 4.986351, 4.988163, 4.989937, 4.99166, 
    4.993255, 4.994709, 4.995702, 4.997621, 4.999029, 4.999756, 4.999607, 
    4.99836, 4.995777, 4.99162, 4.985671, 4.977759, 4.967791, 4.95578, 
    4.941885, 4.926431, 4.909919, 4.893005, 4.876468, 4.861129, 4.847784, 
    4.837109,
  // momentumX(24,6, 0-49)
    4.918346, 4.924214, 4.929765, 4.934965, 4.939806, 4.944293, 4.948441, 
    4.952268, 4.955794, 4.959041, 4.962029, 4.96477, 4.967284, 4.969589, 
    4.971706, 4.972129, 4.975222, 4.976313, 4.97709, 4.977765, 4.978433, 
    4.980412, 4.982152, 4.983939, 4.985767, 4.98762, 4.989464, 4.991274, 
    4.992972, 4.994491, 4.995498, 4.997561, 4.999152, 5.000124, 5.000306, 
    4.999494, 4.997471, 4.994012, 4.988893, 4.98193, 4.972991, 4.96204, 
    4.949162, 4.934595, 4.918754, 4.902222, 4.885718, 4.870051, 4.856028, 
    4.844377,
  // momentumX(24,7, 0-49)
    4.920202, 4.925986, 4.931444, 4.936544, 4.941278, 4.945648, 4.949674, 
    4.953372, 4.956764, 4.959872, 4.962719, 4.965323, 4.967707, 4.969892, 
    4.971903, 4.972137, 4.97493, 4.975934, 4.976643, 4.977257, 4.977875, 
    4.979867, 4.981587, 4.983323, 4.985119, 4.986961, 4.988832, 4.990698, 
    4.992476, 4.994034, 4.995025, 4.997155, 4.998858, 5.000006, 5.000455, 
    5.000026, 4.99852, 4.995724, 4.991423, 4.985418, 4.977546, 4.96772, 
    4.955954, 4.942404, 4.92739, 4.911408, 4.89511, 4.879266, 4.864686, 
    4.852138,
  // momentumX(24,8, 0-49)
    4.922203, 4.927882, 4.933229, 4.938216, 4.942835, 4.947088, 4.95099, 
    4.954564, 4.957827, 4.960806, 4.963521, 4.965996, 4.968257, 4.970326, 
    4.972233, 4.972349, 4.97472, 4.975642, 4.976302, 4.976875, 4.977454, 
    4.979413, 4.981066, 4.982692, 4.984403, 4.986189, 4.988052, 4.989952, 
    4.991802, 4.993388, 4.994358, 4.996493, 4.998249, 4.999518, 5.000184, 
    5.000089, 4.999055, 4.996887, 4.993373, 4.988306, 4.981501, 4.972822, 
    4.962221, 4.949767, 4.935689, 4.92039, 4.904442, 4.888564, 4.873551, 
    4.860202,
  // momentumX(24,9, 0-49)
    4.924329, 4.929885, 4.935111, 4.939977, 4.944474, 4.948607, 4.95239, 
    4.955841, 4.958982, 4.961837, 4.964429, 4.966784, 4.968927, 4.970881, 
    4.972672, 4.972748, 4.974584, 4.975426, 4.976051, 4.9766, 4.977153, 
    4.97903, 4.980568, 4.982034, 4.983612, 4.985303, 4.987132, 4.989051, 
    4.990974, 4.992595, 4.993559, 4.995654, 4.997419, 4.998772, 4.999612, 
    4.999809, 4.999207, 4.997621, 4.994853, 4.990687, 4.98492, 4.977376, 
    4.967946, 4.956625, 4.943548, 4.929025, 4.913544, 4.897759, 4.88244, 
    4.868397,
  // momentumX(24,10, 0-49)
    4.926576, 4.931991, 4.937082, 4.941818, 4.946189, 4.950202, 4.953865, 
    4.957198, 4.960221, 4.962958, 4.965433, 4.967671, 4.969696, 4.971531, 
    4.973192, 4.97331, 4.974496, 4.975257, 4.975863, 4.976406, 4.976948, 
    4.978693, 4.980071, 4.981329, 4.982737, 4.984304, 4.98608, 4.98801, 
    4.990017, 4.99169, 4.992681, 4.994704, 4.996451, 4.997856, 4.998842, 
    4.999298, 4.999086, 4.998041, 4.995966, 4.992651, 4.98787, 4.981419, 
    4.973136, 4.962947, 4.9509, 4.937212, 4.922284, 4.906702, 4.891196, 
    4.876576,
  // momentumX(24,11, 0-49)
    4.928943, 4.934204, 4.939147, 4.943745, 4.947984, 4.95187, 4.955413, 
    4.958628, 4.961534, 4.964156, 4.966515, 4.968637, 4.97054, 4.972244, 
    4.973755, 4.973986, 4.97442, 4.975101, 4.975702, 4.976256, 4.976806, 
    4.978368, 4.97955, 4.980563, 4.981774, 4.983195, 4.984904, 4.986845, 
    4.988947, 4.990697, 4.991765, 4.993696, 4.995408, 4.996849, 4.997957, 
    4.998643, 4.998786, 4.998235, 4.996804, 4.994276, 4.990419, 4.985002, 
    4.977817, 4.968729, 4.957708, 4.944883, 4.930571, 4.91528, 4.899696, 
    4.884621,
  // momentumX(24,12, 0-49)
    4.931442, 4.936534, 4.941318, 4.945765, 4.949864, 4.953617, 4.957031, 
    4.960122, 4.962908, 4.965411, 4.967651, 4.969649, 4.971423, 4.972981, 
    4.974318, 4.974725, 4.974307, 4.974916, 4.975528, 4.976114, 4.976694, 
    4.978027, 4.978982, 4.979725, 4.98072, 4.981984, 4.983621, 4.985569, 
    4.98778, 4.989639, 4.990843, 4.992671, 4.994336, 4.995801, 4.997019, 
    4.997913, 4.998381, 4.998281, 4.997436, 4.995634, 4.992631, 4.988174, 
    4.982021, 4.973984, 4.963962, 4.952005, 4.938346, 4.923423, 4.907864, 
    4.892451,
  // momentumX(24,13, 0-49)
    4.934093, 4.939003, 4.943612, 4.947893, 4.951836, 4.955441, 4.958715, 
    4.961672, 4.964326, 4.966701, 4.968812, 4.970676, 4.972308, 4.973703, 
    4.974848, 4.975464, 4.974095, 4.974648, 4.975296, 4.975943, 4.976576, 
    4.977641, 4.978346, 4.978808, 4.97958, 4.980684, 4.982246, 4.984205, 
    4.986533, 4.988531, 4.989935, 4.991654, 4.993267, 4.994752, 4.996068, 
    4.997155, 4.997918, 4.99823, 4.997921, 4.996779, 4.994556, 4.990984, 
    4.985788, 4.978738, 4.969673, 4.958571, 4.94559, 4.931089, 4.915645, 
    4.900013,
  // momentumX(24,14, 0-49)
    4.936921, 4.94163, 4.946046, 4.950143, 4.953909, 4.957345, 4.96046, 
    4.963262, 4.96577, 4.968, 4.969966, 4.971681, 4.973152, 4.974371, 
    4.975314, 4.976134, 4.973717, 4.97424, 4.974955, 4.975695, 4.976418, 
    4.977182, 4.977629, 4.977811, 4.978366, 4.979317, 4.980805, 4.982772, 
    4.985224, 4.987384, 4.989049, 4.990658, 4.992219, 4.993719, 4.995128, 
    4.996392, 4.997429, 4.998117, 4.998294, 4.997752, 4.996239, 4.993473, 
    4.989157, 4.983024, 4.974865, 4.964593, 4.952296, 4.938266, 4.923021, 
    4.907284,
  // momentumX(24,15, 0-49)
    4.939954, 4.944445, 4.948641, 4.952525, 4.956085, 4.959326, 4.962252, 
    4.964876, 4.967212, 4.969275, 4.971076, 4.972627, 4.973923, 4.974956, 
    4.975694, 4.976676, 4.973099, 4.973635, 4.974455, 4.975329, 4.976182, 
    4.976626, 4.976819, 4.976738, 4.977095, 4.977906, 4.979325, 4.981301, 
    4.983872, 4.986211, 4.988193, 4.98969, 4.991199, 4.992713, 4.994207, 
    4.995636, 4.996924, 4.997959, 4.998579, 4.99858, 4.99771, 4.995675, 
    4.992167, 4.986881, 4.979572, 4.970099, 4.958487, 4.944963, 4.929991, 
    4.914255,
  // momentumX(24,16, 0-49)
    4.943211, 4.947452, 4.951399, 4.955036, 4.958356, 4.961365, 4.964069, 
    4.966485, 4.968622, 4.970495, 4.972114, 4.973482, 4.974594, 4.975438, 
    4.975983, 4.977036, 4.972176, 4.972776, 4.97375, 4.974805, 4.975837, 
    4.975954, 4.975911, 4.9756, 4.975791, 4.976484, 4.977843, 4.979822, 
    4.982503, 4.985028, 4.98737, 4.988751, 4.990204, 4.991729, 4.993303, 
    4.994886, 4.996407, 4.997757, 4.998783, 4.999278, 4.99899, 4.997621, 
    4.994846, 4.990343, 4.983829, 4.97512, 4.964186, 4.9512, 4.936568, 
    4.920935,
  // momentumX(24,17, 0-49)
    4.946694, 4.950654, 4.95431, 4.957654, 4.960692, 4.963429, 4.965877, 
    4.968051, 4.969965, 4.971627, 4.973047, 4.974223, 4.975149, 4.97581, 
    4.976184, 4.977188, 4.970901, 4.971617, 4.972795, 4.974083, 4.975348, 
    4.975148, 4.974903, 4.974407, 4.974476, 4.975085, 4.976398, 4.978378, 
    4.981153, 4.983857, 4.986584, 4.987842, 4.989233, 4.990761, 4.992407, 
    4.994132, 4.995866, 4.997506, 4.998901, 4.999847, 5.000089, 4.999326, 
    4.997222, 4.993437, 4.987666, 4.979686, 4.969424, 4.956998, 4.942767, 
    4.927331,
  // momentumX(24,18, 0-49)
    4.950392, 4.954015, 4.957329, 4.960334, 4.963038, 4.965462, 4.96762, 
    4.969528, 4.9712, 4.972644, 4.973861, 4.974846, 4.975591, 4.976085, 
    4.976321, 4.97714, 4.969261, 4.970144, 4.971568, 4.973141, 4.974692, 
    4.974195, 4.973797, 4.973176, 4.973178, 4.973746, 4.975035, 4.977013, 
    4.97986, 4.982726, 4.985838, 4.986964, 4.988281, 4.9898, 4.991502, 
    4.99335, 4.99528, 4.997187, 4.998922, 5.000279, 5.001005, 5.000793, 
    4.999304, 4.996184, 4.991109, 4.983826, 4.974225, 4.962378, 4.948599, 
    4.933446,
  // momentumX(24,19, 0-49)
    4.954257, 4.957479, 4.960381, 4.962982, 4.965306, 4.967378, 4.969222, 
    4.970854, 4.972284, 4.973517, 4.974545, 4.975358, 4.975943, 4.976294, 
    4.976423, 4.976936, 4.967296, 4.968376, 4.970076, 4.971971, 4.973859, 
    4.973104, 4.972607, 4.971929, 4.971931, 4.972509, 4.973804, 4.975785, 
    4.978683, 4.981678, 4.985153, 4.986128, 4.987349, 4.988836, 4.990572, 
    4.992523, 4.994625, 4.996772, 4.998816, 5.000549, 5.001719, 5.002016, 
    5.001093, 4.99859, 4.994166, 4.98755, 4.978599, 4.967349, 4.954068, 
    4.939276,
  // momentumX(24,20, 0-49)
    4.959174, 4.962858, 4.966164, 4.969108, 4.971708, 4.973982, 4.975949, 
    4.977625, 4.979029, 4.980179, 4.981099, 4.981818, 4.982371, 4.982801, 
    4.983164, 0, 4.964798, 4.966055, 4.967796, 4.969609, 4.971327, 4.969703, 
    4.968443, 4.967083, 4.966592, 4.9669, 4.968161, 4.970348, 4.973696, 
    4.977341, 4.981765, 4.983172, 4.984841, 4.986776, 4.988951, 4.991327, 
    4.993841, 4.996396, 4.998845, 5.000997, 5.002602, 5.003364, 5.002938, 
    5.000969, 4.997112, 4.991087, 4.982724, 4.972033, 4.959246, 4.944842,
  // momentumX(24,21, 0-49)
    4.963408, 4.966722, 4.969628, 4.972158, 4.974346, 4.976221, 4.977811, 
    4.979146, 4.980244, 4.981132, 4.981833, 4.982378, 4.982804, 4.983163, 
    4.983527, 0, 4.959586, 4.9611, 4.963162, 4.96533, 4.967396, 4.965482, 
    4.964082, 4.96265, 4.96222, 4.962704, 4.964239, 4.966779, 4.970561, 
    4.974705, 4.979818, 4.98141, 4.983339, 4.985602, 4.98816, 4.990963, 
    4.993931, 4.996956, 4.999882, 5.002509, 5.004585, 5.00581, 5.005842, 
    5.004326, 5.000915, 4.995324, 4.987371, 4.97705, 4.964567, 4.950371,
  // momentumX(24,22, 0-49)
    4.967702, 4.970664, 4.973182, 4.975305, 4.977076, 4.978538, 4.979732, 
    4.980693, 4.981451, 4.982034, 4.982473, 4.982803, 4.983067, 4.983329, 
    4.983677, 0, 4.955086, 4.956829, 4.959173, 4.961654, 4.964025, 4.961829, 
    4.960271, 4.958739, 4.958321, 4.95891, 4.960636, 4.963431, 4.967537, 
    4.97206, 4.977712, 4.979404, 4.981507, 4.984018, 4.986888, 4.990057, 
    4.993435, 4.9969, 5.000288, 5.003388, 5.00594, 5.007639, 5.008145, 
    5.007098, 5.004148, 4.999008, 4.99149, 4.981569, 4.969436, 4.955513,
  // momentumX(24,23, 0-49)
    4.971951, 4.974577, 4.976721, 4.978443, 4.979802, 4.980852, 4.98164, 
    4.982214, 4.98261, 4.982863, 4.983012, 4.983098, 4.983173, 4.983312, 
    4.983619, 0, 4.951283, 4.953178, 4.955709, 4.958392, 4.960952, 4.958478, 
    4.956745, 4.95508, 4.954624, 4.955256, 4.957099, 4.960074, 4.964422, 
    4.969233, 4.975299, 4.977072, 4.979327, 4.982063, 4.985225, 4.988744, 
    4.992522, 4.996426, 5.000281, 5.003865, 5.006908, 5.009098, 5.010088, 
    5.009516, 5.007031, 5.002338, 4.995245, 4.985715, 4.973922, 4.960277,
  // momentumX(24,24, 0-49)
    4.976042, 4.978349, 4.980137, 4.981477, 4.982438, 4.983085, 4.983476, 
    4.983662, 4.983689, 4.983603, 4.983446, 4.983268, 4.98313, 4.983118, 
    4.983349, 0, 4.948518, 4.95047, 4.953073, 4.955839, 4.958478, 4.955807, 
    4.953943, 4.952183, 4.951692, 4.952342, 4.954256, 4.957346, 4.961858, 
    4.966876, 4.973243, 4.975129, 4.977551, 4.980509, 4.98394, 4.987772, 
    4.991901, 4.996183, 5.000436, 5.004429, 5.007885, 5.010486, 5.011881, 
    5.011705, 5.009609, 5.005295, 4.998567, 4.989384, 4.97791, 4.964542,
  // momentumX(24,25, 0-49)
    4.979859, 4.981875, 4.983335, 4.984321, 4.984909, 4.985174, 4.985183, 
    4.984993, 4.984659, 4.984231, 4.983762, 4.983307, 4.982939, 4.982748, 
    4.982862, 0, 4.94658, 4.948485, 4.951038, 4.953754, 4.956346, 4.953585, 
    4.951666, 4.949878, 4.949385, 4.95006, 4.952026, 4.955197, 4.959819, 
    4.964978, 4.971531, 4.973589, 4.976222, 4.979423, 4.983128, 4.987259, 
    4.991705, 4.996318, 5.000906, 5.005232, 5.009016, 5.011939, 5.013646, 
    5.013772, 5.011967, 5.007938, 5.00149, 4.992584, 4.981378, 4.968261,
  // momentumX(24,26, 0-49)
    4.983298, 4.98506, 4.986228, 4.986894, 4.987146, 4.987062, 4.986718, 
    4.986174, 4.985493, 4.984731, 4.983946, 4.983204, 4.982584, 4.982186, 
    4.982136, 0, 4.945513, 4.947264, 4.949642, 4.952173, 4.954591, 4.951852, 
    4.949958, 4.948216, 4.947764, 4.948481, 4.95049, 4.953713, 4.958396, 
    4.963634, 4.970265, 4.972566, 4.975461, 4.978936, 4.982924, 4.987339, 
    4.992069, 4.996956, 5.001805, 5.006377, 5.010392, 5.013525, 5.015426, 
    5.015734, 5.014105, 5.01025, 5.003979, 4.99526, 4.984254, 4.97135,
  // momentumX(24,27, 0-49)
    4.986259, 4.987812, 4.988739, 4.989136, 4.989098, 4.988709, 4.988045, 
    4.987175, 4.986165, 4.985077, 4.983976, 4.982936, 4.982043, 4.9814, 
    4.981136, 0, 4.94546, 4.946948, 4.949024, 4.951235, 4.95335, 4.950716, 
    4.948902, 4.947252, 4.946861, 4.947614, 4.949643, 4.952878, 4.957563, 
    4.962814, 4.969408, 4.972008, 4.975201, 4.978966, 4.983234, 4.987912, 
    4.99288, 4.997982, 5.003019, 5.007753, 5.011899, 5.015141, 5.017131, 
    5.017511, 5.015946, 5.012156, 5.005963, 4.997341, 4.986464, 4.973726,
  // momentumX(24,28, 0-49)
    4.988665, 4.990068, 4.990814, 4.991004, 4.990735, 4.990089, 4.989146, 
    4.98798, 4.986658, 4.985248, 4.983824, 4.982468, 4.981272, 4.980346, 
    4.979819, 0, 4.946815, 4.947936, 4.949587, 4.951346, 4.953032, 4.950542, 
    4.948813, 4.947252, 4.946893, 4.947637, 4.949623, 4.952797, 4.957403, 
    4.962586, 4.969032, 4.971952, 4.975448, 4.97949, 4.984002, 4.98889, 
    4.994031, 4.999268, 5.004402, 5.0092, 5.013378, 5.016623, 5.018593, 
    5.018941, 5.017337, 5.013512, 5.007304, 4.998701, 4.987891, 4.975283,
  // momentumX(24,29, 0-49)
    4.990462, 4.991789, 4.992432, 4.992489, 4.992052, 4.991203, 4.990024, 
    4.988585, 4.986959, 4.985222, 4.983455, 4.981752, 4.980217, 4.978965, 
    4.978124, 0, 4.949393, 4.950053, 4.951162, 4.952341, 4.953464, 4.951066, 
    4.949343, 4.947788, 4.947369, 4.948007, 4.949859, 4.952889, 4.957327, 
    4.96235, 4.968523, 4.971735, 4.9755, 4.97978, 4.984496, 4.989554, 
    4.994829, 5.000166, 5.005371, 5.010205, 5.014393, 5.01762, 5.019548, 
    5.019832, 5.018151, 5.014245, 5.007967, 4.999325, 4.988527, 4.976,
  // momentumX(24,30, 0-49)
    4.990738, 4.99121, 4.991029, 4.990311, 4.989165, 4.987687, 4.985961, 
    4.984056, 4.982023, 4.979897, 4.977703, 4.975448, 4.973134, 4.970758, 
    4.968334, 4.967433, 4.952801, 4.952506, 4.95306, 4.954014, 4.955168, 
    4.953628, 4.952737, 4.951961, 4.952108, 4.953052, 4.954916, 4.957685, 
    4.961609, 4.965942, 4.971194, 4.974047, 4.977447, 4.981374, 4.985769, 
    4.990544, 4.995582, 5.000725, 5.005774, 5.010484, 5.014568, 5.017704, 
    5.019542, 5.019734, 5.017958, 5.013961, 5.007609, 4.998928, 4.988154, 
    4.975735,
  // momentumX(24,31, 0-49)
    4.991224, 4.991782, 4.991659, 4.990963, 4.989799, 4.988257, 4.986423, 
    4.984369, 4.982151, 4.979816, 4.977396, 4.974913, 4.972373, 4.969775, 
    4.967119, 4.966956, 4.953699, 4.952859, 4.952815, 4.953157, 4.953729, 
    4.952262, 4.951339, 4.950546, 4.950665, 4.951616, 4.953545, 4.956422, 
    4.960444, 4.964846, 4.969977, 4.973281, 4.977116, 4.981448, 4.986209, 
    4.991305, 4.996608, 5.001957, 5.007145, 5.011923, 5.016, 5.01905, 
    5.020725, 5.020681, 5.018607, 5.014267, 5.007555, 4.998531, 4.987468, 
    4.97485,
  // momentumX(24,32, 0-49)
    4.990952, 4.991582, 4.991526, 4.990881, 4.989748, 4.988213, 4.986357, 
    4.984251, 4.981956, 4.979523, 4.976988, 4.974381, 4.971712, 4.968981, 
    4.966177, 4.966247, 4.954534, 4.953211, 4.952619, 4.952398, 4.952437, 
    4.951101, 4.950212, 4.94947, 4.949618, 4.950622, 4.952628, 4.955601, 
    4.959674, 4.964085, 4.969033, 4.97274, 4.976955, 4.98163, 4.986691, 
    4.992035, 4.99753, 5.003008, 5.008257, 5.013021, 5.017007, 5.019885, 
    5.02131, 5.020944, 5.018488, 5.013731, 5.006595, 4.997181, 4.985804, 
    4.972989,
  // momentumX(24,33, 0-49)
    4.989976, 4.990683, 4.990708, 4.990148, 4.98909, 4.987619, 4.985811, 
    4.983734, 4.981448, 4.979006, 4.976447, 4.973802, 4.971087, 4.968307, 
    4.965442, 4.965351, 4.955271, 4.953551, 4.952481, 4.951764, 4.95134, 
    4.950182, 4.949387, 4.948767, 4.949002, 4.950088, 4.952173, 4.955213, 
    4.959281, 4.96364, 4.968359, 4.972418, 4.976954, 4.981907, 4.987197, 
    4.992716, 4.998327, 5.003853, 5.00908, 5.013745, 5.017552, 5.020169, 
    5.021256, 5.020481, 5.017564, 5.012319, 5.004707, 4.994871, 4.983172, 
    4.970181,
  // momentumX(24,34, 0-49)
    4.988362, 4.989154, 4.989285, 4.98884, 4.9879, 4.986543, 4.984841, 
    4.982858, 4.980649, 4.978268, 4.975753, 4.973141, 4.970451, 4.967691, 
    4.964846, 4.964324, 4.955907, 4.953883, 4.95241, 4.951271, 4.950449, 
    4.949511, 4.948865, 4.948426, 4.948793, 4.949985, 4.952144, 4.955214, 
    4.959218, 4.96347, 4.967926, 4.972286, 4.977082, 4.982247, 4.987697, 
    4.993318, 4.998965, 5.004459, 5.009578, 5.014056, 5.017594, 5.019861, 
    5.020521, 5.019255, 5.015803, 5.010012, 5.001885, 4.991614, 4.979609, 
    4.96648,
  // momentumX(24,35, 0-49)
    4.986187, 4.987076, 4.987331, 4.987029, 4.986242, 4.985043, 4.983495, 
    4.981658, 4.979582, 4.977318, 4.974906, 4.972382, 4.969771, 4.967087, 
    4.964324, 4.963235, 4.956457, 4.954219, 4.952422, 4.950934, 4.949782, 
    4.94909, 4.948639, 4.948434, 4.94897, 4.950284, 4.952501, 4.955562, 
    4.959439, 4.963533, 4.967704, 4.972306, 4.977299, 4.98261, 4.988148, 
    4.993796, 4.9994, 5.004778, 5.009702, 5.013903, 5.017081, 5.018907, 
    5.019053, 5.017218, 5.013171, 5.006792, 4.998133, 4.987436, 4.975163, 
    4.961967,
  // momentumX(24,36, 0-49)
    4.983537, 4.98453, 4.984925, 4.98479, 4.984187, 4.983179, 4.981824, 
    4.980174, 4.978276, 4.976174, 4.973908, 4.971516, 4.969026, 4.966462, 
    4.963827, 4.962144, 4.956951, 4.95458, 4.952532, 4.950767, 4.949354, 
    4.948923, 4.9487, 4.948773, 4.949505, 4.950946, 4.953201, 4.956208, 
    4.959899, 4.963787, 4.967659, 4.972442, 4.977566, 4.982953, 4.988503, 
    4.994096, 4.999576, 5.004749, 5.009388, 5.013221, 5.015947, 5.017244, 
    5.016798, 5.014329, 5.009636, 5.002648, 4.993464, 4.982381, 4.969909, 
    4.956739,
  // momentumX(24,37, 0-49)
    4.980508, 4.981606, 4.982151, 4.982196, 4.981798, 4.981007, 4.979875, 
    4.978444, 4.976758, 4.974855, 4.972772, 4.970547, 4.968214, 4.965799, 
    4.963324, 4.9611, 4.957419, 4.954983, 4.952751, 4.950772, 4.949162, 
    4.949, 4.949028, 4.949411, 4.950358, 4.951927, 4.954195, 4.957103, 
    4.96055, 4.96419, 4.967753, 4.97265, 4.977834, 4.983218, 4.988704, 
    4.99416, 4.999428, 5.004307, 5.008569, 5.01194, 5.014123, 5.014809, 
    5.013699, 5.010541, 5.005176, 4.997579, 4.987903, 4.976503, 4.963933, 
    4.950914,
  // momentumX(24,38, 0-49)
    4.977201, 4.978397, 4.979091, 4.979325, 4.979144, 4.978589, 4.977698, 
    4.976512, 4.975065, 4.97339, 4.971519, 4.969489, 4.967337, 4.965096, 
    4.962796, 4.960145, 4.957889, 4.955441, 4.953079, 4.950952, 4.949204, 
    4.949308, 4.949604, 4.950312, 4.951482, 4.953172, 4.955426, 4.958192, 
    4.96134, 4.964695, 4.967939, 4.972879, 4.978047, 4.983353, 4.988689, 
    4.993921, 4.998884, 5.003378, 5.007168, 5.009984, 5.011538, 5.011535, 
    5.0097, 5.005819, 4.999774, 4.991597, 4.981497, 4.96988, 4.957343, 
    4.944621,
  // momentumX(24,39, 0-49)
    4.973715, 4.974999, 4.975837, 4.976258, 4.976297, 4.975984, 4.975348, 
    4.974423, 4.973234, 4.971807, 4.970172, 4.968362, 4.966412, 4.964359, 
    4.962245, 4.959305, 4.958379, 4.955961, 4.953523, 4.9513, 4.949468, 
    4.949832, 4.950396, 4.951439, 4.95283, 4.954629, 4.956837, 4.959415, 
    4.962219, 4.965253, 4.968168, 4.973073, 4.978147, 4.983289, 4.988388, 
    4.993306, 4.997871, 5.001883, 5.005105, 5.007277, 5.00812, 5.007362, 
    5.004759, 5.000136, 4.993432, 4.984732, 4.974305, 4.962605, 4.950256, 
    4.938003,
  // momentumX(24,40, 0-49)
    4.970154, 4.971507, 4.972474, 4.973073, 4.973326, 4.973255, 4.972881, 
    4.972223, 4.971304, 4.970143, 4.968762, 4.967189, 4.965458, 4.963606, 
    4.96168, 4.958601, 4.958908, 4.956546, 4.954076, 4.951808, 4.949941, 
    4.950551, 4.951377, 4.952746, 4.95435, 4.956237, 4.958365, 4.960715, 
    4.96313, 4.96581, 4.968381, 4.973172, 4.978065, 4.982956, 4.987728, 
    4.992238, 4.996309, 4.999742, 5.002305, 5.003745, 5.003803, 5.002235, 
    4.998837, 4.993484, 4.986167, 4.977036, 4.966411, 4.954787, 4.942811, 
    4.931215,
  // momentumX(24,41, 0-49)
    4.966611, 4.968009, 4.969085, 4.969845, 4.970301, 4.970465, 4.970348, 
    4.969962, 4.969318, 4.968431, 4.967318, 4.965998, 4.964501, 4.962861, 
    4.961126, 4.958048, 4.959484, 4.957199, 4.954734, 4.952466, 4.950603, 
    4.951441, 4.952514, 4.954194, 4.955987, 4.957934, 4.959948, 4.96203, 
    4.964015, 4.966311, 4.968513, 4.973105, 4.977732, 4.982281, 4.98663, 
    4.990634, 4.994115, 4.996872, 4.998685, 4.999315, 4.998528, 4.996117, 
    4.99192, 4.985871, 4.978022, 4.96858, 4.957916, 4.946559, 4.935153, 
    4.924411,
  // momentumX(24,42, 0-49)
    4.963175, 4.964589, 4.965748, 4.966649, 4.96729, 4.967675, 4.967805, 
    4.967684, 4.967317, 4.966709, 4.96587, 4.964814, 4.963562, 4.962146, 
    4.960603, 4.957645, 4.960103, 4.957912, 4.955489, 4.953257, 4.951434, 
    4.952474, 4.953773, 4.955733, 4.957686, 4.959659, 4.961521, 4.963294, 
    4.964817, 4.966691, 4.968498, 4.972802, 4.977069, 4.98118, 4.985012, 
    4.988411, 4.991204, 4.993195, 4.994174, 4.993927, 4.992252, 4.988981, 
    4.984013, 4.977334, 4.969066, 4.959468, 4.948955, 4.938068, 4.927447, 
    4.917754,
  // momentumX(24,43, 0-49)
    4.959915, 4.961318, 4.962533, 4.963548, 4.964352, 4.964938, 4.965301, 
    4.965435, 4.965337, 4.965007, 4.964446, 4.963661, 4.962666, 4.96148, 
    4.960136, 4.957391, 4.960761, 4.95868, 4.956325, 4.954162, 4.952404, 
    4.953622, 4.955115, 4.957315, 4.959389, 4.961347, 4.963018, 4.964441, 
    4.965469, 4.966885, 4.968258, 4.972181, 4.975993, 4.979571, 4.982786, 
    4.985485, 4.987495, 4.988636, 4.988711, 4.987537, 4.984951, 4.980837, 
    4.97515, 4.967946, 4.959401, 4.94983, 4.939674, 4.929479, 4.919853, 
    4.911402,
  // momentumX(24,44, 0-49)
    4.956895, 4.958255, 4.959497, 4.960596, 4.961537, 4.962301, 4.962876, 
    4.963249, 4.963411, 4.963352, 4.963067, 4.962556, 4.961821, 4.960875, 
    4.959737, 4.957268, 4.961443, 4.959482, 4.957224, 4.955157, 4.953481, 
    4.954848, 4.956501, 4.958893, 4.961037, 4.962934, 4.964368, 4.965406, 
    4.965909, 4.966825, 4.967713, 4.971162, 4.974424, 4.97737, 4.979871, 
    4.981776, 4.98292, 4.983132, 4.98225, 4.98012, 4.976628, 4.971716, 
    4.965401, 4.957804, 4.949159, 4.93982, 4.930246, 4.920966, 4.912542, 
    4.905505,
  // momentumX(24,45, 0-49)
    4.954153, 4.955442, 4.956679, 4.957835, 4.958883, 4.959798, 4.960562, 
    4.961154, 4.961558, 4.961758, 4.961742, 4.961503, 4.961034, 4.960333, 
    4.959406, 4.957256, 4.962121, 4.960298, 4.958159, 4.956203, 4.954621, 
    4.95611, 4.957882, 4.960408, 4.962569, 4.964353, 4.96551, 4.966124, 
    4.966069, 4.96644, 4.966787, 4.969665, 4.972278, 4.974496, 4.976191, 
    4.977215, 4.977416, 4.976646, 4.974771, 4.971683, 4.967322, 4.961689, 
    4.95487, 4.947047, 4.938503, 4.929619, 4.920855, 4.912706, 4.905671, 
    4.900196,
  // momentumX(24,46, 0-49)
    4.951709, 4.952902, 4.954107, 4.955286, 4.956411, 4.957448, 4.958375, 
    4.959161, 4.959786, 4.960229, 4.960472, 4.960496, 4.96029, 4.959839, 
    4.959132, 4.957314, 4.962758, 4.961088, 4.95909, 4.957263, 4.955777, 
    4.957358, 4.959206, 4.961804, 4.963924, 4.965539, 4.966373, 4.966525, 
    4.965885, 4.965662, 4.965401, 4.967614, 4.969483, 4.970881, 4.971683, 
    4.97175, 4.970951, 4.969162, 4.966289, 4.962273, 4.957111, 4.950871, 
    4.943702, 4.935844, 4.927619, 4.919419, 4.911686, 4.904869, 4.899387, 
    4.895587,
  // momentumX(24,47, 0-49)
    4.949562, 4.950633, 4.951778, 4.952954, 4.954126, 4.955256, 4.956315, 
    4.957269, 4.95809, 4.958755, 4.959237, 4.959513, 4.959562, 4.959362, 
    4.958882, 4.957393, 4.963307, 4.961806, 4.959966, 4.958274, 4.956888, 
    4.958531, 4.960414, 4.963019, 4.965039, 4.966431, 4.966897, 4.96655, 
    4.965296, 4.964425, 4.963489, 4.964943, 4.965979, 4.966473, 4.966308, 
    4.965361, 4.963523, 4.960705, 4.956856, 4.951973, 4.946115, 4.939414, 
    4.932077, 4.924395, 4.916712, 4.90942, 4.902925, 4.897609, 4.893805, 
    4.891757,
  // momentumX(24,48, 0-49)
    4.94768, 4.948614, 4.949677, 4.950824, 4.952013, 4.953206, 4.954365, 
    4.955455, 4.956445, 4.957305, 4.958005, 4.958517, 4.958811, 4.958855, 
    4.958607, 4.95743, 4.963704, 4.962394, 4.960724, 4.959174, 4.957884, 
    4.959568, 4.961443, 4.963991, 4.965849, 4.966964, 4.967022, 4.966144, 
    4.964246, 4.962679, 4.960994, 4.961605, 4.961727, 4.961245, 4.960056, 
    4.958057, 4.95517, 4.951344, 4.946577, 4.940922, 4.934504, 4.927511, 
    4.920208, 4.912917, 4.905994, 4.899813, 4.894729, 4.891049, 4.889009, 
    4.888746,
  // momentumX(24,49, 0-49)
    4.945692, 4.946275, 4.947063, 4.948007, 4.949056, 4.950163, 4.951286, 
    4.952384, 4.953416, 4.954346, 4.955135, 4.95574, 4.956119, 4.956212, 
    4.955952, 4.954215, 4.967573, 4.965439, 4.962609, 4.960008, 4.957872, 
    4.961558, 4.965416, 4.970356, 4.973582, 4.975026, 4.974078, 4.971011, 
    4.965668, 4.960866, 4.955824, 4.955507, 4.954542, 4.952848, 4.950368, 
    4.947054, 4.942887, 4.937885, 4.932127, 4.925748, 4.918957, 4.912019, 
    4.905252, 4.899001, 4.89361, 4.88939, 4.886611, 4.885452, 4.886003, 
    4.888259,
  // momentumX(25,0, 0-49)
    4.925933, 4.931124, 4.936015, 4.940607, 4.944907, 4.948923, 4.952667, 
    4.956147, 4.959369, 4.962331, 4.965029, 4.967461, 4.969619, 4.971503, 
    4.973116, 4.974247, 4.975694, 4.976534, 4.977195, 4.977763, 4.978303, 
    4.97908, 4.979904, 4.98088, 4.98202, 4.983343, 4.984835, 4.986478, 
    4.988221, 4.990023, 4.991735, 4.993485, 4.994883, 4.995748, 4.995881, 
    4.995065, 4.993076, 4.989686, 4.984684, 4.977894, 4.969201, 4.95857, 
    4.946083, 4.931956, 4.916556, 4.9004, 4.884132, 4.868479, 4.854189, 
    4.841959,
  // momentumX(25,1, 0-49)
    4.927026, 4.932236, 4.937124, 4.941692, 4.945944, 4.949895, 4.953556, 
    4.956938, 4.960046, 4.962883, 4.965448, 4.967741, 4.96976, 4.971508, 
    4.972995, 4.97379, 4.975451, 4.976137, 4.976635, 4.977072, 4.977521, 
    4.978458, 4.979441, 4.980615, 4.981967, 4.983503, 4.985191, 4.98702, 
    4.988934, 4.99092, 4.992792, 4.994941, 4.996752, 4.998055, 4.998661, 
    4.998352, 4.996904, 4.994087, 4.98968, 4.983487, 4.975367, 4.965255, 
    4.953193, 4.939358, 4.924083, 4.907857, 4.891315, 4.875189, 4.860251, 
    4.847242,
  // momentumX(25,2, 0-49)
    4.928236, 4.933441, 4.938304, 4.942826, 4.947015, 4.950887, 4.954455, 
    4.95773, 4.960721, 4.963433, 4.965869, 4.968032, 4.969925, 4.971556, 
    4.972939, 4.973425, 4.975278, 4.975841, 4.976205, 4.97653, 4.976901, 
    4.977989, 4.979106, 4.980435, 4.981947, 4.983635, 4.985459, 4.987404, 
    4.989417, 4.991495, 4.993425, 4.995854, 4.997965, 4.999597, 5.000571, 
    5.000686, 4.999723, 4.997451, 4.993648, 4.988107, 4.980661, 4.97122, 
    4.959781, 4.946479, 4.931597, 4.91558, 4.899025, 4.882655, 4.867242, 
    4.853558,
  // momentumX(25,3, 0-49)
    4.929566, 4.934745, 4.939562, 4.944022, 4.948135, 4.951917, 4.955383, 
    4.958548, 4.961421, 4.964013, 4.966328, 4.968372, 4.970154, 4.971688, 
    4.972991, 4.973203, 4.975204, 4.975671, 4.975931, 4.976166, 4.976469, 
    4.977692, 4.978915, 4.980353, 4.981971, 4.983752, 4.985653, 4.987656, 
    4.989704, 4.991798, 4.993697, 4.996298, 4.998598, 5.000453, 5.001705, 
    5.00216, 5.001616, 4.99985, 4.996643, 4.991779, 4.985082, 4.976425, 
    4.965772, 4.953203, 4.938946, 4.923386, 4.907069, 4.890676, 4.874971, 
    4.860731,
  // momentumX(25,4, 0-49)
    4.931008, 4.93614, 4.940896, 4.945281, 4.949308, 4.952993, 4.956354, 
    4.959407, 4.962167, 4.964643, 4.966847, 4.968788, 4.970478, 4.971931, 
    4.973177, 4.973155, 4.975237, 4.975637, 4.975821, 4.975992, 4.976242, 
    4.977576, 4.978874, 4.98037, 4.982038, 4.983856, 4.98578, 4.987794, 
    4.98983, 4.991879, 4.993676, 4.996348, 4.998741, 5.000727, 5.002164, 
    5.002882, 5.002693, 5.001389, 4.998754, 4.994576, 4.988664, 4.980871, 
    4.971121, 4.959445, 4.946002, 4.931112, 4.915251, 4.899047, 4.883229, 
    4.868569,
  // momentumX(25,5, 0-49)
    4.932553, 4.937619, 4.942299, 4.9466, 4.950532, 4.954118, 4.957373, 
    4.960318, 4.962967, 4.965339, 4.967442, 4.969292, 4.970905, 4.9723, 
    4.973505, 4.973295, 4.975376, 4.975733, 4.975873, 4.975999, 4.976211, 
    4.977631, 4.978968, 4.980473, 4.982137, 4.983939, 4.985843, 4.987827, 
    4.98982, 4.991777, 4.993423, 4.996082, 4.998482, 5.000516, 5.002064, 
    5.002976, 5.003079, 5.002186, 5.000093, 4.996589, 4.991478, 4.984593, 
    4.975825, 4.965151, 4.952667, 4.938615, 4.923396, 4.907567, 4.891808, 
    4.876867,
  // momentumX(25,6, 0-49)
    4.934185, 4.93917, 4.943763, 4.94797, 4.951805, 4.955288, 4.95844, 
    4.961281, 4.963829, 4.966102, 4.968116, 4.96989, 4.97144, 4.97279, 
    4.973968, 4.973625, 4.975606, 4.975941, 4.976063, 4.97617, 4.976358, 
    4.977833, 4.979174, 4.980636, 4.982246, 4.983988, 4.985836, 4.987762, 
    4.989691, 4.991532, 4.992995, 4.995569, 4.997908, 4.999924, 5.001517, 
    5.00256, 5.002903, 5.002374, 5.000784, 4.997931, 4.993614, 4.987652, 
    4.979905, 4.970301, 4.958872, 4.945784, 4.931354, 4.916058, 4.900511, 
    4.885429,
  // momentumX(25,7, 0-49)
    4.935893, 4.940784, 4.94528, 4.949388, 4.953124, 4.956505, 4.959556, 
    4.962297, 4.964751, 4.966934, 4.968871, 4.970577, 4.972075, 4.973391, 
    4.974547, 4.974128, 4.975905, 4.976233, 4.976362, 4.976471, 4.976653, 
    4.97815, 4.979456, 4.980828, 4.98234, 4.983981, 4.985743, 4.987593, 
    4.989452, 4.991168, 4.992439, 4.994873, 4.997096, 4.999042, 5.000629, 
    5.001756, 5.002291, 5.002082, 5.000955, 4.998718, 4.995172, 4.990123, 
    4.983405, 4.974901, 4.964583, 4.952542, 4.939005, 4.924366, 4.909166, 
    4.894073,
  // momentumX(25,8, 0-49)
    4.937671, 4.942457, 4.946848, 4.950853, 4.954486, 4.957766, 4.960718, 
    4.963364, 4.965728, 4.96783, 4.969694, 4.971343, 4.972795, 4.974077, 
    4.975214, 4.97478, 4.976242, 4.976571, 4.97673, 4.976866, 4.977058, 
    4.97854, 4.979775, 4.981012, 4.982388, 4.983896, 4.985551, 4.987316, 
    4.98911, 4.990705, 4.991796, 4.994046, 4.996115, 4.997952, 4.999499, 
    5.00067, 5.001359, 5.001431, 5.000728, 4.999069, 4.996257, 4.992092, 
    4.986383, 4.978979, 4.969792, 4.958836, 4.946263, 4.932373, 4.91763, 
    4.902642,
  // momentumX(25,9, 0-49)
    4.939522, 4.944192, 4.948471, 4.952366, 4.955894, 4.959072, 4.961926, 
    4.964479, 4.966755, 4.96878, 4.970574, 4.972166, 4.973575, 4.974823, 
    4.975928, 4.975544, 4.976576, 4.976916, 4.977123, 4.977306, 4.977529, 
    4.978956, 4.980087, 4.981149, 4.982355, 4.983707, 4.985243, 4.986919, 
    4.988662, 4.990154, 4.991093, 4.993133, 4.995021, 4.996726, 4.998206, 
    4.999397, 5.00021, 5.000529, 5.000213, 4.999092, 4.996973, 4.993648, 
    4.988911, 4.982576, 4.974506, 4.964649, 4.953072, 4.939991, 4.92579, 
    4.911009,
  // momentumX(25,10, 0-49)
    4.941456, 4.945998, 4.950157, 4.953936, 4.957352, 4.960425, 4.963178, 
    4.965636, 4.967824, 4.96977, 4.971497, 4.973028, 4.974387, 4.975594, 
    4.976652, 4.976379, 4.976869, 4.977222, 4.977496, 4.977747, 4.978018, 
    4.979352, 4.980344, 4.981201, 4.982213, 4.983394, 4.984804, 4.986394, 
    4.988105, 4.989521, 4.990354, 4.992166, 4.993861, 4.99542, 4.99682, 
    4.998015, 4.998931, 4.999473, 4.999509, 4.998883, 4.997409, 4.994874, 
    4.991057, 4.985744, 4.978755, 4.969977, 4.959402, 4.947165, 4.933567, 
    4.919079,
  // momentumX(25,11, 0-49)
    4.943488, 4.947892, 4.951918, 4.955572, 4.958869, 4.961828, 4.964473, 
    4.96683, 4.968925, 4.970785, 4.972435, 4.973901, 4.975202, 4.976351, 
    4.977344, 4.977236, 4.977071, 4.977445, 4.9778, 4.978139, 4.978481, 
    4.979679, 4.980506, 4.981133, 4.981936, 4.982936, 4.984219, 4.985733, 
    4.98743, 4.988805, 4.98959, 4.991169, 4.992666, 4.994079, 4.995396, 
    4.996587, 4.997594, 4.998336, 4.998695, 4.998528, 4.99765, 4.995848, 
    4.992891, 4.988542, 4.982579, 4.97484, 4.96525, 4.953867, 4.940912, 
    4.926785,
  // momentumX(25,12, 0-49)
    4.94564, 4.949892, 4.953773, 4.957288, 4.960452, 4.963284, 4.965809, 
    4.968053, 4.970044, 4.971808, 4.973372, 4.974759, 4.975985, 4.977059, 
    4.97797, 4.978063, 4.977129, 4.977533, 4.97799, 4.978438, 4.978873, 
    4.979895, 4.980533, 4.980914, 4.981503, 4.982321, 4.983479, 4.984927, 
    4.986634, 4.988007, 4.988809, 4.990157, 4.991462, 4.992733, 4.993971, 
    4.995159, 4.996251, 4.997179, 4.997838, 4.998092, 4.997764, 4.996637, 
    4.994474, 4.991019, 4.986021, 4.979267, 4.970627, 4.960088, 4.947798, 
    4.934089,
  // momentumX(25,13, 0-49)
    4.947933, 4.952016, 4.955732, 4.959089, 4.962103, 4.964792, 4.967181, 
    4.969296, 4.971166, 4.972819, 4.97428, 4.975571, 4.976707, 4.977689, 
    4.978497, 4.978809, 4.976994, 4.977444, 4.978021, 4.978601, 4.979153, 
    4.979963, 4.980396, 4.980526, 4.980901, 4.981544, 4.982584, 4.983975, 
    4.985711, 4.987123, 4.988012, 4.989138, 4.990263, 4.991405, 4.992577, 
    4.993766, 4.994943, 4.996046, 4.996986, 4.997628, 4.997803, 4.997297, 
    4.995863, 4.99323, 4.989122, 4.983292, 4.975555, 4.965837, 4.95422, 
    4.94097,
  // momentumX(25,14, 0-49)
    4.950387, 4.954278, 4.957808, 4.960986, 4.963825, 4.966348, 4.968579, 
    4.970545, 4.972275, 4.973796, 4.975134, 4.976312, 4.977338, 4.97821, 
    4.978907, 4.979425, 4.97661, 4.97713, 4.977851, 4.978589, 4.979284, 
    4.979852, 4.980071, 4.979954, 4.980126, 4.980606, 4.981539, 4.982883, 
    4.984664, 4.98615, 4.987199, 4.988118, 4.989079, 4.990109, 4.991226, 
    4.99243, 4.993695, 4.994971, 4.996171, 4.997174, 4.99781, 4.99787, 
    4.997099, 4.995217, 4.991927, 4.98695, 4.980062, 4.971135, 4.960188, 
    4.947428,
  // momentumX(25,15, 0-49)
    4.953012, 4.956685, 4.960002, 4.96297, 4.965608, 4.967937, 4.969985, 
    4.971778, 4.973346, 4.974717, 4.975914, 4.976958, 4.977856, 4.978607, 
    4.979187, 4.979874, 4.975935, 4.976555, 4.977448, 4.97837, 4.979236, 
    4.979536, 4.979541, 4.979192, 4.97918, 4.979517, 4.980358, 4.981665, 
    4.983503, 4.985093, 4.986369, 4.987097, 4.987914, 4.988852, 4.989933, 
    4.991162, 4.992521, 4.993965, 4.995416, 4.996754, 4.997815, 4.998388, 
    4.998218, 4.997016, 4.99447, 4.990279, 4.98418, 4.976004, 4.965717, 
    4.95347,
  // momentumX(25,16, 0-49)
    4.955808, 4.959229, 4.9623, 4.965026, 4.967431, 4.969538, 4.971376, 
    4.972972, 4.974357, 4.975558, 4.976596, 4.97749, 4.978249, 4.978869, 
    4.979337, 4.980128, 4.974936, 4.975688, 4.976779, 4.977916, 4.978982, 
    4.978996, 4.978796, 4.978239, 4.978075, 4.978295, 4.979061, 4.980342, 
    4.982244, 4.983959, 4.98552, 4.986079, 4.986772, 4.987638, 4.9887, 
    4.989968, 4.99143, 4.993042, 4.994732, 4.996383, 4.997833, 4.998872, 
    4.999245, 4.998656, 4.996783, 4.993306, 4.987936, 4.98047, 4.970826, 
    4.959108,
  // momentumX(25,17, 0-49)
    4.958763, 4.961892, 4.964672, 4.96712, 4.969258, 4.971113, 4.972718, 
    4.974096, 4.975282, 4.976298, 4.977165, 4.9779, 4.978511, 4.979, 
    4.979367, 4.980179, 4.9736, 4.974513, 4.975829, 4.977204, 4.978499, 
    4.97822, 4.977831, 4.977103, 4.976825, 4.976961, 4.977675, 4.978942, 
    4.980911, 4.982769, 4.984655, 4.985065, 4.985654, 4.986466, 4.987527, 
    4.988847, 4.990417, 4.992199, 4.994118, 4.99606, 4.997868, 4.99933, 
    5.000191, 5.000153, 4.998885, 4.996056, 4.991358, 4.984556, 4.975537, 
    4.964358,
  // momentumX(25,18, 0-49)
    4.961843, 4.964629, 4.967072, 4.969197, 4.971034, 4.972611, 4.973962, 
    4.975113, 4.976092, 4.976921, 4.977616, 4.97819, 4.978654, 4.979015, 
    4.979291, 4.980046, 4.971954, 4.973047, 4.974599, 4.976233, 4.977781, 
    4.977211, 4.976659, 4.975799, 4.975451, 4.975545, 4.976236, 4.977504, 
    4.979541, 4.981548, 4.983785, 4.984062, 4.984563, 4.985336, 4.986408, 
    4.98779, 4.989474, 4.991421, 4.993559, 4.995777, 4.997911, 4.999756, 
    5.001056, 5.001511, 5.000786, 4.998543, 4.99446, 4.988282, 4.979865, 
    4.969234,
  // momentumX(25,19, 0-49)
    4.965, 4.967378, 4.969427, 4.971184, 4.972685, 4.973964, 4.975053, 
    4.975977, 4.976758, 4.977411, 4.977946, 4.978371, 4.978695, 4.978937, 
    4.979131, 4.97977, 4.970062, 4.97134, 4.973125, 4.975019, 4.976834, 
    4.975983, 4.975299, 4.974353, 4.973983, 4.974082, 4.974786, 4.976074, 
    4.978185, 4.980337, 4.982932, 4.983087, 4.983509, 4.98425, 4.985336, 
    4.986781, 4.988577, 4.990685, 4.993031, 4.995503, 4.99794, 5.000132, 
    5.001826, 5.002723, 5.002485, 5.000772, 4.997253, 4.991659, 4.983825, 
    4.973745,
  // momentumX(25,20, 0-49)
    4.96907, 4.971853, 4.97428, 4.976379, 4.978179, 4.979703, 4.980981, 
    4.982036, 4.982894, 4.983582, 4.984131, 4.98457, 4.984934, 4.985262, 
    4.9856, 0, 4.967362, 4.968657, 4.970433, 4.97227, 4.973977, 4.972389, 
    4.971055, 4.969516, 4.968708, 4.968553, 4.969211, 4.970665, 4.973172, 
    4.975917, 4.979388, 4.979959, 4.980811, 4.981984, 4.98349, 4.985337, 
    4.98751, 4.989974, 4.992662, 4.995465, 4.99823, 5.000757, 5.002801, 
    5.00407, 5.004237, 5.002963, 4.999919, 4.994827, 4.987511, 4.977941,
  // momentumX(25,21, 0-49)
    4.972409, 4.974806, 4.976856, 4.978595, 4.980055, 4.981269, 4.982268, 
    4.983077, 4.983721, 4.984225, 4.984614, 4.984921, 4.985179, 4.985434, 
    4.985746, 0, 4.962254, 4.963721, 4.965726, 4.967824, 4.969792, 4.9679, 
    4.966414, 4.964807, 4.964072, 4.964111, 4.965068, 4.966903, 4.969873, 
    4.97314, 4.977301, 4.978094, 4.979231, 4.980741, 4.982622, 4.984862, 
    4.987442, 4.990312, 4.993392, 4.996568, 4.999682, 5.002536, 5.004883, 
    5.006442, 5.00689, 5.005895, 5.003135, 4.998338, 4.991322, 4.982051,
  // momentumX(25,22, 0-49)
    4.97575, 4.977777, 4.979461, 4.980845, 4.981971, 4.982874, 4.983584, 
    4.984133, 4.984543, 4.984839, 4.985049, 4.985203, 4.985339, 4.98551, 
    4.985789, 0, 4.957802, 4.959422, 4.961627, 4.96395, 4.966136, 4.963939, 
    4.962275, 4.960557, 4.959836, 4.959994, 4.961162, 4.963283, 4.966613, 
    4.970295, 4.975018, 4.975973, 4.977332, 4.97912, 4.981323, 4.983923, 
    4.986884, 4.990145, 4.993617, 4.997175, 5.000654, 5.003854, 5.006526, 
    5.008392, 5.009137, 5.008434, 5.005967, 5.001472, 4.994767, 4.985815,
  // momentumX(25,23, 0-49)
    4.97903, 4.9807, 4.98203, 4.983072, 4.98387, 4.984463, 4.984885, 
    4.985168, 4.985334, 4.985412, 4.985426, 4.985411, 4.985411, 4.985483, 
    4.985715, 0, 4.953951, 4.955665, 4.95799, 4.960441, 4.962743, 4.960247, 
    4.958386, 4.956528, 4.955769, 4.955982, 4.957291, 4.959627, 4.96324, 
    4.967253, 4.972426, 4.973531, 4.9751, 4.977151, 4.979666, 4.982618, 
    4.98596, 4.98962, 4.993496, 4.997456, 5.001327, 5.004899, 5.007923, 
    5.010116, 5.011169, 5.010761, 5.00858, 5.00437, 4.997954, 4.989296,
  // momentumX(25,24, 0-49)
    4.982182, 4.983513, 4.984507, 4.985221, 4.985703, 4.985996, 4.986135, 
    4.98615, 4.98607, 4.985919, 4.985728, 4.985533, 4.98538, 4.985335, 
    4.985494, 0, 4.951048, 4.95278, 4.955128, 4.957605, 4.959929, 4.957211, 
    4.9552, 4.953234, 4.952438, 4.952682, 4.954084, 4.956569, 4.960389, 
    4.964658, 4.970174, 4.971457, 4.973247, 4.975561, 4.978374, 4.98165, 
    4.985334, 4.989345, 4.993575, 4.997882, 5.002086, 5.005975, 5.009296, 
    5.011769, 5.013084, 5.012925, 5.010993, 5.007029, 5.000869, 4.992476,
  // momentumX(25,25, 0-49)
    4.985147, 4.986164, 4.986844, 4.98725, 4.987433, 4.987438, 4.9873, 
    4.987053, 4.986725, 4.986343, 4.985937, 4.985548, 4.985225, 4.98504, 
    4.985095, 0, 4.948891, 4.950555, 4.952825, 4.955217, 4.957455, 4.95462, 
    4.952531, 4.950522, 4.949719, 4.949996, 4.95147, 4.954067, 4.958037, 
    4.962492, 4.968243, 4.969755, 4.971803, 4.974401, 4.977515, 4.981103, 
    4.985105, 4.989431, 4.993968, 4.998568, 5.003051, 5.007197, 5.010757, 
    5.013449, 5.014969, 5.015006, 5.013266, 5.009499, 5.003544, 4.99537,
  // momentumX(25,26, 0-49)
    4.987865, 4.9886, 4.988998, 4.98912, 4.989028, 4.98876, 4.988358, 
    4.987854, 4.987276, 4.986655, 4.986023, 4.985425, 4.98491, 4.984558, 
    4.98447, 0, 4.947531, 4.949038, 4.951124, 4.95332, 4.955368, 4.952527, 
    4.950438, 4.948456, 4.947687, 4.948007, 4.94954, 4.952215, 4.956279, 
    4.960855, 4.966729, 4.968522, 4.970867, 4.97377, 4.97719, 4.98108, 
    4.985371, 4.989972, 4.994764, 4.999599, 5.004291, 5.008625, 5.01235, 
    5.015193, 5.01685, 5.017016, 5.015405, 5.011773, 5.005966, 4.997958,
  // momentumX(25,27, 0-49)
    4.990288, 4.990781, 4.990932, 4.990807, 4.990461, 4.989943, 4.989286, 
    4.988528, 4.987698, 4.986828, 4.985954, 4.985124, 4.984395, 4.983844, 
    4.983571, 0, 4.947104, 4.948366, 4.950164, 4.952053, 4.953806, 4.951047, 
    4.949018, 4.947112, 4.946393, 4.946748, 4.948308, 4.951011, 4.9551, 
    4.959718, 4.965595, 4.967705, 4.970366, 4.973579, 4.977294, 4.981462, 
    4.986007, 4.990837, 4.995832, 5.000842, 5.005686, 5.010149, 5.013985, 
    5.016919, 5.018657, 5.018899, 5.017364, 5.013811, 5.008099, 5.000204,
  // momentumX(25,28, 0-49)
    4.992364, 4.99267, 4.992622, 4.992288, 4.991722, 4.990971, 4.990073, 
    4.989061, 4.987968, 4.986831, 4.985691, 4.984602, 4.983626, 4.982843, 
    4.982348, 0, 4.947995, 4.94893, 4.950346, 4.951824, 4.953187, 4.950557, 
    4.948601, 4.946773, 4.946075, 4.946415, 4.947931, 4.950579, 4.954597, 
    4.959157, 4.964909, 4.967333, 4.970298, 4.97379, 4.977762, 4.982154, 
    4.986895, 4.991891, 4.997024, 5.002145, 5.00708, 5.011614, 5.015508, 
    5.018489, 5.020265, 5.020542, 5.019038, 5.015524, 5.009858, 5.002028,
  // momentumX(25,29, 0-49)
    4.99406, 4.994244, 4.994057, 4.993563, 4.992815, 4.991854, 4.990718, 
    4.989445, 4.98807, 4.986638, 4.985197, 4.983812, 4.982553, 4.981504, 
    4.980756, 0, 4.950003, 4.95055, 4.951498, 4.952468, 4.953333, 4.950801, 
    4.948859, 4.947036, 4.946271, 4.946498, 4.947872, 4.950364, 4.954204, 
    4.958596, 4.964083, 4.966768, 4.969983, 4.973703, 4.97788, 4.982456, 
    4.98736, 4.992499, 4.997761, 5.002997, 5.008034, 5.012661, 5.016634, 
    5.019682, 5.021515, 5.021831, 5.020354, 5.016856, 5.011202, 5.003389,
  // momentumX(25,30, 0-49)
    4.994519, 4.993861, 4.992861, 4.991597, 4.990131, 4.988516, 4.986785, 
    4.984964, 4.983063, 4.981089, 4.979038, 4.976903, 4.974685, 4.97239, 
    4.970056, 4.968032, 4.954024, 4.95362, 4.953893, 4.954456, 4.955149, 
    4.953227, 4.951905, 4.950692, 4.950378, 4.950848, 4.952226, 4.954489, 
    4.957869, 4.961644, 4.966294, 4.968657, 4.97154, 4.974941, 4.978828, 
    4.983158, 4.987868, 4.99287, 4.998047, 5.00325, 5.008296, 5.012966, 
    5.017006, 5.020132, 5.02204, 5.022424, 5.021001, 5.017544, 5.01192, 
    5.004138,
  // momentumX(25,31, 0-49)
    4.995345, 4.994719, 4.99372, 4.992418, 4.990875, 4.98914, 4.98725, 
    4.985236, 4.983119, 4.98091, 4.978617, 4.976248, 4.9738, 4.97128, 
    4.968707, 4.967444, 4.954495, 4.953582, 4.953315, 4.953332, 4.953514, 
    4.951689, 4.950369, 4.949167, 4.948839, 4.949316, 4.950732, 4.953062, 
    4.956487, 4.960275, 4.964766, 4.967505, 4.970757, 4.974515, 4.978742, 
    4.983388, 4.988389, 4.993653, 4.999059, 5.004455, 5.009655, 5.014433, 
    5.018531, 5.02166, 5.023511, 5.023779, 5.022181, 5.018497, 5.012614, 
    5.004563,
  // momentumX(25,32, 0-49)
    4.995613, 4.995025, 4.99404, 4.992726, 4.991141, 4.989335, 4.987347, 
    4.985208, 4.982944, 4.980573, 4.978112, 4.975571, 4.972955, 4.970267, 
    4.967512, 4.966613, 4.954969, 4.953597, 4.952828, 4.952345, 4.952063, 
    4.950393, 4.949138, 4.948009, 4.947721, 4.948237, 4.949703, 4.952083, 
    4.955504, 4.959243, 4.96351, 4.966569, 4.97013, 4.97418, 4.978678, 
    4.983575, 4.988803, 4.994267, 4.999846, 5.005381, 5.010685, 5.015527, 
    5.019639, 5.022727, 5.024477, 5.024584, 5.022766, 5.018817, 5.01264, 
    5.00429,
  // momentumX(25,33, 0-49)
    4.995334, 4.994799, 4.993851, 4.992554, 4.990967, 4.989133, 4.987097, 
    4.984889, 4.982537, 4.980067, 4.977499, 4.97485, 4.972124, 4.969328, 
    4.966456, 4.965581, 4.955402, 4.953644, 4.952435, 4.951514, 4.95083, 
    4.949367, 4.948236, 4.947248, 4.947051, 4.947638, 4.949155, 4.951556, 
    4.954919, 4.958547, 4.962534, 4.96586, 4.96967, 4.973946, 4.978648, 
    4.983727, 4.989114, 4.994714, 5.000402, 5.006021, 5.011372, 5.016219, 
    5.020291, 5.023284, 5.024884, 5.024779, 5.022697, 5.01844, 5.011938, 
    5.003271,
  // momentumX(25,34, 0-49)
    4.994516, 4.994058, 4.993176, 4.991931, 4.990377, 4.98856, 4.986521, 
    4.984294, 4.981909, 4.979394, 4.976773, 4.974064, 4.971285, 4.968438, 
    4.965515, 4.964412, 4.955777, 4.953714, 4.952136, 4.950844, 4.949824, 
    4.94861, 4.947661, 4.946874, 4.946813, 4.947495, 4.949058, 4.95145, 
    4.954698, 4.95816, 4.961833, 4.965373, 4.969373, 4.97381, 4.978651, 
    4.983845, 4.989325, 4.994994, 5.000727, 5.006361, 5.011694, 5.016483, 
    5.020451, 5.02329, 5.024677, 5.024305, 5.02191, 5.017309, 5.010454, 
    5.001464,
  // momentumX(25,35, 0-49)
    4.993182, 4.992826, 4.992038, 4.990879, 4.989397, 4.987638, 4.985642, 
    4.983441, 4.98107, 4.978556, 4.975928, 4.97321, 4.970424, 4.967576, 
    4.96466, 4.963175, 4.9561, 4.953816, 4.951942, 4.95035, 4.949063, 
    4.948124, 4.947401, 4.946869, 4.946983, 4.94778, 4.949381, 4.95173, 
    4.954807, 4.958058, 4.961395, 4.965098, 4.969231, 4.97377, 4.978685, 
    4.983928, 4.989433, 4.995101, 5.000806, 5.006383, 5.011625, 5.016284, 
    5.020075, 5.022686, 5.023796, 5.023099, 5.02034, 5.015363, 5.008144, 
    4.998838,
  // momentumX(25,36, 0-49)
    4.99136, 4.991127, 4.990465, 4.989424, 4.988052, 4.986389, 4.984475, 
    4.982344, 4.980028, 4.97756, 4.974968, 4.972284, 4.969531, 4.966724, 
    4.963866, 4.961936, 4.956396, 4.953965, 4.951863, 4.950037, 4.948545, 
    4.947903, 4.94744, 4.947205, 4.947526, 4.948452, 4.950078, 4.95235, 
    4.955209, 4.958213, 4.961207, 4.965024, 4.969234, 4.973816, 4.978744, 
    4.983969, 4.989426, 4.995021, 5.000623, 5.006064, 5.011133, 5.01558, 
    5.019113, 5.02142, 5.022179, 5.021094, 5.017928, 5.012548, 5.004965, 
    4.995371,
  // momentumX(25,37, 0-49)
    4.989093, 4.989005, 4.988489, 4.987594, 4.986362, 4.984831, 4.983038, 
    4.981017, 4.9788, 4.976418, 4.973905, 4.97129, 4.968606, 4.965876, 
    4.963112, 4.960749, 4.956685, 4.954175, 4.951907, 4.949906, 4.948266, 
    4.947929, 4.947752, 4.947848, 4.9484, 4.949461, 4.951101, 4.953265, 
    4.955864, 4.958595, 4.961247, 4.96513, 4.969367, 4.973936, 4.978812, 
    4.983953, 4.989293, 4.994737, 5.000153, 5.005373, 5.010181, 5.014324, 
    5.01751, 5.019426, 5.01976, 5.018228, 5.014614, 5.008818, 5.000887, 
    4.991054,
  // momentumX(25,38, 0-49)
    4.986433, 4.986499, 4.986148, 4.985423, 4.98436, 4.982993, 4.981357, 
    4.979482, 4.977402, 4.975144, 4.972745, 4.970237, 4.967655, 4.965031, 
    4.962386, 4.959657, 4.956991, 4.954454, 4.952072, 4.949954, 4.948216, 
    4.948183, 4.948303, 4.948752, 4.949552, 4.950753, 4.952391, 4.954421, 
    4.956728, 4.959168, 4.961491, 4.965396, 4.969607, 4.974107, 4.978873, 
    4.983865, 4.989013, 4.994225, 4.999371, 5.004277, 5.008728, 5.012469, 
    5.015213, 5.016651, 5.016483, 5.014445, 5.010352, 5.00414, 4.995898, 
    4.985897,
  // momentumX(25,39, 0-49)
    4.98344, 4.983667, 4.983495, 4.982955, 4.982084, 4.980909, 4.979459, 
    4.977764, 4.975853, 4.973757, 4.971507, 4.969138, 4.966689, 4.964193, 
    4.961687, 4.95869, 4.957332, 4.954806, 4.952355, 4.950166, 4.948378, 
    4.948637, 4.949059, 4.949871, 4.950925, 4.952264, 4.953889, 4.955763, 
    4.957753, 4.959896, 4.961904, 4.965787, 4.969928, 4.974308, 4.978906, 
    4.983677, 4.988561, 4.99346, 4.998243, 5.002738, 5.006731, 5.009968, 
    5.01217, 5.013039, 5.012294, 5.0097, 5.00511, 4.998499, 4.990002, 4.97993,
  // momentumX(25,40, 0-49)
    4.980185, 4.980569, 4.980579, 4.980239, 4.979576, 4.978613, 4.977376, 
    4.975892, 4.974182, 4.972278, 4.970209, 4.96801, 4.96572, 4.963377, 
    4.961021, 4.957868, 4.957716, 4.955232, 4.952751, 4.950531, 4.948729, 
    4.949263, 4.949982, 4.951154, 4.952459, 4.953933, 4.955529, 4.957229, 
    4.95889, 4.960732, 4.962445, 4.966266, 4.970292, 4.974501, 4.978872, 
    4.983361, 4.987904, 4.992404, 4.996732, 5.000714, 5.004144, 5.006771, 
    5.008329, 5.008542, 5.007154, 5.003967, 4.998874, 4.9919, 4.983227, 
    4.973203,
  // momentumX(25,41, 0-49)
    4.976741, 4.977275, 4.977466, 4.97733, 4.976886, 4.976152, 4.975149, 
    4.973896, 4.972416, 4.970734, 4.968876, 4.966875, 4.964769, 4.962596, 
    4.960401, 4.957204, 4.958153, 4.95573, 4.953249, 4.951032, 4.949247, 
    4.950036, 4.951032, 4.952551, 4.954097, 4.955692, 4.957246, 4.958759, 
    4.960083, 4.96163, 4.963066, 4.966787, 4.970655, 4.974645, 4.978733, 
    4.982875, 4.987002, 4.991017, 4.994792, 4.998161, 5.000918, 5.00283, 
    5.003649, 5.003125, 5.001037, 4.997231, 4.991654, 4.984376, 4.975628, 
    4.965791,
  // momentumX(25,42, 0-49)
    4.973186, 4.973859, 4.974224, 4.97429, 4.974071, 4.973577, 4.972821, 
    4.971821, 4.970592, 4.969154, 4.967532, 4.965755, 4.963854, 4.96187, 
    4.959843, 4.956702, 4.958642, 4.956295, 4.953839, 4.951653, 4.949909, 
    4.950922, 4.952172, 4.954015, 4.955778, 4.957478, 4.958976, 4.96029, 
    4.961278, 4.962534, 4.963706, 4.967291, 4.970962, 4.974685, 4.978436, 
    4.982165, 4.985803, 4.989247, 4.992375, 4.995026, 4.997008, 4.998106, 
    4.998096, 4.996766, 4.993938, 4.989511, 4.983484, 4.975986, 4.967286, 
    4.957791,
  // momentumX(25,43, 0-49)
    4.969604, 4.970394, 4.970921, 4.971184, 4.971187, 4.970936, 4.970438, 
    4.969702, 4.968741, 4.967569, 4.966205, 4.964672, 4.962998, 4.961216, 
    4.959366, 4.956364, 4.959184, 4.95692, 4.954512, 4.952376, 4.950689, 
    4.951897, 4.953369, 4.955495, 4.957449, 4.959227, 4.960651, 4.961758, 
    4.962413, 4.963387, 4.964305, 4.967716, 4.971148, 4.97456, 4.977921, 
    4.981175, 4.984247, 4.987039, 4.989427, 4.991263, 4.992372, 4.992564, 
    4.99165, 4.989461, 4.985876, 4.980847, 4.974436, 4.966821, 4.958312, 
    4.949332,
  // momentumX(25,44, 0-49)
    4.966064, 4.966953, 4.967626, 4.968073, 4.968293, 4.968284, 4.968047, 
    4.967584, 4.966902, 4.966008, 4.964917, 4.963645, 4.962215, 4.960651, 
    4.958984, 4.956183, 4.95977, 4.9576, 4.955254, 4.953185, 4.951562, 
    4.952929, 4.954587, 4.956951, 4.959055, 4.960881, 4.962212, 4.963103, 
    4.963431, 4.964125, 4.96479, 4.967986, 4.971137, 4.974195, 4.977112, 
    4.979828, 4.982265, 4.984324, 4.98589, 4.986822, 4.986973, 4.986184, 
    4.984309, 4.981235, 4.976897, 4.971315, 4.964608, 4.957005, 4.948846, 
    4.940559,
  // momentumX(25,45, 0-49)
    4.962638, 4.963603, 4.964401, 4.965019, 4.965446, 4.965672, 4.965693, 
    4.965505, 4.965105, 4.964497, 4.96369, 4.962691, 4.961516, 4.960183, 
    4.958711, 4.95615, 4.96039, 4.958319, 4.956052, 4.954056, 4.952502, 
    4.953992, 4.955791, 4.95834, 4.960548, 4.962384, 4.963598, 4.964264, 
    4.96427, 4.96468, 4.965085, 4.968025, 4.97085, 4.973502, 4.975922, 
    4.978043, 4.97978, 4.981034, 4.9817, 4.981656, 4.98078, 4.978958, 
    4.976094, 4.972135, 4.967084, 4.961026, 4.954139, 4.946698, 4.939058, 
    4.931637,
  // momentumX(25,46, 0-49)
    4.959384, 4.960401, 4.961304, 4.962074, 4.962692, 4.963142, 4.963412, 
    4.963494, 4.963376, 4.963057, 4.962538, 4.961819, 4.96091, 4.959814, 
    4.958544, 4.956244, 4.961024, 4.959065, 4.956888, 4.954971, 4.95348, 
    4.955057, 4.95695, 4.959622, 4.961882, 4.963686, 4.964756, 4.965185, 
    4.964869, 4.964985, 4.965108, 4.967745, 4.970198, 4.972394, 4.974265, 
    4.975734, 4.97671, 4.977099, 4.976804, 4.975729, 4.973786, 4.970906, 
    4.967056, 4.962245, 4.956552, 4.950125, 4.9432, 4.936079, 4.92913, 
    4.922746,
  // momentumX(25,47, 0-49)
    4.95635, 4.957393, 4.95838, 4.959281, 4.960072, 4.960729, 4.961237, 
    4.961576, 4.961733, 4.961699, 4.961466, 4.961028, 4.960386, 4.959536, 
    4.958477, 4.956443, 4.961648, 4.959813, 4.957735, 4.955901, 4.954465, 
    4.956092, 4.958033, 4.960762, 4.963014, 4.964739, 4.965635, 4.965809, 
    4.965172, 4.964973, 4.964783, 4.967062, 4.969089, 4.970776, 4.972046, 
    4.972809, 4.972975, 4.972452, 4.971157, 4.969021, 4.966, 4.962074, 
    4.957274, 4.951685, 4.945455, 4.938794, 4.931985, 4.925356, 4.919264, 
    4.914069,
  // momentumX(25,48, 0-49)
    4.953563, 4.954612, 4.955658, 4.956668, 4.957611, 4.958456, 4.959181, 
    4.959764, 4.960183, 4.96042, 4.960465, 4.960305, 4.959929, 4.959326, 
    4.958488, 4.956709, 4.96223, 4.960528, 4.958559, 4.956808, 4.955421, 
    4.957064, 4.959004, 4.961722, 4.963907, 4.965501, 4.966192, 4.966093, 
    4.965123, 4.964581, 4.964033, 4.965894, 4.967434, 4.968557, 4.969174, 
    4.969187, 4.968502, 4.967037, 4.964726, 4.961534, 4.957456, 4.952534, 
    4.946867, 4.940608, 4.933976, 4.927238, 4.920715, 4.914744, 4.909664, 
    4.90578,
  // momentumX(25,49, 0-49)
    4.95051, 4.9514, 4.952364, 4.953356, 4.954337, 4.95527, 4.956123, 
    4.956862, 4.957456, 4.957881, 4.95811, 4.958118, 4.957881, 4.957365, 
    4.956535, 4.954092, 4.966395, 4.963832, 4.960638, 4.957756, 4.955451, 
    4.959006, 4.962871, 4.96796, 4.971593, 4.973686, 4.973638, 4.971708, 
    4.96775, 4.964478, 4.961112, 4.962604, 4.963628, 4.964084, 4.963889, 
    4.962953, 4.961198, 4.958563, 4.95502, 4.950583, 4.945317, 4.939349, 
    4.932869, 4.926122, 4.919407, 4.91305, 4.907397, 4.902774, 4.899466, 
    4.897687,
  // momentumX(26,0, 0-49)
    4.94, 4.944391, 4.94844, 4.952157, 4.95555, 4.958627, 4.961393, 4.963849, 
    4.965998, 4.96784, 4.969378, 4.970623, 4.97159, 4.972304, 4.9728, 
    4.972906, 4.973375, 4.973431, 4.973461, 4.973564, 4.973804, 4.974427, 
    4.975248, 4.976345, 4.977716, 4.979355, 4.981232, 4.983315, 4.985551, 
    4.987894, 4.990223, 4.992686, 4.994967, 4.996955, 4.998531, 4.999562, 
    4.999901, 4.999391, 4.997859, 4.995126, 4.991014, 4.985359, 4.978026, 
    4.968945, 4.958121, 4.945682, 4.931883, 4.917126, 4.901945, 4.886976,
  // momentumX(26,1, 0-49)
    4.941255, 4.945621, 4.949628, 4.95329, 4.956614, 4.959611, 4.962287, 
    4.96465, 4.966698, 4.96844, 4.96988, 4.971029, 4.971907, 4.972544, 
    4.972975, 4.97282, 4.973508, 4.973464, 4.973378, 4.973377, 4.973534, 
    4.974285, 4.975206, 4.976415, 4.977892, 4.979619, 4.981553, 4.983666, 
    4.985904, 4.988244, 4.990533, 4.993175, 4.995648, 4.997859, 4.999695, 
    5.00104, 5.001753, 5.001679, 5.000646, 4.998471, 4.994966, 4.989946, 
    4.983253, 4.97478, 4.964502, 4.952498, 4.938988, 4.924335, 4.909052, 
    4.893767,
  // momentumX(26,2, 0-49)
    4.942569, 4.946893, 4.950846, 4.954443, 4.957692, 4.960606, 4.963196, 
    4.965467, 4.967426, 4.969079, 4.970437, 4.971511, 4.972326, 4.97291, 
    4.973302, 4.972916, 4.973806, 4.973686, 4.973504, 4.973412, 4.973489, 
    4.974351, 4.975346, 4.976624, 4.978158, 4.979918, 4.981861, 4.983953, 
    4.986146, 4.988422, 4.990607, 4.993344, 4.995931, 4.998283, 5.000306, 
    5.001887, 5.002901, 5.0032, 5.002613, 5.00096, 4.998045, 4.993671, 
    4.987662, 4.979883, 4.970272, 4.958864, 4.945834, 4.931497, 4.916326, 
    4.900925,
  // momentumX(26,3, 0-49)
    4.943935, 4.948204, 4.952092, 4.955615, 4.958785, 4.961618, 4.964122, 
    4.966311, 4.968189, 4.969768, 4.97106, 4.97208, 4.972853, 4.973409, 
    4.973786, 4.973205, 4.974256, 4.974084, 4.97383, 4.973662, 4.973668, 
    4.974619, 4.975657, 4.976962, 4.978502, 4.98025, 4.982156, 4.984193, 
    4.986302, 4.988472, 4.990499, 4.99326, 4.995889, 4.99831, 5.000443, 
    5.002193, 5.003439, 5.004045, 5.003849, 5.002671, 5.000317, 4.996583, 
    4.991277, 4.984245, 4.975389, 4.964705, 4.952313, 4.938476, 4.923614, 
    4.908288,
  // momentumX(26,4, 0-49)
    4.945349, 4.949549, 4.953363, 4.956806, 4.959896, 4.962646, 4.96507, 
    4.967181, 4.96899, 4.970509, 4.97175, 4.972735, 4.973485, 4.974032, 
    4.974418, 4.973681, 4.974834, 4.974633, 4.974329, 4.974107, 4.97405, 
    4.975069, 4.976121, 4.977407, 4.978909, 4.980601, 4.982437, 4.984389, 
    4.986394, 4.988424, 4.990258, 4.992982, 4.995586, 4.998013, 5.000195, 
    5.002046, 5.003461, 5.004312, 5.004447, 5.003695, 5.001862, 4.998744, 
    4.994145, 4.987888, 4.979846, 4.969979, 4.958351, 4.945166, 4.930783, 
    4.915707,
  // momentumX(26,5, 0-49)
    4.946802, 4.950924, 4.954657, 4.958016, 4.961022, 4.96369, 4.966037, 
    4.968078, 4.969824, 4.971294, 4.9725, 4.973464, 4.974208, 4.974766, 
    4.975174, 4.974328, 4.975505, 4.975296, 4.974972, 4.974713, 4.974607, 
    4.97567, 4.976707, 4.977932, 4.979356, 4.980954, 4.982691, 4.984538, 
    4.986431, 4.988306, 4.989924, 4.992555, 4.995082, 4.997459, 4.999632, 
    5.001528, 5.003053, 5.004092, 5.004505, 5.004128, 5.002773, 5.000243, 
    4.996334, 4.99086, 4.983668, 4.974679, 4.963905, 4.951492, 4.937729, 
    4.923054,
  // momentumX(26,6, 0-49)
    4.948296, 4.952331, 4.955975, 4.959248, 4.962167, 4.964754, 4.967025, 
    4.969, 4.97069, 4.972117, 4.973296, 4.974251, 4.975002, 4.975583, 
    4.976024, 4.975116, 4.97623, 4.976032, 4.975711, 4.975441, 4.975303, 
    4.976385, 4.977377, 4.978502, 4.979811, 4.981283, 4.982903, 4.984636, 
    4.986417, 4.988131, 4.989528, 4.992019, 4.994424, 4.996704, 4.998821, 
    5.000714, 5.002299, 5.003477, 5.004117, 5.004066, 5.00315, 5.001173, 
    4.997931, 4.99323, 4.986898, 4.978821, 4.968964, 4.957409, 4.944374, 
    4.930231,
  // momentumX(26,7, 0-49)
    4.949835, 4.953774, 4.957324, 4.960505, 4.963335, 4.965837, 4.968033, 
    4.96994, 4.971579, 4.972966, 4.974124, 4.975074, 4.97584, 4.976448, 
    4.976927, 4.976012, 4.976964, 4.976792, 4.976501, 4.976244, 4.976095, 
    4.977169, 4.97809, 4.97908, 4.980241, 4.981565, 4.983052, 4.984669, 
    4.986344, 4.987903, 4.98909, 4.991405, 4.993648, 4.995795, 4.997818, 
    4.999667, 5.001273, 5.002547, 5.003373, 5.003607, 5.003088, 5.001628, 
    4.999024, 4.995079, 4.989602, 4.982448, 4.97354, 4.962898, 4.950672, 
    4.93716,
  // momentumX(26,8, 0-49)
    4.951429, 4.955265, 4.958713, 4.961794, 4.96453, 4.966943, 4.969059, 
    4.970898, 4.97248, 4.97383, 4.974967, 4.975914, 4.976696, 4.977333, 
    4.977845, 4.976974, 4.97766, 4.977527, 4.977291, 4.977073, 4.976935, 
    4.977974, 4.978799, 4.979623, 4.980614, 4.98177, 4.983119, 4.98462, 
    4.986207, 4.987626, 4.988623, 4.99073, 4.992783, 4.994769, 4.996668, 
    4.998445, 5.000041, 5.001379, 5.002355, 5.002841, 5.002684, 5.001705, 
    4.99971, 4.99649, 4.991849, 4.985611, 4.97766, 4.967961, 4.956597, 
    4.943792,
  // momentumX(26,9, 0-49)
    4.953088, 4.956812, 4.96015, 4.963123, 4.965757, 4.968074, 4.970102, 
    4.971866, 4.973389, 4.974695, 4.975805, 4.976745, 4.977537, 4.978196, 
    4.978734, 4.97796, 4.97827, 4.978189, 4.978033, 4.97788, 4.97778, 
    4.978755, 4.97946, 4.980095, 4.980895, 4.981874, 4.98308, 4.984471, 
    4.985987, 4.987292, 4.988131, 4.990008, 4.991851, 4.993655, 4.995411, 
    4.997094, 4.998659, 5.000037, 5.00114, 5.001849, 5.002026, 5.001497, 
    5.000074, 4.99755, 4.993714, 4.988372, 4.981369, 4.972619, 4.962144, 
    4.950095,
  // momentumX(26,10, 0-49)
    4.954827, 4.958428, 4.961646, 4.964502, 4.967022, 4.969234, 4.971165, 
    4.972841, 4.974293, 4.975544, 4.97662, 4.977544, 4.978334, 4.979006, 
    4.979555, 4.97893, 4.97875, 4.978733, 4.978679, 4.978618, 4.978583, 
    4.979466, 4.980032, 4.980456, 4.981056, 4.981851, 4.982915, 4.984207, 
    4.985671, 4.986889, 4.987614, 4.989247, 4.990867, 4.992477, 4.99408, 
    4.995658, 4.997178, 4.998582, 4.999794, 5.000707, 5.001192, 5.001086, 
    5.000204, 4.998339, 4.995272, 4.990792, 4.98471, 4.976898, 4.967317, 
    4.956054,
  // momentumX(26,11, 0-49)
    4.956657, 4.960123, 4.963208, 4.965933, 4.968327, 4.970419, 4.972239, 
    4.973818, 4.975185, 4.976367, 4.977395, 4.978288, 4.979064, 4.97973, 
    4.980277, 4.979839, 4.979058, 4.979119, 4.979188, 4.979247, 4.979304, 
    4.980065, 4.980476, 4.980678, 4.981071, 4.981682, 4.982608, 4.983808, 
    4.985242, 4.986406, 4.987069, 4.98845, 4.989841, 4.991255, 4.992701, 
    4.994172, 4.995643, 4.997068, 4.998378, 4.99948, 5.000252, 5.000543, 
    5.00017, 4.998927, 4.996589, 4.992929, 4.987732, 4.98083, 4.972133, 
    4.961664,
  // momentumX(26,12, 0-49)
    4.958586, 4.961901, 4.964838, 4.967417, 4.96967, 4.971628, 4.973322, 
    4.974786, 4.976053, 4.977152, 4.978113, 4.978957, 4.9797, 4.980344, 
    4.98087, 4.980648, 4.979154, 4.979307, 4.979526, 4.97973, 4.979906, 
    4.980518, 4.980759, 4.980734, 4.980921, 4.981354, 4.982149, 4.983266, 
    4.984689, 4.985831, 4.986491, 4.987618, 4.988783, 4.990006, 4.9913, 
    4.992667, 4.994092, 4.995536, 4.996943, 4.998224, 4.99927, 4.999934, 
    5.000038, 4.999378, 4.997725, 4.994837, 4.990478, 4.984446, 4.976607, 
    4.966925,
  // momentumX(26,13, 0-49)
    4.960617, 4.963764, 4.966533, 4.968949, 4.971044, 4.97285, 4.974402, 
    4.975734, 4.976882, 4.97788, 4.978757, 4.979533, 4.980224, 4.980828, 
    4.981322, 4.981328, 4.979001, 4.979272, 4.979662, 4.980037, 4.98036, 
    4.980793, 4.980856, 4.980605, 4.980595, 4.980857, 4.981531, 4.982577, 
    4.984003, 4.985156, 4.985874, 4.986757, 4.987704, 4.988744, 4.989898, 
    4.991172, 4.992559, 4.994028, 4.99553, 4.996988, 4.998293, 4.999307, 
    4.999858, 4.999741, 4.998724, 4.996556, 4.992984, 4.987775, 4.980757, 
    4.971845,
  // momentumX(26,14, 0-49)
    4.962743, 4.965701, 4.968283, 4.970517, 4.972435, 4.974072, 4.975463, 
    4.976647, 4.977662, 4.978541, 4.979313, 4.980003, 4.980623, 4.981172, 
    4.981625, 4.981853, 4.978575, 4.978984, 4.97957, 4.980143, 4.980638, 
    4.980866, 4.980747, 4.980277, 4.980084, 4.980192, 4.980755, 4.98174, 
    4.983183, 4.984377, 4.985216, 4.985863, 4.986608, 4.987482, 4.988513, 
    4.989711, 4.991073, 4.992577, 4.994179, 4.995807, 4.99736, 4.998702, 
    4.999669, 5.000055, 4.999626, 4.998124, 4.995279, 4.99084, 4.984598, 
    4.976427,
  // momentumX(26,15, 0-49)
    4.96495, 4.967693, 4.970068, 4.972099, 4.973822, 4.975271, 4.976488, 
    4.977509, 4.978373, 4.979118, 4.979771, 4.980357, 4.980891, 4.98137, 
    4.981779, 4.982203, 4.977856, 4.978431, 4.979234, 4.980026, 4.980718, 
    4.98072, 4.98042, 4.979746, 4.97939, 4.979363, 4.979831, 4.980763, 
    4.982235, 4.983498, 4.984517, 4.984947, 4.985507, 4.986237, 4.987163, 
    4.988302, 4.989655, 4.991206, 4.992913, 4.99471, 4.996499, 4.998151, 
    4.999502, 5.000349, 5.000455, 4.999561, 4.997384, 4.993657, 4.98814, 
    4.980677,
  // momentumX(26,16, 0-49)
    4.967216, 4.969719, 4.971859, 4.973665, 4.975173, 4.97642, 4.977448, 
    4.978295, 4.979, 4.979597, 4.98012, 4.98059, 4.981026, 4.981429, 4.98179, 
    4.98237, 4.976842, 4.977604, 4.978645, 4.979676, 4.980588, 4.980343, 
    4.979868, 4.979012, 4.978518, 4.978383, 4.978773, 4.979663, 4.981173, 
    4.982527, 4.983779, 4.984013, 4.984412, 4.98502, 4.985863, 4.986963, 
    4.988326, 4.989933, 4.991749, 4.993711, 4.995725, 4.997665, 4.999369, 
    5.000635, 5.001229, 5.000884, 4.999315, 4.996238, 4.991397, 4.984601,
  // momentumX(26,17, 0-49)
    4.969512, 4.97174, 4.973618, 4.975176, 4.976452, 4.977484, 4.978314, 
    4.97898, 4.979518, 4.979966, 4.980352, 4.980701, 4.981031, 4.981352, 
    4.981671, 4.982362, 4.975548, 4.976512, 4.977801, 4.979086, 4.980233, 
    4.979731, 4.979088, 4.978076, 4.977477, 4.977263, 4.977597, 4.978462, 
    4.980017, 4.981482, 4.98301, 4.983071, 4.983333, 4.983841, 4.984626, 
    4.985706, 4.987091, 4.988766, 4.990695, 4.99282, 4.995048, 4.997253, 
    4.999278, 5.000922, 5.001952, 5.002101, 5.001079, 4.998593, 4.994374, 
    4.988206,
  // momentumX(26,18, 0-49)
    4.971802, 4.973717, 4.975297, 4.976582, 4.977609, 4.978417, 4.979047, 
    4.979535, 4.979914, 4.980217, 4.98047, 4.980698, 4.980921, 4.981159, 
    4.981435, 4.982197, 4.974019, 4.975191, 4.976727, 4.978267, 4.979657, 
    4.978886, 4.978089, 4.97695, 4.976281, 4.976023, 4.97633, 4.977189, 
    4.978799, 4.980386, 4.982221, 4.982135, 4.982282, 4.982712, 4.983455, 
    4.984532, 4.985951, 4.9877, 4.989746, 4.992026, 4.994454, 4.996904, 
    4.999218, 5.001203, 5.002622, 5.003211, 5.00268, 5.00073, 4.99708, 
    4.991498,
  // momentumX(26,19, 0-49)
    4.974044, 4.975593, 4.976839, 4.977823, 4.978588, 4.979169, 4.979604, 
    4.979926, 4.980161, 4.980335, 4.98047, 4.980588, 4.98071, 4.980864, 
    4.981096, 4.981905, 4.972337, 4.973706, 4.975469, 4.977249, 4.978876, 
    4.977831, 4.976893, 4.975658, 4.974956, 4.974691, 4.975004, 4.975879, 
    4.977556, 4.979274, 4.981433, 4.981222, 4.981273, 4.981641, 4.982354, 
    4.983438, 4.984897, 4.986722, 4.98888, 4.991309, 4.993922, 4.996593, 
    4.999171, 5.001457, 5.003224, 5.004207, 5.004115, 5.00265, 4.999523, 
    4.994492,
  // momentumX(26,20, 0-49)
    4.977043, 4.979004, 4.980653, 4.982024, 4.983145, 4.984046, 4.984755, 
    4.985302, 4.985719, 4.986032, 4.986275, 4.986479, 4.986677, 4.986904, 
    4.987205, 0, 4.969875, 4.971127, 4.972816, 4.974531, 4.976083, 4.974407, 
    4.972915, 4.971169, 4.97008, 4.969584, 4.969836, 4.970838, 4.972848, 
    4.975082, 4.978014, 4.978158, 4.978577, 4.979314, 4.980385, 4.981804, 
    4.983576, 4.985689, 4.988112, 4.990792, 4.993645, 4.996556, 4.999379, 
    5.001928, 5.003983, 5.005283, 5.005549, 5.004485, 5.001798, 4.997241,
  // momentumX(26,21, 0-49)
    4.97925, 4.980883, 4.98223, 4.983332, 4.984216, 4.984912, 4.985448, 
    4.985849, 4.986141, 4.98635, 4.9865, 4.986621, 4.986745, 4.986916, 
    4.987184, 0, 4.965111, 4.966493, 4.968369, 4.970301, 4.97207, 4.970103, 
    4.968467, 4.966664, 4.965661, 4.965364, 4.965918, 4.967295, 4.969753, 
    4.972483, 4.976055, 4.976404, 4.977072, 4.978096, 4.979475, 4.981217, 
    4.983313, 4.985742, 4.988464, 4.991421, 4.994527, 4.997666, 5.000692, 
    5.003428, 5.005657, 5.007132, 5.007581, 5.006714, 5.004252, 4.999951,
  // momentumX(26,22, 0-49)
    4.981404, 4.982722, 4.983783, 4.984627, 4.985284, 4.985783, 4.986148, 
    4.986403, 4.986568, 4.986663, 4.986715, 4.986749, 4.986797, 4.986908, 
    4.98714, 0, 4.96099, 4.962482, 4.964514, 4.966624, 4.968567, 4.966304, 
    4.964496, 4.962591, 4.961608, 4.961434, 4.962199, 4.963859, 4.966667, 
    4.969792, 4.973887, 4.974385, 4.975251, 4.976512, 4.978163, 4.980196, 
    4.982597, 4.985335, 4.988364, 4.991613, 4.994995, 4.998389, 5.00165, 
    5.004604, 5.007035, 5.008707, 5.009351, 5.008693, 5.006459, 5.002415,
  // momentumX(26,23, 0-49)
    4.983479, 4.984495, 4.985284, 4.985883, 4.986323, 4.986632, 4.986832, 
    4.98694, 4.986977, 4.986959, 4.986909, 4.98685, 4.986816, 4.986859, 
    4.987047, 0, 4.957404, 4.958957, 4.961073, 4.96328, 4.965307, 4.962757, 
    4.96076, 4.958724, 4.957712, 4.957599, 4.958509, 4.960382, 4.963464, 
    4.966908, 4.971419, 4.972058, 4.973106, 4.974591, 4.9765, 4.978821, 
    4.981529, 4.984586, 4.987936, 4.991505, 4.995192, 4.998876, 5.002409, 
    5.00561, 5.008269, 5.010154, 5.011004, 5.010548, 5.008529, 5.004719,
  // momentumX(26,24, 0-49)
    4.985459, 4.986189, 4.98672, 4.987087, 4.98732, 4.987445, 4.987481, 
    4.987444, 4.987351, 4.987216, 4.987059, 4.986901, 4.986779, 4.986742, 
    4.986866, 0, 4.954684, 4.956232, 4.958356, 4.960571, 4.962602, 4.959841, 
    4.957701, 4.955566, 4.954525, 4.954449, 4.955456, 4.957479, 4.960763, 
    4.964447, 4.969274, 4.970074, 4.971316, 4.973023, 4.975178, 4.977761, 
    4.980742, 4.984078, 4.98771, 4.991553, 4.995505, 4.999441, 5.003209, 
    5.006629, 5.009492, 5.011566, 5.012599, 5.012326, 5.010496, 5.006893,
  // momentumX(26,25, 0-49)
    4.987332, 4.987795, 4.988081, 4.988227, 4.98826, 4.988207, 4.988082, 
    4.987899, 4.987672, 4.987413, 4.98714, 4.986873, 4.986648, 4.986516, 
    4.986553, 0, 4.952617, 4.954093, 4.956138, 4.958269, 4.960216, 4.957344, 
    4.955132, 4.95296, 4.95192, 4.951881, 4.952963, 4.955096, 4.958523, 
    4.962382, 4.96742, 4.968424, 4.96989, 4.971837, 4.974241, 4.977078, 
    4.980317, 4.983906, 4.987782, 4.991862, 4.996039, 5.000186, 5.004151, 
    5.007753, 5.010787, 5.013021, 5.014207, 5.014087, 5.012415, 5.008984,
  // momentumX(26,26, 0-49)
    4.989085, 4.989303, 4.989362, 4.989299, 4.989142, 4.988912, 4.988623, 
    4.988289, 4.987917, 4.98752, 4.987116, 4.986723, 4.986379, 4.986131, 
    4.986053, 0, 4.951242, 4.952576, 4.954455, 4.95641, 4.958189, 4.955317, 
    4.953111, 4.950973, 4.949968, 4.949975, 4.951116, 4.953321, 4.956832, 
    4.960795, 4.965936, 4.967187, 4.96891, 4.971114, 4.973774, 4.976858, 
    4.980333, 4.984146, 4.988233, 4.992505, 4.996861, 5.001172, 5.005288, 
    5.009029, 5.012194, 5.014551, 5.015856, 5.015856, 5.014309, 5.011011,
  // momentumX(26,27, 0-49)
    4.990705, 4.990705, 4.990558, 4.990302, 4.989961, 4.989553, 4.989096, 
    4.988595, 4.988062, 4.987507, 4.986948, 4.986408, 4.985921, 4.985535, 
    4.985317, 0, 4.950675, 4.9518, 4.953434, 4.955128, 4.956655, 4.953875, 
    4.951737, 4.949679, 4.948724, 4.948766, 4.949928, 4.952152, 4.955673, 
    4.959657, 4.964782, 4.966302, 4.968293, 4.970756, 4.97366, 4.976973, 
    4.980659, 4.984664, 4.988923, 4.993354, 4.997853, 5.002294, 5.00653, 
    5.010384, 5.013654, 5.016113, 5.017517, 5.017615, 5.016166, 5.012967,
  // momentumX(26,28, 0-49)
    4.992178, 4.991997, 4.991673, 4.991239, 4.990721, 4.990136, 4.989495, 
    4.988809, 4.988087, 4.987344, 4.9866, 4.985881, 4.985225, 4.984678, 
    4.984301, 0, 4.951277, 4.95214, 4.953459, 4.954813, 4.956015, 4.953386, 
    4.95134, 4.949368, 4.948436, 4.948458, 4.949565, 4.951716, 4.955142, 
    4.959041, 4.964017, 4.965793, 4.968029, 4.970719, 4.973828, 4.977328, 
    4.981176, 4.985326, 4.989712, 4.994259, 4.998865, 5.003407, 5.007742, 
    5.011695, 5.015062, 5.017617, 5.019115, 5.019303, 5.017936, 5.014811,
  // momentumX(26,29, 0-49)
    4.993492, 4.993173, 4.992706, 4.992117, 4.991431, 4.990662, 4.989821, 
    4.98892, 4.987972, 4.987, 4.986029, 4.985097, 4.984242, 4.98352, 
    4.982977, 0, 4.952824, 4.953395, 4.954348, 4.955293, 4.95609, 4.953598, 
    4.951597, 4.949647, 4.948653, 4.948557, 4.949506, 4.951476, 4.95469, 
    4.958384, 4.963066, 4.965036, 4.967458, 4.970321, 4.97359, 4.977238, 
    4.981226, 4.985511, 4.990031, 4.994714, 4.999458, 5.004147, 5.00863, 
    5.012733, 5.016247, 5.018942, 5.020564, 5.020856, 5.019571, 5.016503,
  // momentumX(26,30, 0-49)
    4.99386, 4.992723, 4.991463, 4.990121, 4.988725, 4.987293, 4.985828, 
    4.984329, 4.982784, 4.98118, 4.979504, 4.977741, 4.975895, 4.973988, 
    4.972077, 4.969747, 4.956999, 4.956827, 4.957161, 4.957656, 4.958186, 
    4.95614, 4.954606, 4.953129, 4.952481, 4.952558, 4.953475, 4.955208, 
    4.957977, 4.961077, 4.964963, 4.966609, 4.968697, 4.971236, 4.974212, 
    4.977611, 4.981407, 4.985562, 4.990018, 4.994699, 4.999503, 5.004301, 
    5.008934, 5.013212, 5.016919, 5.019805, 5.021607, 5.022055, 5.020894, 
    5.017915,
  // momentumX(26,31, 0-49)
    4.994776, 4.99362, 4.992315, 4.990895, 4.989389, 4.987814, 4.986178, 
    4.984484, 4.982728, 4.980905, 4.979011, 4.977039, 4.974996, 4.972894, 
    4.97077, 4.969105, 4.957089, 4.956472, 4.956341, 4.956375, 4.956476, 
    4.954564, 4.953073, 4.951636, 4.950986, 4.951061, 4.95199, 4.953743, 
    4.956496, 4.959546, 4.963222, 4.965158, 4.96754, 4.970372, 4.973639, 
    4.977323, 4.981398, 4.985823, 4.99054, 4.995468, 5.000506, 5.005515, 
    5.010334, 5.014765, 5.01858, 5.021528, 5.023334, 5.023723, 5.022443, 
    5.01929,
  // momentumX(26,32, 0-49)
    4.995375, 4.994205, 4.99286, 4.991376, 4.989777, 4.988082, 4.986303, 
    4.984447, 4.982514, 4.980509, 4.978431, 4.976282, 4.974068, 4.971794, 
    4.969482, 4.968209, 4.95724, 4.956205, 4.955632, 4.955235, 4.954943, 
    4.953212, 4.951815, 4.950471, 4.949865, 4.949964, 4.950908, 4.952662, 
    4.955353, 4.958293, 4.961698, 4.963876, 4.966497, 4.969563, 4.973063, 
    4.976978, 4.981282, 4.985934, 4.990874, 4.996023, 5.001267, 5.006473, 
    5.011462, 5.016034, 5.019948, 5.022943, 5.024738, 5.025053, 5.023633, 
    5.020279,
  // momentumX(26,33, 0-49)
    4.995639, 4.99447, 4.9931, 4.991568, 4.989897, 4.988105, 4.98621, 
    4.984221, 4.982143, 4.979988, 4.97776, 4.975465, 4.973111, 4.970702, 
    4.968242, 4.967098, 4.957392, 4.955994, 4.955024, 4.954244, 4.95361, 
    4.952107, 4.950858, 4.949664, 4.949143, 4.949293, 4.950252, 4.951982, 
    4.954559, 4.957333, 4.960416, 4.962787, 4.965594, 4.96884, 4.972515, 
    4.976605, 4.981087, 4.985918, 4.991039, 4.996368, 5.001789, 5.007158, 
    5.012293, 5.01698, 5.020972, 5.023992, 5.025752, 5.025967, 5.02438, 
    5.020803,
  // momentumX(26,34, 0-49)
    4.995543, 4.994396, 4.993027, 4.99147, 4.98975, 4.98789, 4.985905, 
    4.983811, 4.98162, 4.979345, 4.976997, 4.97459, 4.97213, 4.969624, 
    4.967066, 4.965834, 4.957517, 4.955821, 4.954513, 4.953405, 4.952485, 
    4.951245, 4.95019, 4.9492, 4.948807, 4.949031, 4.950005, 4.951681, 
    4.954097, 4.956656, 4.959386, 4.961906, 4.964849, 4.968222, 4.972019, 
    4.97623, 4.980836, 4.985796, 4.991051, 4.996513, 5.002068, 5.007562, 
    5.012805, 5.017571, 5.021602, 5.024612, 5.026301, 5.026382, 5.024599, 
    5.020772,
  // momentumX(26,35, 0-49)
    4.995066, 4.99397, 4.992628, 4.991074, 4.989336, 4.987434, 4.985391, 
    4.983224, 4.98095, 4.978586, 4.976151, 4.97366, 4.971129, 4.968563, 
    4.965956, 4.964484, 4.957617, 4.955689, 4.954103, 4.952727, 4.951577, 
    4.950626, 4.949806, 4.949069, 4.948839, 4.949157, 4.950138, 4.951736, 
    4.953943, 4.956252, 4.958614, 4.961243, 4.964278, 4.967728, 4.971596, 
    4.975876, 4.980554, 4.985588, 4.990923, 4.996468, 5.002102, 5.007667, 
    5.012964, 5.017759, 5.02178, 5.024729, 5.026304, 5.026208, 5.024194, 
    5.02009,
  // momentumX(26,36, 0-49)
    4.99419, 4.993175, 4.991889, 4.99037, 4.988643, 4.986734, 4.984667, 
    4.98246, 4.980136, 4.977716, 4.975226, 4.972688, 4.970117, 4.967527, 
    4.964915, 4.96312, 4.957703, 4.95561, 4.953803, 4.952217, 4.950887, 
    4.950241, 4.949687, 4.949242, 4.949209, 4.949636, 4.95062, 4.952115, 
    4.954077, 4.95611, 4.958105, 4.960808, 4.963894, 4.967376, 4.971268, 
    4.975566, 4.98026, 4.985313, 4.990666, 4.996232, 5.001882, 5.007453, 
    5.012741, 5.017495, 5.021441, 5.024268, 5.025669, 5.02535, 5.023067, 
    5.018667,
  // momentumX(26,37, 0-49)
    4.992908, 4.991998, 4.9908, 4.989348, 4.987668, 4.985786, 4.983728, 
    4.981519, 4.979182, 4.976744, 4.974233, 4.971678, 4.969099, 4.966518, 
    4.963937, 4.961798, 4.957793, 4.955594, 4.953619, 4.951871, 4.950411, 
    4.950073, 4.949806, 4.949687, 4.949876, 4.950426, 4.951407, 4.952781, 
    4.954471, 4.956215, 4.957856, 4.9606, 4.963703, 4.967181, 4.971049, 
    4.975317, 4.979972, 4.984982, 4.990291, 4.995806, 5.001399, 5.006898, 
    5.012094, 5.01673, 5.020518, 5.023149, 5.024311, 5.023713, 5.021127, 
    5.016415,
  // momentumX(26,38, 0-49)
    4.991222, 4.990443, 4.98936, 4.988006, 4.986406, 4.984589, 4.98258, 
    4.980407, 4.978095, 4.975675, 4.97318, 4.970641, 4.968087, 4.965544, 
    4.963021, 4.960566, 4.957904, 4.955646, 4.953547, 4.951684, 4.950138, 
    4.950104, 4.950134, 4.950362, 4.950793, 4.951478, 4.952455, 4.953692, 
    4.955092, 4.956546, 4.957858, 4.960621, 4.96371, 4.967146, 4.970952, 
    4.975142, 4.979702, 4.98461, 4.989802, 4.995189, 5.000639, 5.005978, 
    5.010987, 5.015409, 5.01895, 5.021299, 5.022146, 5.021213, 5.018287, 
    5.013258,
  // momentumX(26,39, 0-49)
    4.989146, 4.988517, 4.987576, 4.98635, 4.984865, 4.983149, 4.981227, 
    4.979128, 4.976882, 4.974522, 4.972079, 4.969591, 4.967091, 4.96461, 
    4.962165, 4.959454, 4.95805, 4.955768, 4.953585, 4.951646, 4.950048, 
    4.950306, 4.950636, 4.951224, 4.951909, 4.952735, 4.953708, 4.954801, 
    4.955904, 4.957078, 4.958095, 4.960857, 4.963908, 4.967274, 4.970981, 
    4.975045, 4.979459, 4.984196, 4.9892, 4.994374, 4.999588, 5.004664, 
    5.009383, 5.013483, 5.016672, 5.018644, 5.019099, 5.017773, 5.014479, 
    5.009132,
  // momentumX(26,40, 0-49)
    4.986707, 4.986245, 4.985466, 4.984396, 4.983058, 4.981478, 4.979682, 
    4.977698, 4.975558, 4.973294, 4.970941, 4.968537, 4.966121, 4.963724, 
    4.961371, 4.958483, 4.95824, 4.95596, 4.953722, 4.951737, 4.950122, 
    4.950653, 4.951275, 4.952221, 4.953166, 4.954142, 4.955109, 4.956059, 
    4.956869, 4.957781, 4.958541, 4.961287, 4.964283, 4.967553, 4.97113, 
    4.975026, 4.979239, 4.983742, 4.988476, 4.993349, 4.998224, 5.002929, 
    5.007241, 5.010903, 5.013631, 5.015126, 5.015107, 5.013333, 5.009647, 
    5.004004,
  // momentumX(26,41, 0-49)
    4.983946, 4.983662, 4.983064, 4.982172, 4.981009, 4.979598, 4.977962, 
    4.976132, 4.974137, 4.972007, 4.969779, 4.967493, 4.965187, 4.962894, 
    4.960647, 4.957664, 4.958471, 4.956212, 4.953946, 4.951943, 4.950333, 
    4.951114, 4.952014, 4.953312, 4.954513, 4.955637, 4.9566, 4.957409, 
    4.957942, 4.95862, 4.959163, 4.961884, 4.964809, 4.967964, 4.97138, 
    4.97507, 4.97903, 4.983232, 4.987618, 4.992094, 4.996525, 5.000741, 
    5.004525, 5.007628, 5.009777, 5.010693, 5.010121, 5.007853, 5.003766, 
    4.997855,
  // momentumX(26,42, 0-49)
    4.980917, 4.980814, 4.98041, 4.979715, 4.978751, 4.977537, 4.976097, 
    4.974453, 4.972636, 4.970678, 4.968611, 4.966472, 4.964302, 4.962132, 
    4.959999, 4.957001, 4.958748, 4.95652, 4.954246, 4.952245, 4.950657, 
    4.95166, 4.952818, 4.954448, 4.955894, 4.957162, 4.958123, 4.958803, 
    4.95908, 4.959553, 4.959918, 4.962606, 4.965451, 4.968475, 4.971704, 
    4.97515, 4.978807, 4.982642, 4.986598, 4.990582, 4.994461, 4.998068, 
    5.0012, 5.003619, 5.005074, 5.005314, 5.004117, 5.001315, 4.996832, 
    4.990704,
  // momentumX(26,43, 0-49)
    4.977679, 4.97776, 4.977554, 4.977072, 4.976327, 4.975336, 4.974116, 
    4.972692, 4.971086, 4.969328, 4.967451, 4.965489, 4.963478, 4.961449, 
    4.959437, 4.956493, 4.959065, 4.956875, 4.954607, 4.952624, 4.951071, 
    4.952264, 4.953651, 4.955585, 4.95726, 4.958661, 4.959623, 4.960185, 
    4.960233, 4.960534, 4.960759, 4.963408, 4.966163, 4.96904, 4.97206, 
    4.975228, 4.978531, 4.981936, 4.985381, 4.988777, 4.991995, 4.994875, 
    4.99723, 4.998845, 4.999496, 4.998971, 4.997089, 4.993732, 4.988872, 
    4.982594,
  // momentumX(26,44, 0-49)
    4.974301, 4.974561, 4.974557, 4.974297, 4.973784, 4.973035, 4.972059, 
    4.970877, 4.96951, 4.967981, 4.966322, 4.964559, 4.962726, 4.960854, 
    4.958971, 4.956134, 4.959414, 4.957269, 4.955017, 4.953065, 4.951551, 
    4.952901, 4.954484, 4.956686, 4.958561, 4.960083, 4.961043, 4.961501, 
    4.961351, 4.961507, 4.961627, 4.964231, 4.966889, 4.969604, 4.972392, 
    4.975247, 4.97815, 4.981063, 4.983919, 4.986634, 4.989085, 4.991127, 
    4.992589, 4.993289, 4.99304, 4.991673, 4.989062, 4.985146, 4.979949, 
    4.973607,
  // momentumX(26,45, 0-49)
    4.970855, 4.971286, 4.971483, 4.971446, 4.971176, 4.970679, 4.969965, 
    4.969045, 4.967938, 4.96666, 4.965239, 4.963696, 4.962062, 4.960358, 
    4.958611, 4.955917, 4.95979, 4.957693, 4.955468, 4.95355, 4.952076, 
    4.95355, 4.955291, 4.957713, 4.959756, 4.961379, 4.962333, 4.9627, 
    4.962382, 4.962423, 4.96246, 4.965011, 4.967559, 4.970098, 4.972632, 
    4.97514, 4.977598, 4.979958, 4.982154, 4.984101, 4.985687, 4.986785, 
    4.987253, 4.986942, 4.985713, 4.983451, 4.980091, 4.975633, 4.970161, 
    4.963855,
  // momentumX(26,46, 0-49)
    4.967414, 4.968003, 4.968394, 4.968578, 4.968554, 4.968318, 4.967876, 
    4.967232, 4.9664, 4.96539, 4.964222, 4.962915, 4.961491, 4.959968, 
    4.958365, 4.955836, 4.960183, 4.95814, 4.955951, 4.954069, 4.952631, 
    4.954192, 4.956049, 4.95864, 4.960809, 4.962502, 4.963447, 4.963733, 
    4.963276, 4.963221, 4.963187, 4.965672, 4.968098, 4.970442, 4.972695, 
    4.974825, 4.976792, 4.978544, 4.980013, 4.981115, 4.981754, 4.981822, 
    4.98121, 4.979815, 4.977552, 4.974366, 4.970264, 4.965308, 4.959643, 
    4.953489,
  // momentumX(26,47, 0-49)
    4.964046, 4.964777, 4.965352, 4.965752, 4.96597, 4.965997, 4.965829, 
    4.96547, 4.96492, 4.964187, 4.963284, 4.962223, 4.961019, 4.959685, 
    4.958235, 4.955878, 4.960584, 4.958601, 4.956454, 4.954607, 4.953197, 
    4.954808, 4.956738, 4.959435, 4.961684, 4.963416, 4.964339, 4.964552, 
    4.96398, 4.963842, 4.963738, 4.966136, 4.968418, 4.970546, 4.972489, 
    4.974205, 4.975642, 4.976735, 4.977419, 4.977613, 4.977237, 4.976211, 
    4.974462, 4.97194, 4.968619, 4.964515, 4.959707, 4.954324, 4.948567, 
    4.942689,
  // momentumX(26,48, 0-49)
    4.96081, 4.961668, 4.962411, 4.963017, 4.963469, 4.963753, 4.96386, 
    4.963782, 4.963516, 4.963064, 4.962431, 4.961621, 4.960644, 4.959507, 
    4.958216, 4.956029, 4.960979, 4.959066, 4.956965, 4.955151, 4.953761, 
    4.955386, 4.957339, 4.960083, 4.962356, 4.964089, 4.964973, 4.965117, 
    4.964446, 4.964223, 4.964039, 4.966322, 4.968429, 4.970309, 4.971912, 
    4.973177, 4.974042, 4.974437, 4.974288, 4.973528, 4.972093, 4.969935, 
    4.967025, 4.963368, 4.959004, 4.954024, 4.948578, 4.942863, 4.937129, 
    4.93166,
  // momentumX(26,49, 0-49)
    4.957191, 4.958059, 4.958873, 4.959602, 4.960219, 4.9607, 4.961027, 
    4.961179, 4.961144, 4.960912, 4.960473, 4.959821, 4.95895, 4.957851, 
    4.956515, 4.953525, 4.964903, 4.962058, 4.958658, 4.955644, 4.953284, 
    4.956749, 4.960586, 4.965696, 4.969499, 4.971891, 4.972278, 4.970906, 
    4.967642, 4.965106, 4.962541, 4.964893, 4.966942, 4.968615, 4.969858, 
    4.970594, 4.970757, 4.97027, 4.969067, 4.967099, 4.964337, 4.960783, 
    4.956475, 4.951499, 4.945994, 4.940145, 4.934196, 4.928425, 4.923135, 
    4.918625,
  // momentumX(27,0, 0-49)
    4.952485, 4.956017, 4.95919, 4.962013, 4.964487, 4.966623, 4.968421, 
    4.969888, 4.971034, 4.971874, 4.972427, 4.972726, 4.972806, 4.972714, 
    4.972504, 4.972033, 4.971988, 4.9717, 4.971503, 4.971475, 4.971662, 
    4.97227, 4.973104, 4.974205, 4.975557, 4.977133, 4.978898, 4.980816, 
    4.982846, 4.984953, 4.987058, 4.989343, 4.991569, 4.993695, 4.995677, 
    4.997463, 4.998989, 5.00017, 5.000906, 5.001068, 5.000506, 4.999043, 
    4.996487, 4.992639, 4.987311, 4.98035, 4.971671, 4.961278, 4.9493, 
    4.936006,
  // momentumX(27,1, 0-49)
    4.953785, 4.957267, 4.960383, 4.963142, 4.965549, 4.967614, 4.969344, 
    4.970743, 4.971827, 4.97261, 4.973116, 4.973373, 4.973421, 4.973308, 
    4.973083, 4.972408, 4.972571, 4.972211, 4.971914, 4.971784, 4.971873, 
    4.97256, 4.97343, 4.974563, 4.975933, 4.977504, 4.979235, 4.981091, 
    4.983034, 4.985042, 4.987011, 4.989357, 4.991658, 4.993884, 4.995999, 
    4.997962, 4.999713, 5.001177, 5.002253, 5.002817, 5.002716, 5.001765, 
    4.999763, 4.996496, 4.991755, 4.985361, 4.977194, 4.967225, 4.955546, 
    4.942395,
  // momentumX(27,2, 0-49)
    4.9551, 4.958522, 4.961576, 4.964267, 4.96661, 4.96861, 4.970279, 
    4.971625, 4.97266, 4.973405, 4.97388, 4.974118, 4.974155, 4.974039, 
    4.97382, 4.972966, 4.973311, 4.972891, 4.972506, 4.972278, 4.972264, 
    4.973009, 4.97389, 4.975019, 4.976368, 4.9779, 4.979566, 4.981339, 
    4.983176, 4.985064, 4.98687, 4.989237, 4.991573, 4.993855, 4.996058, 
    4.998144, 5.000066, 5.00175, 5.003102, 5.003998, 5.004288, 5.003786, 
    5.002285, 4.999563, 4.995397, 4.989588, 4.981988, 4.972539, 4.961292, 
    4.948447,
  // momentumX(27,3, 0-49)
    4.956424, 4.959782, 4.962767, 4.965392, 4.967669, 4.969612, 4.971227, 
    4.972527, 4.973528, 4.974247, 4.97471, 4.974946, 4.974991, 4.974892, 
    4.974695, 4.973688, 4.974173, 4.973708, 4.973245, 4.972928, 4.972816, 
    4.973597, 4.974463, 4.975552, 4.976844, 4.978302, 4.979884, 4.981561, 
    4.983288, 4.985043, 4.986671, 4.989024, 4.991359, 4.993658, 4.995905, 
    4.99807, 5.000108, 5.001954, 5.003517, 5.004678, 5.00529, 5.005171, 
    5.004114, 5.001892, 4.998278, 4.993056, 4.986063, 4.977203, 4.966496, 
    4.9541,
  // momentumX(27,4, 0-49)
    4.957763, 4.961049, 4.963962, 4.966518, 4.968731, 4.970614, 4.97218, 
    4.973444, 4.974419, 4.975125, 4.975588, 4.975837, 4.975906, 4.975838, 
    4.975676, 4.974549, 4.975114, 4.974617, 4.974098, 4.973704, 4.973499, 
    4.974296, 4.97512, 4.976135, 4.977338, 4.978698, 4.980179, 4.981754, 
    4.983374, 4.984993, 4.986437, 4.988748, 4.991049, 4.993332, 4.995584, 
    4.997785, 4.999891, 5.001845, 5.003561, 5.004924, 5.005792, 5.005991, 
    5.00532, 5.003553, 5.000459, 4.995819, 4.98945, 4.981233, 4.971154, 
    4.959323,
  // momentumX(27,5, 0-49)
    4.959124, 4.96233, 4.965165, 4.967649, 4.969796, 4.971621, 4.973139, 
    4.974367, 4.975321, 4.976024, 4.976496, 4.976768, 4.976871, 4.976844, 
    4.976726, 4.975518, 4.976087, 4.975574, 4.975018, 4.974565, 4.97428, 
    4.975071, 4.975831, 4.976738, 4.977826, 4.979064, 4.980437, 4.981911, 
    4.983433, 4.984925, 4.986189, 4.988428, 4.990667, 4.992902, 4.995128, 
    4.997325, 4.999457, 5.001471, 5.003284, 5.004794, 5.005862, 5.006324, 
    5.005984, 5.004626, 5.002022, 4.997947, 4.992211, 4.984674, 4.975287, 
    4.964118,
  // momentumX(27,6, 0-49)
    4.960515, 4.963633, 4.966385, 4.96879, 4.970866, 4.972629, 4.974098, 
    4.975291, 4.976225, 4.976924, 4.97741, 4.977711, 4.977855, 4.977876, 
    4.977808, 4.976558, 4.977046, 4.976531, 4.97596, 4.975471, 4.975124, 
    4.975888, 4.976562, 4.977334, 4.978279, 4.979381, 4.980637, 4.982016, 
    4.983459, 4.984834, 4.985934, 4.988077, 4.990227, 4.992387, 4.994555, 
    4.996716, 4.998837, 5.000868, 5.002738, 5.004347, 5.005566, 5.006243, 
    5.006188, 5.005199, 5.003053, 4.999527, 4.994426, 4.987591, 4.978942, 
    4.968504,
  // momentumX(27,7, 0-49)
    4.961944, 4.964969, 4.96763, 4.969948, 4.971945, 4.97364, 4.975054, 
    4.976207, 4.977119, 4.977812, 4.978312, 4.978641, 4.978827, 4.978899, 
    4.97888, 4.977633, 4.977947, 4.977446, 4.976884, 4.976382, 4.975995, 
    4.976711, 4.97728, 4.977891, 4.978675, 4.97963, 4.980768, 4.982057, 
    4.98344, 4.984717, 4.985673, 4.987694, 4.989734, 4.991795, 4.99388, 
    4.995977, 4.998057, 5.000075, 5.001965, 5.003634, 5.004968, 5.005818, 
    5.006014, 5.00536, 5.003646, 5.000652, 4.996178, 4.990054, 4.982172, 
    4.972516,
  // momentumX(27,8, 0-49)
    4.96342, 4.966343, 4.968904, 4.971127, 4.973035, 4.974654, 4.976002, 
    4.977108, 4.977989, 4.978671, 4.979177, 4.979532, 4.979758, 4.979877, 
    4.979905, 4.978708, 4.978746, 4.978274, 4.97775, 4.977262, 4.976861, 
    4.977507, 4.977953, 4.978384, 4.978992, 4.979788, 4.980811, 4.982022, 
    4.983364, 4.984567, 4.985405, 4.987285, 4.989192, 4.991133, 4.993113, 
    4.995123, 4.997139, 4.999117, 5.001001, 5.002707, 5.004125, 5.005124, 
    5.005543, 5.005198, 5.003892, 5.001414, 4.997559, 4.992144, 4.985043, 
    4.976196,
  // momentumX(27,9, 0-49)
    4.964952, 4.967762, 4.970212, 4.972329, 4.974138, 4.975667, 4.976941, 
    4.977984, 4.978825, 4.979486, 4.97999, 4.980362, 4.98062, 4.980781, 
    4.980847, 4.979746, 4.979405, 4.97898, 4.978518, 4.978075, 4.977688, 
    4.978245, 4.978553, 4.978786, 4.97921, 4.979844, 4.980752, 4.981893, 
    4.983215, 4.984366, 4.985122, 4.98684, 4.988597, 4.990402, 4.992261, 
    4.994167, 4.9961, 4.998025, 4.999886, 5.001608, 5.003094, 5.004222, 
    5.004846, 5.004794, 5.003879, 5.001898, 4.998647, 4.993936, 4.987614, 
    4.979589,
  // momentumX(27,10, 0-49)
    4.966544, 4.969228, 4.971554, 4.973551, 4.975248, 4.976675, 4.977859, 
    4.97883, 4.979616, 4.980243, 4.980734, 4.981112, 4.98139, 4.981582, 
    4.981678, 4.980717, 4.979891, 4.979529, 4.979159, 4.978791, 4.978449, 
    4.978896, 4.979054, 4.97908, 4.979313, 4.979784, 4.980581, 4.981661, 
    4.982981, 4.984105, 4.984818, 4.986358, 4.987952, 4.989606, 4.991331, 
    4.993123, 4.994964, 4.996823, 4.998651, 5.000382, 5.001927, 5.003174, 
    5.003991, 5.00422, 5.003681, 5.002182, 4.999519, 4.995496, 4.989943, 
    4.982737,
  // momentumX(27,11, 0-49)
    4.968184, 4.970732, 4.972922, 4.974787, 4.976358, 4.97767, 4.978752, 
    4.979636, 4.980354, 4.980931, 4.981393, 4.981763, 4.982052, 4.982261, 
    4.982378, 4.981594, 4.980174, 4.979899, 4.979648, 4.979387, 4.979123, 
    4.979436, 4.979437, 4.979248, 4.979291, 4.979603, 4.980292, 4.981318, 
    4.98265, 4.983774, 4.984485, 4.985836, 4.987253, 4.988749, 4.990333, 
    4.992004, 4.993749, 4.995539, 4.997333, 4.99907, 5.000671, 5.002034, 
    5.00304, 5.00354, 5.003365, 5.00233, 5.000237, 4.996881, 4.992076, 
    4.985673,
  // momentumX(27,12, 0-49)
    4.969869, 4.972264, 4.974305, 4.976025, 4.977458, 4.978641, 4.979606, 
    4.98039, 4.981024, 4.981538, 4.981959, 4.982306, 4.982589, 4.982803, 
    4.982933, 4.982355, 4.980234, 4.98007, 4.979968, 4.979845, 4.979689, 
    4.97985, 4.979685, 4.979283, 4.979139, 4.979298, 4.979885, 4.980863, 
    4.982218, 4.983363, 4.984119, 4.985269, 4.986504, 4.987836, 4.989278, 
    4.990828, 4.992476, 4.9942, 4.995962, 4.997709, 4.999368, 5.000849, 
    5.002039, 5.002804, 5.002984, 5.002398, 5.00085, 4.998134, 4.99405, 
    4.988423,
  // momentumX(27,13, 0-49)
    4.971578, 4.973805, 4.975684, 4.977247, 4.978529, 4.979571, 4.980408, 
    4.98108, 4.981618, 4.982056, 4.982419, 4.982728, 4.982991, 4.983199, 
    4.983337, 4.982982, 4.980053, 4.980028, 4.980104, 4.980148, 4.980134, 
    4.980123, 4.97979, 4.979178, 4.978858, 4.978872, 4.979362, 4.980295, 
    4.981681, 4.982868, 4.983716, 4.984661, 4.98571, 4.986878, 4.988178, 
    4.989611, 4.991169, 4.992833, 4.994571, 4.996334, 4.998056, 4.999658, 
    5.001034, 5.002057, 5.002578, 5.002422, 5.001395, 4.999288, 4.995888, 
    4.991003,
  // momentumX(27,14, 0-49)
    4.973285, 4.975332, 4.977035, 4.978428, 4.979551, 4.980443, 4.981143, 
    4.981692, 4.982125, 4.982474, 4.982768, 4.983025, 4.983253, 4.983449, 
    4.983591, 4.983465, 4.979623, 4.979764, 4.980047, 4.980291, 4.980448, 
    4.980245, 4.979743, 4.978934, 4.978452, 4.978334, 4.978735, 4.979624, 
    4.981044, 4.98229, 4.983274, 4.984014, 4.98488, 4.985888, 4.987052, 
    4.988374, 4.98985, 4.991462, 4.993183, 4.994971, 4.996765, 4.998491, 
    5.000052, 5.001328, 5.002178, 5.002431, 5.001897, 5.000363, 4.99761, 
    4.993423,
  // momentumX(27,15, 0-49)
    4.974969, 4.976818, 4.97833, 4.979544, 4.980499, 4.981234, 4.981791, 
    4.982209, 4.982529, 4.98278, 4.982994, 4.983189, 4.983375, 4.983549, 
    4.983696, 4.983794, 4.978942, 4.979278, 4.979795, 4.980265, 4.98062, 
    4.980211, 4.979545, 4.978554, 4.977929, 4.977694, 4.978014, 4.978863, 
    4.980318, 4.981638, 4.982798, 4.983336, 4.984023, 4.984879, 4.985915, 
    4.987135, 4.988539, 4.990111, 4.991827, 4.993648, 4.99552, 4.997373, 
    4.999117, 5.000638, 5.001802, 5.002442, 5.002368, 5.00137, 4.999219, 
    4.995688,
  // momentumX(27,16, 0-49)
    4.9766, 4.978232, 4.979541, 4.980565, 4.981343, 4.981917, 4.982327, 
    4.982615, 4.982817, 4.982967, 4.983095, 4.98322, 4.983356, 4.983504, 
    4.983661, 4.983968, 4.978021, 4.978576, 4.979346, 4.980065, 4.980643, 
    4.980015, 4.979194, 4.97804, 4.977294, 4.976964, 4.977215, 4.978029, 
    4.979517, 4.980919, 4.982292, 4.982636, 4.983153, 4.983865, 4.984783, 
    4.985914, 4.987255, 4.988797, 4.990517, 4.992379, 4.994334, 4.996316, 
    4.99824, 4.999999, 5.001459, 5.002461, 5.002818, 5.002316, 5.000722, 
    4.997799,
  // momentumX(27,17, 0-49)
    4.97815, 4.979545, 4.980634, 4.981458, 4.982053, 4.982463, 4.982728, 
    4.982884, 4.982973, 4.983024, 4.983063, 4.983118, 4.983199, 4.983321, 
    4.983489, 4.983988, 4.976887, 4.977677, 4.978717, 4.979698, 4.980515, 
    4.97966, 4.978692, 4.977397, 4.976559, 4.976156, 4.976355, 4.977139, 
    4.97866, 4.980151, 4.981763, 4.981924, 4.982281, 4.982859, 4.983669, 
    4.98472, 4.986009, 4.987531, 4.989263, 4.991172, 4.993215, 4.995326, 
    4.997425, 4.999409, 5.001151, 5.00249, 5.003245, 5.0032, 5.002119, 
    4.999754,
  // momentumX(27,18, 0-49)
    4.979592, 4.980724, 4.981576, 4.982186, 4.982595, 4.982841, 4.982964, 
    4.983, 4.982983, 4.982941, 4.9829, 4.982886, 4.982915, 4.983007, 
    4.983186, 4.983865, 4.975588, 4.976619, 4.977927, 4.979177, 4.980241, 
    4.979152, 4.978045, 4.976635, 4.97573, 4.975284, 4.975449, 4.976212, 
    4.977769, 4.979352, 4.981221, 4.981211, 4.981418, 4.981871, 4.982583, 
    4.983562, 4.984807, 4.986314, 4.988064, 4.990025, 4.992156, 4.994394, 
    4.996664, 4.998864, 5.000867, 5.002522, 5.003644, 5.004018, 5.003407, 
    5.001557,
  // momentumX(27,19, 0-49)
    4.980903, 4.98174, 4.98233, 4.982714, 4.982932, 4.983019, 4.98301, 
    4.982938, 4.982831, 4.982711, 4.982603, 4.982526, 4.982506, 4.982572, 
    4.982763, 4.983617, 4.9742, 4.975467, 4.977031, 4.978539, 4.979841, 
    4.978513, 4.97728, 4.975773, 4.974828, 4.974364, 4.974518, 4.975278, 
    4.976873, 4.978549, 4.980679, 4.98051, 4.980577, 4.980914, 4.981531, 
    4.982439, 4.983643, 4.985138, 4.986907, 4.988921, 4.991139, 4.993503, 
    4.995936, 4.998341, 5.000593, 5.002542, 5.004004, 5.004765, 5.004586, 
    5.00321,
  // momentumX(27,20, 0-49)
    4.982862, 4.984146, 4.985185, 4.986007, 4.98664, 4.987111, 4.987448, 
    4.987677, 4.987826, 4.987921, 4.987986, 4.988048, 4.988135, 4.988278, 
    4.988526, 0, 4.972143, 4.973258, 4.97473, 4.976183, 4.977445, 4.975578, 
    4.973876, 4.971932, 4.970649, 4.969963, 4.970038, 4.970872, 4.97272, 
    4.974809, 4.977582, 4.977671, 4.978006, 4.978611, 4.979485, 4.980634, 
    4.982059, 4.983755, 4.985709, 4.987898, 4.990287, 4.992825, 4.995441, 
    4.998047, 5.000524, 5.002726, 5.004475, 5.005559, 5.005739, 5.004762,
  // momentumX(27,21, 0-49)
    4.984021, 4.985055, 4.985878, 4.986519, 4.987, 4.98735, 4.987592, 
    4.987746, 4.987836, 4.987881, 4.987903, 4.987926, 4.987977, 4.98809, 
    4.988317, 0, 4.96787, 4.969113, 4.970778, 4.972454, 4.973938, 4.971829, 
    4.970017, 4.96804, 4.966849, 4.966359, 4.966709, 4.967876, 4.970111, 
    4.97262, 4.975931, 4.976147, 4.976643, 4.977433, 4.978511, 4.979876, 
    4.981517, 4.983426, 4.985584, 4.987966, 4.990533, 4.993235, 4.996002, 
    4.998747, 5.001359, 5.003693, 5.005579, 5.006813, 5.007162, 5.006378,
  // momentumX(27,22, 0-49)
    4.9851, 4.985905, 4.986529, 4.987001, 4.987345, 4.987583, 4.987735, 
    4.987818, 4.987849, 4.987846, 4.987824, 4.987807, 4.987818, 4.987895, 
    4.988095, 0, 4.96427, 4.965615, 4.967438, 4.969296, 4.970961, 4.968601, 
    4.96665, 4.964593, 4.963428, 4.963049, 4.963583, 4.964988, 4.96751, 
    4.970334, 4.974064, 4.974349, 4.974948, 4.975873, 4.977114, 4.978661, 
    4.980502, 4.982621, 4.984995, 4.987593, 4.990371, 4.993275, 4.996236, 
    4.999167, 5.001956, 5.004463, 5.006518, 5.007926, 5.008459, 5.007876,
  // momentumX(27,23, 0-49)
    4.986108, 4.986693, 4.987132, 4.98745, 4.987665, 4.987799, 4.987868, 
    4.987884, 4.987857, 4.987806, 4.987741, 4.98768, 4.987649, 4.987686, 
    4.987846, 0, 4.961174, 4.962575, 4.964491, 4.966458, 4.968225, 4.965626, 
    4.963521, 4.961361, 4.960176, 4.959849, 4.960501, 4.962069, 4.964801, 
    4.96786, 4.971903, 4.972238, 4.972919, 4.973962, 4.97535, 4.977074, 
    4.979115, 4.981455, 4.984063, 4.986903, 4.989927, 4.993075, 4.996275, 
    4.999434, 5.00244, 5.005151, 5.007399, 5.008994, 5.009711, 5.00932,
  // momentumX(27,24, 0-49)
    4.987052, 4.987432, 4.987696, 4.987866, 4.987962, 4.987997, 4.987984, 
    4.987933, 4.987851, 4.98775, 4.987639, 4.987533, 4.987454, 4.987441, 
    4.987548, 0, 4.958886, 4.960289, 4.962229, 4.964231, 4.966028, 4.963264, 
    4.961052, 4.958817, 4.957613, 4.957313, 4.958032, 4.959703, 4.962571, 
    4.965787, 4.970043, 4.970445, 4.971216, 4.972371, 4.973891, 4.975769, 
    4.977979, 4.980506, 4.983313, 4.986362, 4.989601, 4.992966, 4.996381, 
    4.99975, 5.002959, 5.005866, 5.0083, 5.010072, 5.010966, 5.010753,
  // momentumX(27,25, 0-49)
    4.987951, 4.988135, 4.988231, 4.988259, 4.988237, 4.988174, 4.98808, 
    4.987959, 4.987818, 4.987662, 4.987497, 4.987339, 4.987206, 4.987133, 
    4.987175, 0, 4.957164, 4.958512, 4.960404, 4.962363, 4.964118, 4.961286, 
    4.959035, 4.956786, 4.955588, 4.955317, 4.956082, 4.957819, 4.960765, 
    4.964076, 4.968446, 4.968953, 4.969841, 4.971123, 4.972783, 4.974807, 
    4.977177, 4.979869, 4.98285, 4.986078, 4.989499, 4.993052, 4.996652, 
    5.000207, 5.003596, 5.006678, 5.009283, 5.011218, 5.01227, 5.012215,
  // momentumX(27,26, 0-49)
    4.988813, 4.988812, 4.98875, 4.988639, 4.9885, 4.988336, 4.988153, 
    4.987953, 4.987741, 4.987518, 4.98729, 4.987069, 4.986872, 4.986731, 
    4.986691, 0, 4.956017, 4.957257, 4.959034, 4.960871, 4.962512, 4.95972, 
    4.957509, 4.955312, 4.954154, 4.953917, 4.954714, 4.956479, 4.959447, 
    4.962788, 4.967175, 4.967828, 4.968863, 4.970294, 4.972103, 4.974275, 
    4.976792, 4.979629, 4.982756, 4.986129, 4.989699, 4.9934, 4.997152, 
    5.000857, 5.004397, 5.007628, 5.010381, 5.01246, 5.013651, 5.013734,
  // momentumX(27,27, 0-49)
    4.98965, 4.989479, 4.989264, 4.98902, 4.988759, 4.988484, 4.9882, 
    4.987906, 4.987603, 4.987295, 4.986986, 4.986688, 4.986415, 4.986197, 
    4.986067, 0, 4.955529, 4.956617, 4.958216, 4.959864, 4.961324, 4.958663, 
    4.956551, 4.954452, 4.95335, 4.953136, 4.95393, 4.955672, 4.958594, 
    4.961887, 4.966184, 4.967004, 4.968203, 4.969788, 4.971744, 4.974054, 
    4.976701, 4.979663, 4.98291, 4.986403, 4.990092, 4.993917, 4.997795, 
    5.001633, 5.005309, 5.008677, 5.011567, 5.013782, 5.015105, 5.01531,
  // momentumX(27,28, 0-49)
    4.990469, 4.990145, 4.989788, 4.989411, 4.989022, 4.988625, 4.988218, 
    4.987805, 4.987385, 4.986967, 4.986554, 4.98616, 4.985801, 4.9855, 
    4.985283, 0, 4.956028, 4.956934, 4.958307, 4.959707, 4.96093, 4.958463, 
    4.956476, 4.954484, 4.953412, 4.953169, 4.953884, 4.955516, 4.958292, 
    4.961439, 4.965523, 4.966502, 4.967848, 4.969568, 4.971642, 4.974057, 
    4.976798, 4.979848, 4.983181, 4.986762, 4.990545, 4.994473, 4.998466, 
    5.002428, 5.006239, 5.009749, 5.012783, 5.015139, 5.016596, 5.016923,
  // momentumX(27,29, 0-49)
    4.991272, 4.99082, 4.990334, 4.989828, 4.989304, 4.988763, 4.988209, 
    4.987643, 4.987072, 4.986504, 4.985958, 4.985448, 4.984994, 4.984619, 
    4.984338, 0, 4.957261, 4.957983, 4.959101, 4.960205, 4.96113, 4.958851, 
    4.956955, 4.955013, 4.953891, 4.953528, 4.954064, 4.955482, 4.958002, 
    4.960886, 4.964627, 4.965713, 4.967158, 4.968967, 4.971126, 4.973623, 
    4.976449, 4.979589, 4.983022, 4.986718, 4.990633, 4.994709, 4.998869, 
    5.003012, 5.00701, 5.010713, 5.013935, 5.016467, 5.018081, 5.018536,
  // momentumX(27,30, 0-49)
    4.991342, 4.990104, 4.98886, 4.987627, 4.986415, 4.985223, 4.984044, 
    4.982868, 4.981678, 4.980457, 4.979197, 4.977892, 4.976555, 4.975228, 
    4.973989, 4.972118, 4.961142, 4.961493, 4.962195, 4.962931, 4.963588, 
    4.961671, 4.96014, 4.958567, 4.957699, 4.957439, 4.957901, 4.95906, 
    4.961126, 4.963423, 4.966387, 4.96713, 4.968222, 4.969685, 4.971525, 
    4.973748, 4.976355, 4.979339, 4.982685, 4.986363, 4.990328, 4.994513, 
    4.998833, 5.003178, 5.007408, 5.011355, 5.014824, 5.017593, 5.019419, 
    5.020052,
  // momentumX(27,31, 0-49)
    4.992085, 4.990796, 4.989485, 4.988165, 4.986845, 4.985525, 4.9842, 
    4.982865, 4.981511, 4.980129, 4.978714, 4.977267, 4.975796, 4.974329, 
    4.972923, 4.971511, 4.96095, 4.960932, 4.961246, 4.961601, 4.961905, 
    4.960153, 4.958697, 4.957186, 4.956329, 4.956063, 4.956516, 4.957662, 
    4.959669, 4.961869, 4.964588, 4.965552, 4.966871, 4.968566, 4.970642, 
    4.973103, 4.975951, 4.979178, 4.982767, 4.986686, 4.990888, 4.995302, 
    4.99984, 5.004383, 5.008787, 5.012877, 5.016449, 5.019275, 5.021107, 
    5.021693,
  // momentumX(27,32, 0-49)
    4.992704, 4.991362, 4.989981, 4.988571, 4.987143, 4.985699, 4.984235, 
    4.982752, 4.981244, 4.979711, 4.978148, 4.976559, 4.974949, 4.97334, 
    4.971759, 4.970668, 4.96088, 4.960486, 4.96041, 4.960387, 4.96035, 
    4.958791, 4.957444, 4.956033, 4.955215, 4.954963, 4.95541, 4.956527, 
    4.958438, 4.960497, 4.962925, 4.964082, 4.965597, 4.967487, 4.969763, 
    4.972429, 4.975488, 4.97893, 4.982742, 4.986887, 4.991313, 4.995951, 
    5.000702, 5.005444, 5.010021, 5.014254, 5.017927, 5.020806, 5.022637, 
    5.023165,
  // momentumX(27,33, 0-49)
    4.993176, 4.991786, 4.990337, 4.988843, 4.987313, 4.98575, 4.984156, 
    4.982533, 4.980882, 4.979203, 4.977501, 4.975778, 4.97404, 4.972296, 
    4.97056, 4.969613, 4.960853, 4.960111, 4.959667, 4.95929, 4.95894, 
    4.957603, 4.956401, 4.955134, 4.954391, 4.954172, 4.954613, 4.955681, 
    4.957458, 4.959333, 4.961436, 4.962754, 4.964429, 4.966482, 4.968922, 
    4.971757, 4.974994, 4.978625, 4.982632, 4.986979, 4.991614, 4.996459, 
    5.001411, 5.006339, 5.011081, 5.015445, 5.019209, 5.022128, 5.023943, 
    5.024394,
  // momentumX(27,34, 0-49)
    4.993468, 4.992046, 4.990543, 4.988973, 4.98735, 4.985679, 4.983964, 
    4.982211, 4.980426, 4.978615, 4.976783, 4.974936, 4.973081, 4.971223, 
    4.96936, 4.968389, 4.960826, 4.959777, 4.958998, 4.958305, 4.957679, 
    4.956588, 4.955568, 4.954486, 4.953852, 4.953686, 4.95412, 4.955118, 
    4.956721, 4.958376, 4.960136, 4.961588, 4.963395, 4.965575, 4.968145, 
    4.971118, 4.974501, 4.978288, 4.98246, 4.986983, 4.9918, 4.996827, 
    5.001957, 5.00705, 5.011934, 5.016407, 5.020238, 5.023174, 5.024948, 
    5.025294,
  // momentumX(27,35, 0-49)
    4.993543, 4.992109, 4.990572, 4.988945, 4.987246, 4.98548, 4.983659, 
    4.98179, 4.979885, 4.977952, 4.976004, 4.97405, 4.972095, 4.970143, 
    4.968186, 4.967057, 4.960784, 4.959477, 4.958406, 4.957438, 4.956577, 
    4.955748, 4.954938, 4.954085, 4.953589, 4.953495, 4.953919, 4.954828, 
    4.956221, 4.957632, 4.959045, 4.960607, 4.962515, 4.964794, 4.967463, 
    4.970541, 4.974034, 4.977944, 4.982249, 4.986913, 4.991876, 4.997052, 
    5.002326, 5.007547, 5.012538, 5.017087, 5.020951, 5.023866, 5.025561, 
    5.025771,
  // momentumX(27,36, 0-49)
    4.993363, 4.991943, 4.990395, 4.988733, 4.986978, 4.985139, 4.983231, 
    4.981265, 4.979257, 4.977222, 4.975175, 4.973129, 4.971095, 4.969073, 
    4.967054, 4.965679, 4.960728, 4.959213, 4.957893, 4.956695, 4.95564, 
    4.955082, 4.954507, 4.953914, 4.953588, 4.953581, 4.953995, 4.954797, 
    4.955952, 4.957104, 4.958177, 4.959828, 4.961814, 4.964163, 4.966903, 
    4.970053, 4.973625, 4.977619, 4.982017, 4.986782, 4.991848, 4.997127, 
    5.002496, 5.007801, 5.012851, 5.017424, 5.021269, 5.024117, 5.025689, 
    5.025723,
  // momentumX(27,37, 0-49)
    4.992894, 4.991515, 4.989983, 4.988314, 4.986529, 4.984643, 4.982672, 
    4.980633, 4.978547, 4.97643, 4.974305, 4.972188, 4.970094, 4.968026, 
    4.965975, 4.964311, 4.960664, 4.958989, 4.957465, 4.956078, 4.95487, 
    4.954582, 4.954257, 4.953956, 4.953823, 4.953918, 4.954322, 4.955003, 
    4.955902, 4.956789, 4.957542, 4.959267, 4.961312, 4.963708, 4.96649, 
    4.969682, 4.973296, 4.977336, 4.981783, 4.986598, 4.991717, 4.997042, 
    5.00245, 5.007774, 5.01282, 5.017355, 5.021121, 5.02384, 5.025236, 
    5.025045,
  // momentumX(27,38, 0-49)
    4.992102, 4.990796, 4.989309, 4.987664, 4.985879, 4.983975, 4.981972, 
    4.979889, 4.977752, 4.97558, 4.973402, 4.971236, 4.969102, 4.967009, 
    4.964951, 4.962999, 4.960605, 4.958811, 4.957121, 4.955583, 4.954257, 
    4.954235, 4.954173, 4.954182, 4.954263, 4.954476, 4.954871, 4.955422, 
    4.956054, 4.956684, 4.957149, 4.958934, 4.961021, 4.963445, 4.966245, 
    4.969447, 4.97307, 4.977113, 4.981561, 4.986373, 4.991481, 4.996788, 
    5.002161, 5.007431, 5.012395, 5.016815, 5.020426, 5.022949, 5.024106, 
    5.023642,
  // momentumX(27,39, 0-49)
    4.990971, 4.989764, 4.988355, 4.986764, 4.985014, 4.983126, 4.981123, 
    4.97903, 4.976871, 4.974676, 4.97247, 4.970282, 4.968132, 4.966033, 
    4.963985, 4.961775, 4.960558, 4.95868, 4.956858, 4.955204, 4.953793, 
    4.954025, 4.954226, 4.954561, 4.954874, 4.955217, 4.955606, 4.956029, 
    4.956393, 4.956779, 4.956996, 4.958832, 4.960948, 4.963384, 4.966179, 
    4.969365, 4.972958, 4.976961, 4.981358, 4.986107, 4.991138, 4.99635, 
    5.001607, 5.006737, 5.011529, 5.015744, 5.019113, 5.021358, 5.022209, 
    5.021421,
  // momentumX(27,40, 0-49)
    4.989492, 4.988411, 4.987108, 4.985605, 4.983923, 4.982087, 4.980121, 
    4.978053, 4.975909, 4.973721, 4.971519, 4.969333, 4.96719, 4.965103, 
    4.963079, 4.960662, 4.960529, 4.958594, 4.956668, 4.954926, 4.953461, 
    4.953931, 4.954395, 4.955062, 4.955615, 4.956097, 4.956487, 4.956788, 
    4.956896, 4.957064, 4.957074, 4.958955, 4.961094, 4.963527, 4.966299, 
    4.96944, 4.972969, 4.976889, 4.98118, 4.9858, 4.990678, 4.995711, 
    5.000761, 5.005651, 5.010171, 5.01408, 5.017112, 5.018996, 5.019468, 
    5.018303,
  // momentumX(27,41, 0-49)
    4.98767, 4.986738, 4.98557, 4.984185, 4.982606, 4.98086, 4.978968, 
    4.97696, 4.974867, 4.972721, 4.970555, 4.9684, 4.966283, 4.964226, 
    4.962235, 4.959669, 4.96052, 4.958544, 4.956538, 4.954738, 4.95324, 
    4.953933, 4.95465, 4.955646, 4.956444, 4.957076, 4.957476, 4.957663, 
    4.957536, 4.957518, 4.957366, 4.959292, 4.961448, 4.963868, 4.9666, 
    4.969671, 4.973102, 4.976892, 4.98102, 4.985444, 4.99009, 4.994852, 
    4.999594, 5.004138, 5.008276, 5.01177, 5.014363, 5.015793, 5.015814, 
    5.014226,
  // momentumX(27,42, 0-49)
    4.985522, 4.98476, 4.983753, 4.982516, 4.981074, 4.97945, 4.977669, 
    4.975759, 4.973754, 4.971684, 4.969582, 4.967484, 4.965418, 4.963405, 
    4.961457, 4.958804, 4.960528, 4.958524, 4.956461, 4.954623, 4.953115, 
    4.954007, 4.954963, 4.956277, 4.957321, 4.958108, 4.958529, 4.958621, 
    4.958286, 4.958118, 4.957849, 4.959821, 4.961989, 4.96439, 4.967066, 
    4.970046, 4.973344, 4.976959, 4.980868, 4.985023, 4.989351, 4.993749, 
    4.998077, 5.002162, 5.005802, 5.008768, 5.010814, 5.011698, 5.011199, 
    5.009146,
  // momentumX(27,43, 0-49)
    4.983078, 4.982504, 4.981679, 4.980618, 4.979343, 4.977874, 4.976239, 
    4.974464, 4.972579, 4.970617, 4.968614, 4.966598, 4.964602, 4.962647, 
    4.96075, 4.958064, 4.960546, 4.958526, 4.956423, 4.954565, 4.953062, 
    4.954131, 4.955307, 4.956923, 4.958204, 4.959147, 4.959601, 4.959621, 
    4.959113, 4.958833, 4.958492, 4.960511, 4.962692, 4.965067, 4.967675, 
    4.97054, 4.973672, 4.977067, 4.980697, 4.984512, 4.988438, 4.992373, 
    4.996177, 4.999687, 5.00271, 5.00503, 5.006423, 5.006673, 5.005592, 
    5.003043,
  // momentumX(27,44, 0-49)
    4.980382, 4.980007, 4.979383, 4.978521, 4.97744, 4.976157, 4.974699, 
    4.973089, 4.971357, 4.969535, 4.967654, 4.965747, 4.963842, 4.961959, 
    4.960116, 4.957444, 4.96057, 4.958542, 4.956412, 4.954548, 4.953062, 
    4.954283, 4.955656, 4.957548, 4.959053, 4.960151, 4.960651, 4.960621, 
    4.959981, 4.95963, 4.959256, 4.961325, 4.963518, 4.965861, 4.968388, 
    4.971116, 4.974051, 4.97718, 4.980473, 4.983876, 4.987314, 4.990685, 
    4.993859, 4.996679, 4.998967, 5.000529, 5.001168, 5.000703, 4.998985, 
    4.995923,
  // momentumX(27,45, 0-49)
    4.977487, 4.977318, 4.976908, 4.976263, 4.975397, 4.974328, 4.973073, 
    4.971658, 4.970108, 4.968452, 4.96672, 4.964941, 4.963143, 4.961346, 
    4.959565, 4.956938, 4.960594, 4.958564, 4.956421, 4.954561, 4.953098, 
    4.954445, 4.955987, 4.958123, 4.959834, 4.961078, 4.961632, 4.961581, 
    4.960852, 4.960466, 4.960093, 4.962214, 4.964419, 4.966725, 4.969159, 
    4.971728, 4.974432, 4.977252, 4.980149, 4.983069, 4.985935, 4.988648, 
    4.991086, 4.993104, 4.994545, 4.995243, 4.995037, 4.993789, 4.991396, 
    4.987819,
  // momentumX(27,46, 0-49)
    4.974452, 4.974493, 4.974304, 4.97389, 4.973258, 4.972421, 4.971393, 
    4.970196, 4.968852, 4.967385, 4.965823, 4.964191, 4.962515, 4.960814, 
    4.959103, 4.956544, 4.960613, 4.958589, 4.956441, 4.954591, 4.953156, 
    4.954598, 4.956281, 4.95862, 4.960506, 4.961886, 4.962506, 4.96246, 
    4.961684, 4.961299, 4.960954, 4.963126, 4.965339, 4.9676, 4.969926, 
    4.972314, 4.974755, 4.97722, 4.979667, 4.982036, 4.98425, 4.986214, 
    4.987817, 4.988932, 4.989427, 4.989168, 4.988042, 4.98596, 4.982873, 
    4.9788,
  // momentumX(27,47, 0-49)
    4.971342, 4.971589, 4.971627, 4.971451, 4.971065, 4.970476, 4.969693, 
    4.968733, 4.967612, 4.966353, 4.964977, 4.963507, 4.961967, 4.960371, 
    4.958735, 4.956259, 4.960622, 4.95861, 4.956469, 4.954632, 4.953219, 
    4.954731, 4.956517, 4.959014, 4.961045, 4.962544, 4.963233, 4.963216, 
    4.962434, 4.962078, 4.961781, 4.963998, 4.966213, 4.96842, 4.970622, 
    4.972805, 4.974948, 4.977016, 4.978959, 4.98071, 4.982198, 4.983331, 
    4.98401, 4.984134, 4.9836, 4.982316, 4.980217, 4.977271, 4.973495, 
    4.968967,
  // momentumX(27,48, 0-49)
    4.968221, 4.96867, 4.968932, 4.968997, 4.968864, 4.968532, 4.968005, 
    4.967294, 4.966412, 4.965373, 4.964195, 4.962899, 4.961504, 4.960023, 
    4.958469, 4.956077, 4.960622, 4.958631, 4.9565, 4.954679, 4.953285, 
    4.954834, 4.956685, 4.959286, 4.961421, 4.963017, 4.963776, 4.963808, 
    4.963056, 4.96275, 4.962512, 4.964767, 4.96697, 4.969106, 4.971163, 
    4.973114, 4.974928, 4.976556, 4.977943, 4.97902, 4.979716, 4.979949, 
    4.979635, 4.978698, 4.977073, 4.974717, 4.971618, 4.96781, 4.963374, 
    4.958452,
  // momentumX(27,49, 0-49)
    4.964688, 4.965261, 4.965686, 4.965944, 4.966022, 4.965912, 4.965609, 
    4.96511, 4.964419, 4.963542, 4.962485, 4.96126, 4.959875, 4.958338, 
    4.95665, 4.953324, 4.963948, 4.960972, 4.957505, 4.954463, 4.952101, 
    4.95546, 4.959188, 4.964164, 4.967905, 4.970287, 4.97073, 4.969472, 
    4.966397, 4.964046, 4.961688, 4.964251, 4.966651, 4.968855, 4.970845, 
    4.972581, 4.974022, 4.975112, 4.975787, 4.975982, 4.975631, 4.974669, 
    4.973047, 4.97073, 4.967712, 4.964019, 4.959729, 4.954966, 4.949904, 
    4.944765,
  // momentumX(28,0, 0-49)
    4.963037, 4.965694, 4.96799, 4.96993, 4.971521, 4.972774, 4.973701, 
    4.974322, 4.97466, 4.974749, 4.974625, 4.974331, 4.973917, 4.973434, 
    4.972936, 4.972286, 4.972091, 4.971761, 4.971567, 4.971555, 4.971744, 
    4.972298, 4.973012, 4.97391, 4.974973, 4.97617, 4.977477, 4.978871, 
    4.980332, 4.981852, 4.983389, 4.985156, 4.986973, 4.988846, 4.990781, 
    4.992773, 4.99481, 4.99686, 4.998869, 5.000762, 5.002431, 5.003738, 
    5.00451, 5.00454, 5.003603, 5.00145, 4.997844, 4.992567, 4.985462, 
    4.976461,
  // momentumX(28,1, 0-49)
    4.964329, 4.966931, 4.969166, 4.971049, 4.972588, 4.973791, 4.974676, 
    4.975263, 4.975576, 4.975647, 4.975512, 4.975218, 4.974807, 4.97433, 
    4.973841, 4.973016, 4.97299, 4.972588, 4.972288, 4.972158, 4.972225, 
    4.97281, 4.973512, 4.974387, 4.975416, 4.976565, 4.977803, 4.979111, 
    4.980468, 4.981872, 4.983257, 4.985047, 4.986896, 4.988817, 4.990819, 
    4.992906, 4.995065, 4.997271, 4.999474, 5.001599, 5.003541, 5.005161, 
    5.006287, 5.006708, 5.006192, 5.004486, 5.001334, 4.996506, 4.989824, 
    4.981192,
  // momentumX(28,2, 0-49)
    4.965621, 4.968162, 4.970339, 4.972167, 4.973656, 4.974818, 4.975669, 
    4.976233, 4.976532, 4.976597, 4.976467, 4.976181, 4.975784, 4.975326, 
    4.974851, 4.973862, 4.973973, 4.973501, 4.973098, 4.972849, 4.972789, 
    4.973388, 4.974058, 4.974888, 4.97586, 4.976943, 4.978105, 4.979328, 
    4.98059, 4.981882, 4.983115, 4.984918, 4.986787, 4.988737, 4.990783, 
    4.992933, 4.995179, 4.997493, 4.999833, 5.002124, 5.004266, 5.00612, 
    5.007517, 5.00825, 5.008084, 5.006764, 5.004031, 4.999646, 4.993412, 
    4.985214,
  // momentumX(28,3, 0-49)
    4.966917, 4.969394, 4.971512, 4.973285, 4.974725, 4.975849, 4.976673, 
    4.977219, 4.97751, 4.977582, 4.977464, 4.977196, 4.976823, 4.976389, 
    4.975935, 4.974799, 4.974998, 4.974462, 4.973961, 4.973601, 4.973414, 
    4.97401, 4.974627, 4.975387, 4.976283, 4.977287, 4.978371, 4.979517, 
    4.980698, 4.981891, 4.98298, 4.984787, 4.986662, 4.988626, 4.990697, 
    4.992883, 4.995177, 4.997558, 4.999983, 5.002381, 5.004653, 5.00667, 
    5.008263, 5.009232, 5.009345, 5.008354, 5.006002, 5.002043, 4.996274, 
    4.988564,
  // momentumX(28,4, 0-49)
    4.968223, 4.970632, 4.972686, 4.974402, 4.975794, 4.97688, 4.977679, 
    4.97821, 4.978501, 4.97858, 4.978481, 4.97824, 4.977897, 4.977489, 
    4.97706, 4.975801, 4.976025, 4.975429, 4.974844, 4.97438, 4.974075, 
    4.974649, 4.975199, 4.975864, 4.976665, 4.977577, 4.978583, 4.979664, 
    4.980787, 4.981899, 4.982858, 4.984657, 4.986529, 4.988494, 4.99057, 
    4.992767, 4.99508, 4.997489, 4.999952, 5.002404, 5.004749, 5.006863, 
    5.008582, 5.00972, 5.010053, 5.009339, 5.007329, 5.00378, 4.998486, 
    4.991301,
  // momentumX(28,5, 0-49)
    4.969545, 4.971881, 4.973867, 4.975522, 4.976862, 4.977907, 4.978678, 
    4.979195, 4.979484, 4.979575, 4.979497, 4.979285, 4.978973, 4.978598, 
    4.978193, 4.976839, 4.977013, 4.976367, 4.975714, 4.975161, 4.97475, 
    4.975285, 4.975749, 4.976297, 4.976986, 4.977798, 4.978731, 4.979761, 
    4.980849, 4.981899, 4.982753, 4.984535, 4.986391, 4.988342, 4.990406, 
    4.992593, 4.994897, 4.997301, 4.999764, 5.002223, 5.00459, 5.006744, 
    5.008537, 5.009789, 5.010285, 5.009804, 5.008102, 5.004949, 5.000133, 
    4.993503,
  // momentumX(28,6, 0-49)
    4.970886, 4.97314, 4.975051, 4.976639, 4.977922, 4.978922, 4.979661, 
    4.98016, 4.980445, 4.980545, 4.980488, 4.980305, 4.980027, 4.979684, 
    4.979302, 4.977885, 4.977926, 4.977243, 4.97654, 4.975917, 4.975418, 
    4.975897, 4.97626, 4.976669, 4.977231, 4.977938, 4.978801, 4.979794, 
    4.980872, 4.981885, 4.982657, 4.984412, 4.986242, 4.988164, 4.990201, 
    4.992358, 4.994633, 4.997004, 4.999434, 5.001863, 5.00421, 5.006363, 
    5.008183, 5.0095, 5.010123, 5.009836, 5.008419, 5.005644, 5.001309, 
    4.995253,
  // momentumX(28,7, 0-49)
    4.97225, 4.974414, 4.976242, 4.977755, 4.978972, 4.979918, 4.980618, 
    4.981094, 4.98137, 4.981475, 4.981435, 4.981279, 4.981033, 4.980721, 
    4.98036, 4.978918, 4.978734, 4.978028, 4.977297, 4.976627, 4.976062, 
    4.976467, 4.976714, 4.976967, 4.977389, 4.977985, 4.978783, 4.979753, 
    4.980847, 4.981849, 4.982569, 4.984282, 4.986072, 4.987955, 4.989949, 
    4.992061, 4.994284, 4.996599, 4.998971, 5.001343, 5.003639, 5.005757, 
    5.007569, 5.008923, 5.00964, 5.009525, 5.00837, 5.005964, 5.002109, 
    4.996638,
  // momentumX(28,8, 0-49)
    4.973632, 4.975698, 4.977432, 4.978859, 4.980003, 4.980888, 4.981541, 
    4.981984, 4.982244, 4.982347, 4.98232, 4.982186, 4.981969, 4.981684, 
    4.98134, 4.979915, 4.979413, 4.978697, 4.977963, 4.977275, 4.97667, 
    4.976981, 4.977097, 4.97718, 4.977454, 4.977934, 4.978669, 4.97963, 
    4.980763, 4.981778, 4.982479, 4.984136, 4.985872, 4.987704, 4.989642, 
    4.991693, 4.99385, 4.996092, 4.998385, 5.00068, 5.002903, 5.004966, 
    5.006748, 5.008116, 5.00891, 5.00895, 5.008045, 5.005998, 5.00262, 
    4.997739,
  // momentumX(28,9, 0-49)
    4.975026, 4.976983, 4.978614, 4.979947, 4.981006, 4.98182, 4.982415, 
    4.982818, 4.983053, 4.983148, 4.983126, 4.983008, 4.982814, 4.982553, 
    4.982228, 4.980858, 4.979939, 4.979236, 4.978528, 4.977848, 4.977229, 
    4.97743, 4.977406, 4.977305, 4.977422, 4.977784, 4.978463, 4.979421, 
    4.980612, 4.981666, 4.98238, 4.983967, 4.985638, 4.987401, 4.989273, 
    4.991251, 4.993327, 4.995483, 4.997686, 4.999889, 5.002028, 5.004021, 
    5.005765, 5.007137, 5.007996, 5.008182, 5.00752, 5.005828, 5.002922, 
    4.998632,
  // momentumX(28,10, 0-49)
    4.976417, 4.978255, 4.979773, 4.981001, 4.981967, 4.9827, 4.98323, 
    4.983584, 4.983787, 4.983865, 4.98384, 4.983733, 4.983557, 4.983315, 
    4.983003, 4.981734, 4.980297, 4.979631, 4.978978, 4.97834, 4.977737, 
    4.977809, 4.977633, 4.977343, 4.9773, 4.977544, 4.978166, 4.979129, 
    4.980392, 4.981504, 4.982268, 4.983768, 4.985357, 4.987044, 4.988835, 
    4.990729, 4.992716, 4.994777, 4.996881, 4.998987, 5.001035, 5.002955, 
    5.004656, 5.00603, 5.006954, 5.007286, 5.006864, 5.005523, 5.003084, 
    4.999376,
  // momentumX(28,11, 0-49)
    4.977788, 4.979498, 4.980894, 4.982008, 4.982872, 4.983517, 4.983973, 
    4.984268, 4.984429, 4.984483, 4.984451, 4.984347, 4.984181, 4.983957, 
    4.983658, 4.98253, 4.980477, 4.979874, 4.979309, 4.978745, 4.978193, 
    4.978118, 4.977784, 4.977296, 4.977094, 4.977222, 4.97779, 4.978761, 
    4.980103, 4.981291, 4.982141, 4.983537, 4.985031, 4.986626, 4.988327, 
    4.990128, 4.992017, 4.993978, 4.995981, 4.997988, 4.999948, 5.001796, 
    5.00346, 5.004842, 5.005836, 5.006314, 5.006134, 5.005139, 5.003159, 
    5.000023,
  // momentumX(28,12, 0-49)
    4.979121, 4.98069, 4.981956, 4.982948, 4.983704, 4.984252, 4.984627, 
    4.984859, 4.984973, 4.984995, 4.984945, 4.984837, 4.984681, 4.984471, 
    4.984189, 4.983234, 4.980469, 4.979962, 4.979518, 4.979064, 4.978595, 
    4.978358, 4.977861, 4.977178, 4.976821, 4.976835, 4.97735, 4.978325, 
    4.979751, 4.981029, 4.981995, 4.983273, 4.984656, 4.986147, 4.987747, 
    4.989446, 4.991234, 4.993092, 4.994994, 4.996906, 4.998783, 5.000571, 
    5.002206, 5.003607, 5.004677, 5.00531, 5.005374, 5.004723, 5.003193, 
    5.000611,
  // momentumX(28,13, 0-49)
    4.980392, 4.981812, 4.982938, 4.983803, 4.984443, 4.98489, 4.985179, 
    4.985341, 4.985403, 4.985387, 4.985314, 4.985199, 4.985044, 4.984848, 
    4.984589, 4.983837, 4.980271, 4.979891, 4.979608, 4.979298, 4.978949, 
    4.978534, 4.977874, 4.977001, 4.976495, 4.976401, 4.976861, 4.977839, 
    4.979345, 4.980719, 4.981833, 4.982975, 4.984235, 4.98561, 4.987098, 
    4.988689, 4.990372, 4.992128, 4.993932, 4.995756, 4.997561, 4.999301, 
    5.00092, 5.002353, 5.003514, 5.00431, 5.004621, 5.004309, 5.003215, 
    5.001168,
  // momentumX(28,14, 0-49)
    4.981575, 4.982839, 4.983819, 4.984552, 4.985072, 4.985415, 4.985616, 
    4.985703, 4.985707, 4.98565, 4.98555, 4.985421, 4.985268, 4.985085, 
    4.984856, 4.98433, 4.97988, 4.979667, 4.979576, 4.979448, 4.979251, 
    4.97865, 4.977829, 4.976778, 4.976137, 4.975942, 4.976348, 4.97732, 
    4.978895, 4.98037, 4.981659, 4.982649, 4.98377, 4.985018, 4.986386, 
    4.987864, 4.989438, 4.991094, 4.992805, 4.99455, 4.996294, 4.998002, 
    4.999622, 5.001102, 5.002368, 5.003336, 5.003896, 5.003918, 5.003249, 
    5.001713,
  // momentumX(28,15, 0-49)
    4.982654, 4.983751, 4.984578, 4.985173, 4.985571, 4.985808, 4.985918, 
    4.98593, 4.985873, 4.985772, 4.985643, 4.985499, 4.985344, 4.985178, 
    4.984991, 4.984704, 4.979304, 4.979292, 4.979429, 4.979517, 4.979506, 
    4.978709, 4.977736, 4.976521, 4.975759, 4.975474, 4.975827, 4.976785, 
    4.978418, 4.979989, 4.981472, 4.982297, 4.983266, 4.984376, 4.985615, 
    4.986974, 4.988441, 4.989997, 4.991624, 4.993299, 4.994998, 4.996687, 
    4.998328, 4.999872, 5.001257, 5.002406, 5.003217, 5.003567, 5.003305, 
    5.002254,
  // momentumX(28,16, 0-49)
    4.983608, 4.984528, 4.985196, 4.98565, 4.985922, 4.986052, 4.98607, 
    4.986007, 4.98589, 4.985743, 4.985583, 4.985423, 4.985268, 4.985124, 
    4.984986, 4.984951, 4.978553, 4.978775, 4.979172, 4.979506, 4.979712, 
    4.978718, 4.977604, 4.976244, 4.975379, 4.975018, 4.975318, 4.976254, 
    4.977931, 4.979589, 4.981279, 4.981926, 4.98273, 4.983689, 4.984793, 
    4.986029, 4.987384, 4.988845, 4.990394, 4.992012, 4.993679, 4.995368, 
    4.997046, 4.998671, 5.000189, 5.001527, 5.002593, 5.003264, 5.003393, 
    5.002801,
  // momentumX(28,17, 0-49)
    4.984422, 4.985153, 4.985654, 4.985961, 4.986106, 4.986128, 4.986056, 
    4.985919, 4.985743, 4.985553, 4.985363, 4.985186, 4.985034, 4.984914, 
    4.984838, 4.985061, 4.977653, 4.978134, 4.978813, 4.97942, 4.979869, 
    4.978677, 4.977434, 4.975953, 4.975008, 4.974584, 4.974835, 4.975744, 
    4.977448, 4.979182, 4.981081, 4.981539, 4.982168, 4.982968, 4.983927, 
    4.985033, 4.986276, 4.987643, 4.98912, 4.990694, 4.992342, 4.994048, 
    4.995781, 4.997505, 4.999168, 5.000705, 5.002026, 5.00301, 5.003512, 
    5.003355,
  // momentumX(28,18, 0-49)
    4.985089, 4.985617, 4.985938, 4.98609, 4.986105, 4.986018, 4.985858, 
    4.985652, 4.985424, 4.985193, 4.984977, 4.984787, 4.98464, 4.984551, 
    4.984545, 4.985033, 4.976648, 4.977406, 4.978383, 4.979276, 4.979985, 
    4.978594, 4.977239, 4.975657, 4.97465, 4.974179, 4.974391, 4.975267, 
    4.976982, 4.978776, 4.980881, 4.981141, 4.981584, 4.982214, 4.98302, 
    4.983992, 4.985119, 4.986394, 4.987806, 4.989342, 4.990986, 4.992723, 
    4.994529, 4.996365, 4.998188, 4.999933, 5.00151, 5.002803, 5.003664, 
    5.003913,
  // momentumX(28,19, 0-49)
    4.985601, 4.985903, 4.986029, 4.986017, 4.985898, 4.985704, 4.985462, 
    4.985194, 4.98492, 4.984657, 4.984419, 4.984222, 4.984084, 4.984033, 
    4.984104, 4.984866, 4.975602, 4.976647, 4.977926, 4.979109, 4.980078, 
    4.978496, 4.977036, 4.975368, 4.974319, 4.973816, 4.973994, 4.974836, 
    4.976551, 4.978387, 4.980682, 4.980737, 4.980986, 4.981435, 4.982077, 
    4.982903, 4.983911, 4.985092, 4.986441, 4.987948, 4.989601, 4.991385, 
    4.993277, 4.995243, 4.997238, 4.999198, 5.001037, 5.002635, 5.003841, 
    5.004478,
  // momentumX(28,20, 0-49)
    4.986712, 4.987498, 4.98811, 4.988571, 4.988906, 4.989136, 4.989282, 
    4.98936, 4.98939, 4.989389, 4.989371, 4.989356, 4.989365, 4.989432, 
    4.989607, 0, 4.973971, 4.974906, 4.976127, 4.977295, 4.978267, 4.976232, 
    4.974376, 4.972327, 4.970971, 4.970251, 4.970322, 4.971179, 4.973058, 
    4.975195, 4.977999, 4.978202, 4.978607, 4.979215, 4.980005, 4.980972, 
    4.982105, 4.983404, 4.984862, 4.986478, 4.988243, 4.990149, 4.992177, 
    4.994302, 4.996484, 4.998657, 5.000737, 5.002606, 5.004115, 5.005083,
  // momentumX(28,21, 0-49)
    4.987054, 4.987665, 4.988129, 4.988471, 4.988711, 4.988868, 4.988958, 
    4.989, 4.989004, 4.988986, 4.988958, 4.988937, 4.988944, 4.989013, 
    4.989195, 0, 4.970282, 4.971366, 4.97281, 4.974231, 4.975453, 4.973234, 
    4.971309, 4.969253, 4.967992, 4.967446, 4.967751, 4.968876, 4.971061, 
    4.973518, 4.976734, 4.976965, 4.977419, 4.978096, 4.978973, 4.980039, 
    4.981282, 4.982694, 4.984271, 4.986003, 4.987885, 4.989907, 4.992052, 
    4.994292, 4.996589, 4.998882, 5.001087, 5.003087, 5.004737, 5.00586,
  // momentumX(28,22, 0-49)
    4.987328, 4.98778, 4.988113, 4.988348, 4.988502, 4.988594, 4.988635, 
    4.98864, 4.988618, 4.988581, 4.988539, 4.988505, 4.988502, 4.988559, 
    4.988728, 0, 4.967324, 4.968526, 4.970151, 4.971785, 4.973213, 4.970802, 
    4.968777, 4.96666, 4.965425, 4.964967, 4.965406, 4.966697, 4.969078, 
    4.97174, 4.975243, 4.975431, 4.975869, 4.976557, 4.977474, 4.978605, 
    4.979939, 4.981463, 4.98317, 4.985048, 4.987089, 4.989276, 4.991593, 
    4.994008, 4.996481, 4.99895, 5.001328, 5.003502, 5.005326, 5.006629,
  // momentumX(28,23, 0-49)
    4.987549, 4.987857, 4.98807, 4.988206, 4.988283, 4.988314, 4.98831, 
    4.988281, 4.988234, 4.988175, 4.988117, 4.988068, 4.988048, 4.988085, 
    4.988226, 0, 4.964871, 4.966145, 4.967893, 4.969668, 4.971232, 4.968641, 
    4.966502, 4.964304, 4.963049, 4.962618, 4.963121, 4.964503, 4.966997, 
    4.96978, 4.973461, 4.973578, 4.97397, 4.974645, 4.975582, 4.976766, 
    4.978186, 4.979832, 4.981688, 4.983741, 4.985978, 4.988378, 4.990917, 
    4.993559, 4.996259, 4.998947, 5.001537, 5.003915, 5.005933, 5.007423,
  // momentumX(28,24, 0-49)
    4.98774, 4.98791, 4.988009, 4.988055, 4.98806, 4.988034, 4.987987, 
    4.987925, 4.987851, 4.987772, 4.987696, 4.987629, 4.987588, 4.987599, 
    4.987702, 0, 4.963188, 4.964485, 4.966293, 4.968147, 4.969785, 4.967083, 
    4.964877, 4.962627, 4.961349, 4.960917, 4.961437, 4.962847, 4.965379, 
    4.968204, 4.971961, 4.972018, 4.972366, 4.973018, 4.973957, 4.975173, 
    4.976654, 4.97839, 4.980366, 4.982566, 4.984974, 4.987565, 4.990309, 
    4.993167, 4.996087, 4.998994, 5.001799, 5.004381, 5.006594, 5.00827,
  // momentumX(28,25, 0-49)
    4.987918, 4.987956, 4.987947, 4.987906, 4.98784, 4.98776, 4.987669, 
    4.987572, 4.98747, 4.98737, 4.987273, 4.987188, 4.987124, 4.987105, 
    4.987164, 0, 4.961998, 4.963271, 4.96508, 4.966942, 4.96859, 4.965873, 
    4.963664, 4.961417, 4.960142, 4.95971, 4.960229, 4.96163, 4.964145, 
    4.966951, 4.9707, 4.97073, 4.971062, 4.971709, 4.972658, 4.973903, 
    4.975436, 4.977246, 4.979321, 4.981645, 4.984196, 4.986951, 4.989874, 
    4.992926, 4.996044, 4.999156, 5.002161, 5.00494, 5.007341, 5.009192,
  // momentumX(28,26, 0-49)
    4.988102, 4.988014, 4.9879, 4.98777, 4.987633, 4.987494, 4.987355, 
    4.987218, 4.987085, 4.986959, 4.98684, 4.986735, 4.98665, 4.986601, 
    4.986614, 0, 4.96127, 4.962483, 4.964233, 4.96604, 4.967638, 4.965005, 
    4.962867, 4.960688, 4.95945, 4.959028, 4.95953, 4.960891, 4.963342, 
    4.966077, 4.969729, 4.969779, 4.970129, 4.970798, 4.971775, 4.973054, 
    4.974634, 4.976504, 4.978654, 4.98107, 4.983733, 4.986615, 4.989684, 
    4.992893, 4.996181, 4.99947, 5.002655, 5.005613, 5.008188, 5.010205,
  // momentumX(28,27, 0-49)
    4.988311, 4.988101, 4.987882, 4.987662, 4.987448, 4.987243, 4.987047, 
    4.986861, 4.986687, 4.986527, 4.986381, 4.986256, 4.986153, 4.986082, 
    4.986058, 0, 4.961052, 4.962173, 4.963817, 4.96551, 4.967003, 4.964544, 
    4.962538, 4.960472, 4.959287, 4.958868, 4.959324, 4.960605, 4.962934, 
    4.965534, 4.969001, 4.969101, 4.969494, 4.970201, 4.971213, 4.972528, 
    4.974146, 4.97606, 4.978265, 4.980749, 4.983495, 4.986478, 4.989666, 
    4.993008, 4.996446, 4.999894, 5.003249, 5.006377, 5.009121, 5.011301,
  // momentumX(28,28, 0-49)
    4.988558, 4.98823, 4.987906, 4.987594, 4.987296, 4.987011, 4.986745, 
    4.986495, 4.986266, 4.986061, 4.985881, 4.985734, 4.98562, 4.985543, 
    4.985505, 0, 4.961629, 4.962648, 4.964153, 4.965688, 4.967029, 4.964806, 
    4.962961, 4.961018, 4.959865, 4.959403, 4.959753, 4.960879, 4.963003, 
    4.965382, 4.968564, 4.968718, 4.969153, 4.969889, 4.97092, 4.97225, 
    4.973881, 4.975813, 4.978045, 4.980568, 4.983372, 4.986431, 4.989717, 
    4.993181, 4.996759, 5.000366, 5.003891, 5.007196, 5.010116, 5.012463,
  // momentumX(28,29, 0-49)
    4.988853, 4.988415, 4.987991, 4.98758, 4.987185, 4.986807, 4.986447, 
    4.986111, 4.985805, 4.985536, 4.985315, 4.985149, 4.985041, 4.984988, 
    4.984979, 0, 4.96272, 4.963651, 4.965005, 4.966348, 4.967486, 4.965503, 
    4.96379, 4.961924, 4.960732, 4.960146, 4.960302, 4.961183, 4.963007, 
    4.965075, 4.967861, 4.968034, 4.96848, 4.969221, 4.970254, 4.97159, 
    4.973233, 4.975191, 4.977465, 4.980054, 4.982945, 4.986122, 4.989549, 
    4.993178, 4.996941, 5.000747, 5.004481, 5.007996, 5.01112, 5.013654,
  // momentumX(28,30, 0-49)
    4.98853, 4.987349, 4.986206, 4.985108, 4.984058, 4.983053, 4.98209, 
    4.981159, 4.980254, 4.979371, 4.978508, 4.977676, 4.976903, 4.976246, 
    4.975795, 4.974938, 4.965952, 4.966966, 4.968203, 4.969349, 4.970299, 
    4.968656, 4.967254, 4.965686, 4.964678, 4.964137, 4.964175, 4.964772, 
    4.966136, 4.967617, 4.969641, 4.969453, 4.969526, 4.969896, 4.970581, 
    4.971605, 4.972989, 4.974744, 4.976882, 4.979402, 4.982292, 4.98553, 
    4.989075, 4.992872, 4.996842, 5.000887, 5.004877, 5.008653, 5.012033, 
    5.014809,
  // momentumX(28,31, 0-49)
    4.988934, 4.987695, 4.986489, 4.98532, 4.98419, 4.983098, 4.982041, 
    4.981017, 4.980021, 4.979056, 4.978122, 4.977229, 4.976397, 4.975665, 
    4.975098, 4.974432, 4.965597, 4.966311, 4.967228, 4.96806, 4.968717, 
    4.96726, 4.965956, 4.96447, 4.963483, 4.962937, 4.96296, 4.963528, 
    4.964809, 4.96617, 4.967934, 4.96792, 4.968172, 4.968722, 4.969593, 
    4.970803, 4.972375, 4.97432, 4.976649, 4.979359, 4.982438, 4.985861, 
    4.989586, 4.993555, 4.997685, 5.001874, 5.005987, 5.009863, 5.013318, 
    5.016133,
  // momentumX(28,32, 0-49)
    4.989329, 4.988023, 4.986743, 4.985494, 4.984277, 4.983092, 4.98194, 
    4.980819, 4.979729, 4.978675, 4.977658, 4.976685, 4.97577, 4.974939, 
    4.974227, 4.97373, 4.965408, 4.965789, 4.966353, 4.966842, 4.96719, 
    4.965924, 4.964731, 4.963346, 4.9624, 4.961866, 4.961875, 4.962408, 
    4.963588, 4.964805, 4.966289, 4.966444, 4.96687, 4.967595, 4.96864, 
    4.970027, 4.971777, 4.973903, 4.976413, 4.979305, 4.982565, 4.986166, 
    4.990065, 4.994201, 4.998487, 5.002816, 5.007049, 5.011023, 5.014543, 
    5.017394,
  // momentumX(28,33, 0-49)
    4.989703, 4.988327, 4.986968, 4.985633, 4.984324, 4.983045, 4.981792, 
    4.980573, 4.979386, 4.978236, 4.977127, 4.976064, 4.975055, 4.974112, 
    4.973249, 4.97283, 4.965299, 4.96534, 4.965545, 4.96569, 4.965733, 
    4.964666, 4.963603, 4.962349, 4.961465, 4.960958, 4.96096, 4.961446, 
    4.962501, 4.963549, 4.96474, 4.96506, 4.965649, 4.966537, 4.967746, 
    4.969299, 4.971216, 4.973511, 4.976191, 4.979255, 4.982684, 4.986455, 
    4.990518, 4.994809, 4.99924, 5.003698, 5.008042, 5.0121, 5.015676, 
    5.018547,
  // momentumX(28,34, 0-49)
    4.990031, 4.988589, 4.987155, 4.985735, 4.984336, 4.982958, 4.981607, 
    4.980285, 4.978996, 4.977746, 4.976541, 4.975382, 4.974274, 4.973217, 
    4.972211, 4.971758, 4.965207, 4.964923, 4.964778, 4.964593, 4.964345, 
    4.963485, 4.962573, 4.961481, 4.960687, 4.960222, 4.960217, 4.960645, 
    4.961547, 4.962411, 4.963303, 4.963782, 4.964528, 4.965569, 4.966932, 
    4.96864, 4.970713, 4.973166, 4.976003, 4.979225, 4.982812, 4.986735, 
    4.990946, 4.995378, 4.999937, 5.004506, 5.008938, 5.013061, 5.01667, 
    5.019539,
  // momentumX(28,35, 0-49)
    4.990283, 4.988789, 4.987288, 4.985792, 4.984304, 4.982832, 4.981381, 
    4.979957, 4.978567, 4.977216, 4.97591, 4.974653, 4.973446, 4.97228, 
    4.971144, 4.970554, 4.965104, 4.964519, 4.964046, 4.963553, 4.96304, 
    4.962392, 4.96165, 4.960749, 4.960071, 4.959666, 4.959654, 4.960008, 
    4.960733, 4.961397, 4.961999, 4.96263, 4.963524, 4.964712, 4.966218, 
    4.96807, 4.970286, 4.972882, 4.975864, 4.979228, 4.982954, 4.987012, 
    4.991352, 4.995899, 5.000561, 5.005215, 5.009709, 5.013865, 5.017476, 
    5.020309,
  // momentumX(28,36, 0-49)
    4.990426, 4.988896, 4.987345, 4.985782, 4.984218, 4.982658, 4.981112, 
    4.97959, 4.9781, 4.976649, 4.975245, 4.973891, 4.972588, 4.971323, 
    4.970076, 4.969267, 4.964972, 4.964121, 4.963349, 4.962579, 4.961828, 
    4.961393, 4.960837, 4.960156, 4.959619, 4.959288, 4.959268, 4.959536, 
    4.960064, 4.96052, 4.960848, 4.961624, 4.962659, 4.963984, 4.965623, 
    4.967606, 4.969953, 4.972678, 4.975785, 4.979272, 4.983116, 4.987284, 
    4.991723, 4.996358, 5.001091, 5.005792, 5.010311, 5.014461, 5.01803, 
    5.020787,
  // momentumX(28,37, 0-49)
    4.99042, 4.988878, 4.987295, 4.985683, 4.984055, 4.98242, 4.980792, 
    4.97918, 4.977595, 4.97605, 4.974551, 4.973106, 4.971712, 4.970358, 
    4.969019, 4.967945, 4.964811, 4.963729, 4.962691, 4.961675, 4.960719, 
    4.960494, 4.960138, 4.959701, 4.959327, 4.959084, 4.959058, 4.959228, 
    4.959541, 4.959791, 4.959871, 4.960784, 4.961951, 4.963401, 4.965164, 
    4.967265, 4.969728, 4.972565, 4.975777, 4.979362, 4.983298, 4.987546, 
    4.992053, 4.996737, 5.001498, 5.006205, 5.0107, 5.014793, 5.018272, 5.0209,
  // momentumX(28,38, 0-49)
    4.99023, 4.988701, 4.987109, 4.98547, 4.983797, 4.982105, 4.980407, 
    4.978717, 4.977051, 4.97542, 4.973835, 4.972305, 4.97083, 4.969398, 
    4.967984, 4.966624, 4.964621, 4.963344, 4.962071, 4.960845, 4.959713, 
    4.959695, 4.959548, 4.959376, 4.959183, 4.959043, 4.959011, 4.959078, 
    4.959167, 4.959216, 4.959079, 4.960124, 4.961415, 4.962979, 4.964853, 
    4.967059, 4.969621, 4.972549, 4.975846, 4.979504, 4.983499, 4.98779, 
    4.992322, 4.997014, 5.001755, 5.006413, 5.010828, 5.014806, 5.018132, 
    5.020571,
  // momentumX(28,39, 0-49)
    4.98982, 4.988333, 4.986758, 4.985115, 4.983422, 4.981692, 4.979945, 
    4.978195, 4.976461, 4.974759, 4.973101, 4.971496, 4.969948, 4.968448, 
    4.966973, 4.965341, 4.964407, 4.962965, 4.961492, 4.960084, 4.958814, 
    4.958994, 4.959059, 4.959167, 4.959174, 4.959148, 4.959116, 4.959077, 
    4.958942, 4.958804, 4.958484, 4.959653, 4.96106, 4.962731, 4.964701, 
    4.966998, 4.96964, 4.972637, 4.975991, 4.979691, 4.983709, 4.988005, 
    4.992517, 4.997162, 5.001826, 5.006374, 5.010642, 5.014437, 5.017542, 
    5.019726,
  // momentumX(28,40, 0-49)
    4.989163, 4.987743, 4.986215, 4.984596, 4.982908, 4.981167, 4.979392, 
    4.977604, 4.975822, 4.974064, 4.972347, 4.970681, 4.969072, 4.967516, 
    4.965992, 4.964116, 4.964172, 4.962595, 4.960951, 4.959398, 4.958017, 
    4.958385, 4.958663, 4.959061, 4.959281, 4.959382, 4.959355, 4.959212, 
    4.958863, 4.958557, 4.95809, 4.959379, 4.960891, 4.962658, 4.964714, 
    4.967083, 4.969785, 4.972829, 4.97621, 4.979917, 4.983921, 4.988175, 
    4.992615, 4.997153, 5.001677, 5.006044, 5.010092, 5.013627, 5.016435, 
    5.018291,
  // momentumX(28,41, 0-49)
    4.988236, 4.986912, 4.985459, 4.983894, 4.982239, 4.980513, 4.978737, 
    4.976935, 4.975128, 4.973335, 4.971576, 4.969865, 4.968209, 4.966607, 
    4.965042, 4.962963, 4.963916, 4.962226, 4.960443, 4.958775, 4.957313, 
    4.957856, 4.958346, 4.959037, 4.959479, 4.959718, 4.959705, 4.959471, 
    4.958921, 4.958473, 4.957899, 4.959299, 4.96091, 4.962762, 4.96489, 
    4.967316, 4.970056, 4.973118, 4.976497, 4.980174, 4.984117, 4.988278, 
    4.992589, 4.996957, 5.001267, 5.005378, 5.009124, 5.012317, 5.014746, 
    5.016197,
  // momentumX(28,42, 0-49)
    4.98703, 4.98583, 4.984478, 4.982997, 4.981404, 4.979722, 4.977974, 
    4.976183, 4.974374, 4.97257, 4.97079, 4.96905, 4.96736, 4.965723, 
    4.964126, 4.961891, 4.963639, 4.961859, 4.95996, 4.958206, 4.956691, 
    4.957398, 4.958096, 4.959077, 4.959745, 4.96013, 4.960144, 4.959831, 
    4.959105, 4.958547, 4.957901, 4.959409, 4.961112, 4.963038, 4.965222, 
    4.967688, 4.970444, 4.973498, 4.976838, 4.980443, 4.98428, 4.988293, 
    4.992411, 4.996538, 5.000558, 5.00433, 5.007689, 5.010449, 5.012415, 
    5.013385,
  // momentumX(28,43, 0-49)
    4.98554, 4.984489, 4.983268, 4.981898, 4.980398, 4.978789, 4.977099, 
    4.975349, 4.973565, 4.971771, 4.96999, 4.96824, 4.96653, 4.964868, 
    4.963245, 4.9609, 4.963339, 4.961486, 4.959499, 4.957683, 4.956139, 
    4.956997, 4.957892, 4.959154, 4.960049, 4.960588, 4.96064, 4.960272, 
    4.959402, 4.958764, 4.958083, 4.959694, 4.961483, 4.963474, 4.965702, 
    4.968185, 4.970934, 4.973947, 4.977213, 4.980706, 4.984384, 4.988188, 
    4.992046, 4.99586, 4.999508, 5.002852, 5.005733, 5.007973, 5.009391, 
    5.009803,
  // momentumX(28,44, 0-49)
    4.983782, 4.982901, 4.981836, 4.980603, 4.979224, 4.977719, 4.976113, 
    4.974431, 4.972697, 4.970939, 4.969179, 4.967435, 4.965723, 4.964047, 
    4.962406, 4.959991, 4.963014, 4.961103, 4.959048, 4.957194, 4.955643, 
    4.956639, 4.95772, 4.959247, 4.960364, 4.961061, 4.961168, 4.960768, 
    4.95979, 4.959107, 4.958425, 4.960135, 4.962002, 4.964049, 4.966306, 
    4.968788, 4.971504, 4.974445, 4.977598, 4.980931, 4.984395, 4.987931, 
    4.991458, 4.994877, 4.99807, 5.000897, 5.003209, 5.00484, 5.005627, 
    5.005414,
  // momentumX(28,45, 0-49)
    4.981774, 4.981083, 4.980196, 4.979126, 4.977894, 4.97652, 4.975028, 
    4.973438, 4.971782, 4.970082, 4.968363, 4.966645, 4.964943, 4.963265, 
    4.961613, 4.959162, 4.962658, 4.960703, 4.958603, 4.956729, 4.955187, 
    4.956307, 4.957557, 4.959331, 4.960659, 4.961514, 4.961693, 4.961289, 
    4.960246, 4.959553, 4.958898, 4.960707, 4.962646, 4.964738, 4.967009, 
    4.969471, 4.972126, 4.974962, 4.977961, 4.981081, 4.984278, 4.987478, 
    4.990602, 4.993547, 4.996198, 4.998419, 5.000072, 5.001008, 5.001089, 
    5.000189,
  // momentumX(28,46, 0-49)
    4.979548, 4.979063, 4.978371, 4.977488, 4.976427, 4.975208, 4.973854, 
    4.972385, 4.970828, 4.969208, 4.96755, 4.965873, 4.964198, 4.96253, 
    4.960874, 4.958412, 4.962271, 4.960286, 4.958158, 4.95628, 4.95476, 
    4.955986, 4.957387, 4.959378, 4.960902, 4.961915, 4.96218, 4.961805, 
    4.96074, 4.960072, 4.959472, 4.961374, 4.96338, 4.965507, 4.967777, 
    4.970197, 4.972763, 4.975461, 4.978261, 4.981122, 4.983987, 4.986786, 
    4.989431, 4.991823, 4.993845, 4.995374, 4.996282, 4.996446, 4.995755, 
    4.994122,
  // momentumX(28,47, 0-49)
    4.977147, 4.976876, 4.976397, 4.975716, 4.974848, 4.973806, 4.972611, 
    4.971286, 4.96985, 4.968332, 4.966752, 4.965134, 4.963496, 4.961848, 
    4.960196, 4.957739, 4.96185, 4.959847, 4.957707, 4.955839, 4.95435, 
    4.955663, 4.957192, 4.959366, 4.961065, 4.962229, 4.962596, 4.962281, 
    4.96124, 4.96063, 4.960107, 4.962099, 4.964166, 4.966316, 4.96857, 
    4.970924, 4.973373, 4.975894, 4.978453, 4.981, 4.983474, 4.985802, 
    4.987894, 4.98965, 4.990963, 4.991716, 4.991806, 4.991132, 4.989618, 
    4.987222,
  // momentumX(28,48, 0-49)
    4.974618, 4.974567, 4.974308, 4.973845, 4.973186, 4.972341, 4.971326, 
    4.970162, 4.968867, 4.967466, 4.965981, 4.964435, 4.962846, 4.961228, 
    4.959587, 4.957145, 4.961398, 4.959391, 4.957252, 4.9554, 4.953947, 
    4.955328, 4.956959, 4.959277, 4.961123, 4.962427, 4.962908, 4.962682, 
    4.96171, 4.961189, 4.960761, 4.962839, 4.964956, 4.967119, 4.969338, 
    4.971605, 4.973905, 4.976213, 4.978484, 4.980662, 4.982685, 4.984473, 
    4.98594, 4.986984, 4.987511, 4.987416, 4.986622, 4.985056, 4.982687, 
    4.979521,
  // momentumX(28,49, 0-49)
    4.971751, 4.97187, 4.971794, 4.971513, 4.971032, 4.970352, 4.969482, 
    4.968434, 4.96722, 4.965861, 4.964369, 4.962768, 4.961073, 4.959293, 
    4.957433, 4.953966, 4.963982, 4.960976, 4.957507, 4.954463, 4.952083, 
    4.955269, 4.95878, 4.963472, 4.966963, 4.969119, 4.969381, 4.967987, 
    4.964842, 4.962405, 4.959975, 4.962437, 4.964849, 4.967206, 4.969516, 
    4.971771, 4.973949, 4.976017, 4.977924, 4.979613, 4.981015, 4.982051, 
    4.98264, 4.982693, 4.982131, 4.980882, 4.978908, 4.976194, 4.972773, 
    4.968725,
  // momentumX(29,0, 0-49)
    4.971556, 4.973361, 4.974815, 4.975937, 4.976742, 4.97725, 4.977488, 
    4.977488, 4.977288, 4.976929, 4.976456, 4.97591, 4.975338, 4.97478, 
    4.974274, 4.973676, 4.973505, 4.973238, 4.973083, 4.97306, 4.973165, 
    4.973533, 4.973971, 4.974497, 4.975105, 4.975779, 4.976512, 4.977307, 
    4.978165, 4.979098, 4.980094, 4.981372, 4.982794, 4.984384, 4.986169, 
    4.988163, 4.99037, 4.992781, 4.995366, 4.998078, 5.000845, 5.003565, 
    5.00611, 5.008316, 5.009995, 5.010931, 5.010883, 5.009605, 5.006854, 
    5.002412,
  // momentumX(29,1, 0-49)
    4.97285, 4.9746, 4.976003, 4.977079, 4.977844, 4.97832, 4.978535, 
    4.978521, 4.978314, 4.977955, 4.977486, 4.976948, 4.976385, 4.975832, 
    4.975327, 4.974553, 4.974493, 4.974136, 4.97386, 4.973703, 4.973669, 
    4.97404, 4.974442, 4.974925, 4.975485, 4.976109, 4.976785, 4.977513, 
    4.978296, 4.979141, 4.980009, 4.981315, 4.982766, 4.984389, 4.986212, 
    4.988253, 4.990514, 4.992992, 4.995659, 4.998469, 5.001352, 5.00421, 
    5.006918, 5.009318, 5.011222, 5.012416, 5.012663, 5.011715, 5.009322, 
    5.005255,
  // momentumX(29,2, 0-49)
    4.974152, 4.975846, 4.977199, 4.978231, 4.97896, 4.979407, 4.979604, 
    4.979578, 4.979369, 4.979012, 4.978549, 4.978021, 4.977464, 4.976915, 
    4.976405, 4.97546, 4.975474, 4.975027, 4.974627, 4.974336, 4.974163, 
    4.974525, 4.97488, 4.975307, 4.975816, 4.976388, 4.977014, 4.977693, 
    4.978423, 4.979195, 4.979949, 4.981287, 4.982766, 4.984417, 4.986269, 
    4.988337, 4.990631, 4.993144, 4.995852, 4.998711, 5.001653, 5.004588, 
    5.007389, 5.009909, 5.011964, 5.013349, 5.013828, 5.013155, 5.011086, 
    5.007389,
  // momentumX(29,3, 0-49)
    4.975455, 4.977093, 4.978398, 4.979385, 4.98008, 4.980501, 4.980679, 
    4.980646, 4.980434, 4.980083, 4.979627, 4.979106, 4.978555, 4.978006, 
    4.977489, 4.976379, 4.976416, 4.975876, 4.975358, 4.974937, 4.97463, 
    4.974973, 4.975272, 4.975631, 4.976077, 4.976596, 4.977183, 4.977833, 
    4.978536, 4.979261, 4.979921, 4.981289, 4.982796, 4.98447, 4.98634, 
    4.988424, 4.990729, 4.993248, 4.995963, 4.998829, 5.001781, 5.004733, 
    5.007569, 5.010144, 5.012286, 5.013795, 5.014449, 5.014008, 5.01223, 
    5.008885,
  // momentumX(29,4, 0-49)
    4.976765, 4.978344, 4.979596, 4.980538, 4.981195, 4.981589, 4.981749, 
    4.981706, 4.981493, 4.981143, 4.980695, 4.980181, 4.979634, 4.979084, 
    4.978553, 4.977294, 4.977292, 4.976662, 4.976037, 4.975495, 4.975061, 
    4.975371, 4.975604, 4.975881, 4.976256, 4.976723, 4.97728, 4.97792, 
    4.978625, 4.979328, 4.979919, 4.98132, 4.982853, 4.984545, 4.986426, 
    4.988512, 4.990811, 4.993315, 4.996003, 4.99884, 5.00176, 5.004683, 
    5.0075, 5.010075, 5.012246, 5.013824, 5.0146, 5.014348, 5.012831, 5.009826,
  // momentumX(29,5, 0-49)
    4.978075, 4.97959, 4.980784, 4.981678, 4.982295, 4.98266, 4.9828, 
    4.982745, 4.982529, 4.982182, 4.981737, 4.981228, 4.980682, 4.980126, 
    4.979578, 4.978192, 4.978077, 4.977365, 4.976644, 4.975996, 4.975449, 
    4.975712, 4.975867, 4.976048, 4.976345, 4.976757, 4.977293, 4.977944, 
    4.978681, 4.97939, 4.979939, 4.981371, 4.982926, 4.984634, 4.986518, 
    4.988595, 4.990872, 4.99334, 4.995981, 4.998755, 5.001609, 5.004463, 
    5.007217, 5.009746, 5.0119, 5.013502, 5.014358, 5.014255, 5.012973, 
    5.010293,
  // momentumX(29,6, 0-49)
    4.979375, 4.980821, 4.981953, 4.982794, 4.983367, 4.983699, 4.983816, 
    4.983747, 4.983525, 4.983177, 4.982736, 4.982229, 4.981682, 4.981119, 
    4.980551, 4.979065, 4.978755, 4.977969, 4.97717, 4.976434, 4.975792, 
    4.975995, 4.976058, 4.976129, 4.976338, 4.976693, 4.977218, 4.977898, 
    4.978695, 4.979438, 4.979978, 4.981435, 4.98301, 4.984728, 4.986608, 
    4.988667, 4.990908, 4.993323, 4.995894, 4.998584, 5.00134, 5.004094, 
    5.006751, 5.009197, 5.011295, 5.012885, 5.013788, 5.013808, 5.012739, 
    5.010373,
  // momentumX(29,7, 0-49)
    4.980656, 4.982026, 4.983089, 4.983871, 4.984396, 4.98469, 4.984782, 
    4.984697, 4.984466, 4.984116, 4.983675, 4.98317, 4.982621, 4.982047, 
    4.981458, 4.979904, 4.979315, 4.978468, 4.977612, 4.976809, 4.976092, 
    4.976218, 4.97618, 4.976123, 4.976236, 4.976532, 4.977053, 4.977777, 
    4.978659, 4.979466, 4.980029, 4.981503, 4.983092, 4.984814, 4.986686, 
    4.988718, 4.99091, 4.993259, 4.995742, 4.998327, 5.000965, 5.003592, 
    5.006126, 5.008463, 5.010478, 5.012031, 5.012955, 5.013077, 5.012204, 
    5.010143,
  // momentumX(29,8, 0-49)
    4.981897, 4.983184, 4.984174, 4.984893, 4.985365, 4.98562, 4.985681, 
    4.985578, 4.985337, 4.984982, 4.984541, 4.984036, 4.983485, 4.982903, 
    4.982292, 4.980708, 4.979747, 4.978858, 4.977969, 4.977125, 4.976357, 
    4.976388, 4.976235, 4.976039, 4.976047, 4.976282, 4.976804, 4.977584, 
    4.978576, 4.979469, 4.980087, 4.981573, 4.983167, 4.984883, 4.986736, 
    4.988731, 4.990869, 4.993138, 4.99552, 4.997984, 5.000488, 5.002973, 
    5.005363, 5.007573, 5.009488, 5.010984, 5.011919, 5.012128, 5.011442, 
    5.009677,
  // momentumX(29,9, 0-49)
    4.983086, 4.984283, 4.985192, 4.985842, 4.986258, 4.986469, 4.986499, 
    4.986375, 4.986122, 4.985764, 4.985322, 4.984818, 4.984266, 4.983675, 
    4.983043, 4.981473, 4.980051, 4.97914, 4.978247, 4.977389, 4.976596, 
    4.976516, 4.976236, 4.97589, 4.975786, 4.975957, 4.976483, 4.977327, 
    4.978443, 4.979445, 4.980153, 4.981635, 4.983224, 4.984926, 4.986752, 
    4.988701, 4.990771, 4.992952, 4.995222, 4.997556, 4.999913, 5.002243, 
    5.004482, 5.006552, 5.008358, 5.009792, 5.010726, 5.011018, 5.010513, 
    5.009043,
  // momentumX(29,10, 0-49)
    4.984201, 4.9853, 4.986125, 4.986701, 4.987059, 4.987222, 4.987219, 
    4.987072, 4.986808, 4.986445, 4.986005, 4.985502, 4.984953, 4.984358, 
    4.983712, 4.982196, 4.980223, 4.979319, 4.978451, 4.977612, 4.976825, 
    4.976614, 4.976199, 4.975692, 4.975474, 4.975579, 4.976107, 4.977016, 
    4.978267, 4.979397, 4.980227, 4.981689, 4.983257, 4.984932, 4.986719, 
    4.988612, 4.990606, 4.992688, 4.99484, 4.997035, 4.99924, 5.001411, 
    5.003496, 5.005424, 5.007121, 5.008492, 5.009428, 5.009802, 5.009476, 
    5.008297,
  // momentumX(29,11, 0-49)
    4.985221, 4.986217, 4.986951, 4.987451, 4.987747, 4.987863, 4.987825, 
    4.987659, 4.987381, 4.987016, 4.986578, 4.986081, 4.985535, 4.984943, 
    4.984293, 4.982874, 4.980265, 4.979398, 4.978592, 4.977806, 4.977054, 
    4.9767, 4.976141, 4.975471, 4.975133, 4.975172, 4.9757, 4.976673, 
    4.978061, 4.979329, 4.980305, 4.981731, 4.983263, 4.984897, 4.98663, 
    4.988455, 4.990363, 4.992339, 4.994365, 4.996418, 4.998469, 5.000483, 
    5.002415, 5.004209, 5.005803, 5.007117, 5.008061, 5.008524, 5.008382, 
    5.00749,
  // momentumX(29,12, 0-49)
    4.986129, 4.987016, 4.987657, 4.988077, 4.98831, 4.988379, 4.988306, 
    4.988117, 4.987829, 4.987461, 4.98703, 4.986541, 4.986005, 4.985423, 
    4.984781, 4.983505, 4.980176, 4.979388, 4.978679, 4.977983, 4.977303, 
    4.976789, 4.976083, 4.975247, 4.974793, 4.974764, 4.975285, 4.976314, 
    4.977836, 4.979246, 4.980394, 4.981762, 4.983236, 4.98481, 4.986475, 
    4.98822, 4.99003, 4.991893, 4.99379, 4.9957, 4.997602, 4.999462, 5.00125, 
    5.002921, 5.004425, 5.005697, 5.00666, 5.007222, 5.007267, 5.006666,
  // momentumX(29,13, 0-49)
    4.98691, 4.987683, 4.988225, 4.988565, 4.988734, 4.988751, 4.988646, 
    4.988435, 4.988138, 4.98777, 4.987345, 4.98687, 4.986352, 4.985789, 
    4.985172, 4.984077, 4.97996, 4.979289, 4.978722, 4.978153, 4.97758, 
    4.976897, 4.976046, 4.975048, 4.974481, 4.974383, 4.974892, 4.975965, 
    4.977607, 4.979157, 4.980497, 4.98178, 4.983175, 4.984669, 4.986247, 
    4.987896, 4.989599, 4.991342, 4.993107, 4.994876, 4.996633, 4.998353, 
    5.000012, 5.001576, 5.003008, 5.004256, 5.005257, 5.005929, 5.00617, 
    5.005861,
  // momentumX(29,14, 0-49)
    4.987552, 4.988207, 4.988649, 4.988905, 4.989006, 4.988974, 4.988832, 
    4.988601, 4.988295, 4.987929, 4.987513, 4.987056, 4.986562, 4.986031, 
    4.985457, 4.984582, 4.97962, 4.979108, 4.978724, 4.978326, 4.977896, 
    4.977039, 4.976047, 4.974896, 4.974222, 4.974059, 4.974547, 4.975648, 
    4.977391, 4.979072, 4.980613, 4.981785, 4.983075, 4.984465, 4.985938, 
    4.987476, 4.989061, 4.990677, 4.992309, 4.993942, 4.995565, 4.997159, 
    4.998707, 5.000188, 5.001571, 5.002817, 5.003875, 5.004673, 5.00512, 
    5.005102,
  // momentumX(29,15, 0-49)
    4.988047, 4.988579, 4.988916, 4.989087, 4.989118, 4.989033, 4.988854, 
    4.988601, 4.988286, 4.987922, 4.98752, 4.987084, 4.986623, 4.986136, 
    4.985628, 4.985004, 4.979161, 4.978853, 4.978694, 4.978505, 4.978258, 
    4.977225, 4.976098, 4.97481, 4.974041, 4.973814, 4.974275, 4.975384, 
    4.977204, 4.978997, 4.980742, 4.981776, 4.982933, 4.984197, 4.985542, 
    4.986952, 4.988406, 4.989891, 4.991391, 4.992896, 4.994396, 4.995882, 
    4.997343, 4.998764, 5.000125, 5.001397, 5.002533, 5.003475, 5.004138, 
    5.004411,
  // momentumX(29,16, 0-49)
    4.988392, 4.988796, 4.989022, 4.989101, 4.98906, 4.98892, 4.988703, 
    4.988425, 4.988101, 4.987741, 4.987353, 4.986944, 4.986523, 4.986093, 
    4.985668, 4.985326, 4.978594, 4.978531, 4.978637, 4.978697, 4.978667, 
    4.977459, 4.976213, 4.974801, 4.973953, 4.973667, 4.974092, 4.975191, 
    4.977059, 4.978941, 4.980883, 4.98175, 4.982749, 4.983858, 4.985055, 
    4.986319, 4.987631, 4.988978, 4.990348, 4.991733, 4.993127, 4.994525, 
    4.995924, 4.997314, 4.998682, 5.000005, 5.001247, 5.002351, 5.00324, 
    5.003806,
  // momentumX(29,17, 0-49)
    4.988588, 4.988854, 4.988962, 4.988945, 4.988825, 4.988625, 4.988366, 
    4.988063, 4.987727, 4.98737, 4.986999, 4.986622, 4.986247, 4.985889, 
    4.985566, 4.98553, 4.977942, 4.97816, 4.978563, 4.978907, 4.979125, 
    4.977752, 4.9764, 4.974884, 4.973968, 4.973629, 4.97401, 4.97508, 
    4.976967, 4.978909, 4.981034, 4.981708, 4.982517, 4.983448, 4.984474, 
    4.985574, 4.986732, 4.987938, 4.98918, 4.990454, 4.991757, 4.99309, 
    4.994452, 4.995841, 4.997247, 4.998652, 5.000022, 5.001309, 5.002435, 
    5.003295,
  // momentumX(29,18, 0-49)
    4.988639, 4.988755, 4.988736, 4.98861, 4.988406, 4.988142, 4.987838, 
    4.987507, 4.987159, 4.986805, 4.986453, 4.986112, 4.985792, 4.985513, 
    4.98531, 4.985602, 4.977243, 4.977769, 4.978495, 4.979146, 4.979639, 
    4.978107, 4.976663, 4.97506, 4.974088, 4.973702, 4.974034, 4.975058, 
    4.976934, 4.978906, 4.981187, 4.981641, 4.982238, 4.982964, 4.983794, 
    4.984714, 4.985708, 4.986764, 4.987881, 4.989054, 4.990283, 4.991574, 
    4.992928, 4.994346, 4.995821, 4.997337, 4.998865, 5.000354, 5.001728, 
    5.002884,
  // momentumX(29,19, 0-49)
    4.98855, 4.988499, 4.988338, 4.988094, 4.987796, 4.987462, 4.987109, 
    4.986747, 4.986388, 4.986039, 4.985707, 4.985406, 4.985149, 4.984963, 
    4.984892, 4.98553, 4.976555, 4.977411, 4.978475, 4.979445, 4.980222, 
    4.978542, 4.977019, 4.975341, 4.974323, 4.973892, 4.974168, 4.975128, 
    4.976965, 4.978934, 4.981341, 4.981552, 4.981909, 4.982407, 4.983021, 
    4.98374, 4.984555, 4.985459, 4.98645, 4.98753, 4.988702, 4.989972, 
    4.991343, 4.99282, 4.994395, 4.996053, 4.997765, 4.999477, 5.001114, 
    5.002572,
  // momentumX(29,20, 0-49)
    4.989048, 4.989503, 4.989847, 4.990098, 4.99027, 4.990378, 4.990433, 
    4.990442, 4.990415, 4.99036, 4.990286, 4.990209, 4.990146, 4.990134, 
    4.990227, 0, 4.975359, 4.976153, 4.977207, 4.978203, 4.979018, 4.976952, 
    4.975087, 4.973069, 4.971763, 4.971109, 4.97125, 4.972173, 4.974099, 
    4.976275, 4.979077, 4.979346, 4.979769, 4.980332, 4.98101, 4.981788, 
    4.982655, 4.983606, 4.984644, 4.985774, 4.987006, 4.988348, 4.98981, 
    4.991399, 4.993111, 4.994935, 4.996837, 4.99877, 5.000656, 5.002386,
  // momentumX(29,21, 0-49)
    4.988827, 4.98916, 4.989402, 4.98957, 4.989676, 4.989734, 4.989754, 
    4.989744, 4.989711, 4.98966, 4.9896, 4.989542, 4.989507, 4.989525, 
    4.989647, 0, 4.972302, 4.973264, 4.974558, 4.975825, 4.976907, 4.974704, 
    4.972797, 4.970784, 4.969567, 4.96906, 4.969389, 4.970522, 4.972679, 
    4.975086, 4.978195, 4.978409, 4.978792, 4.979332, 4.980003, 4.980789, 
    4.981676, 4.98266, 4.983741, 4.984922, 4.986211, 4.987618, 4.989153, 
    4.990819, 4.992617, 4.994532, 4.996534, 4.998575, 5.000577, 5.002439,
  // momentumX(29,22, 0-49)
    4.988561, 4.988786, 4.988936, 4.989029, 4.989077, 4.989089, 4.989075, 
    4.989043, 4.988997, 4.988944, 4.988889, 4.988842, 4.988819, 4.988848, 
    4.988978, 0, 4.970036, 4.971129, 4.972622, 4.974118, 4.975419, 4.973063, 
    4.971076, 4.969011, 4.967807, 4.967357, 4.967772, 4.969004, 4.971275, 
    4.973795, 4.977079, 4.977161, 4.977431, 4.977885, 4.978497, 4.979252, 
    4.980139, 4.981151, 4.982288, 4.983549, 4.98494, 4.986465, 4.988132, 
    4.989944, 4.991897, 4.993972, 4.996139, 4.998345, 5.000515, 5.002546,
  // momentumX(29,23, 0-49)
    4.988266, 4.988394, 4.988463, 4.988487, 4.988479, 4.988449, 4.988403, 
    4.988348, 4.988288, 4.988229, 4.988175, 4.988132, 4.988114, 4.988146, 
    4.988268, 0, 4.968285, 4.969466, 4.971102, 4.972762, 4.974215, 4.971715, 
    4.969638, 4.967495, 4.966257, 4.9658, 4.966229, 4.967482, 4.969783, 
    4.972326, 4.975673, 4.975587, 4.97571, 4.976046, 4.976573, 4.977282, 
    4.978163, 4.979208, 4.980416, 4.981785, 4.983315, 4.985008, 4.986862, 
    4.988875, 4.991038, 4.993327, 4.995707, 4.998123, 5.000495, 5.002719,
  // momentumX(29,24, 0-49)
    4.987961, 4.987996, 4.987988, 4.98795, 4.987892, 4.987821, 4.987746, 
    4.98767, 4.987597, 4.987533, 4.987478, 4.987438, 4.987423, 4.987453, 
    4.987559, 0, 4.967278, 4.968503, 4.970228, 4.971992, 4.973543, 4.970967, 
    4.968838, 4.966646, 4.96537, 4.964878, 4.96527, 4.966482, 4.968736, 
    4.971223, 4.974539, 4.974289, 4.974264, 4.97447, 4.974896, 4.975535, 
    4.976382, 4.977432, 4.978685, 4.980134, 4.981779, 4.98362, 4.985648, 
    4.987854, 4.990224, 4.992731, 4.995331, 4.997964, 5.000548, 5.002974,
  // momentumX(29,25, 0-49)
    4.98766, 4.987607, 4.987528, 4.98743, 4.987325, 4.987216, 4.987114, 
    4.987021, 4.986938, 4.986869, 4.986818, 4.986785, 4.986776, 4.986806, 
    4.986895, 0, 4.966704, 4.967937, 4.969695, 4.971504, 4.973098, 4.970532, 
    4.968414, 4.966226, 4.964935, 4.964411, 4.964749, 4.965886, 4.968045, 
    4.970422, 4.973626, 4.973247, 4.973096, 4.973194, 4.973528, 4.974099, 
    4.974905, 4.975947, 4.977223, 4.97873, 4.980465, 4.982426, 4.984601, 
    4.986979, 4.989538, 4.992245, 4.995053, 4.997897, 5.000687, 5.003313,
  // momentumX(29,26, 0-49)
    4.987382, 4.987242, 4.987093, 4.986938, 4.986787, 4.986643, 4.986514, 
    4.986403, 4.986313, 4.986247, 4.986204, 4.986186, 4.986193, 4.986231, 
    4.986312, 0, 4.966497, 4.967708, 4.969454, 4.971251, 4.972836, 4.970378, 
    4.968344, 4.96622, 4.96495, 4.964405, 4.96468, 4.965718, 4.967741, 
    4.969964, 4.972982, 4.972522, 4.972288, 4.972305, 4.972567, 4.97308, 
    4.973845, 4.974867, 4.976147, 4.977685, 4.979478, 4.981522, 4.983808, 
    4.986319, 4.989032, 4.991911, 4.994902, 4.997937, 5.000921, 5.003737,
  // momentumX(29,27, 0-49)
    4.987139, 4.986915, 4.986696, 4.986484, 4.986285, 4.986104, 4.98595, 
    4.985823, 4.985728, 4.985668, 4.985642, 4.98565, 4.985687, 4.985753, 
    4.985845, 0, 4.966663, 4.967835, 4.969529, 4.971269, 4.972798, 4.970535, 
    4.968647, 4.966635, 4.965405, 4.964836, 4.965031, 4.96594, 4.967781, 
    4.969799, 4.972559, 4.972056, 4.971772, 4.971733, 4.971939, 4.972399, 
    4.97312, 4.974112, 4.975377, 4.97692, 4.978742, 4.980838, 4.983202, 
    4.985818, 4.98866, 4.991688, 4.994846, 4.998058, 5.001228, 5.00423,
  // momentumX(29,28, 0-49)
    4.986944, 4.986639, 4.986349, 4.986075, 4.985826, 4.985606, 4.985421, 
    4.985277, 4.985176, 4.985127, 4.985129, 4.985179, 4.985272, 4.985394, 
    4.985533, 0, 4.967456, 4.968589, 4.970207, 4.971852, 4.973289, 4.971285, 
    4.969576, 4.967695, 4.966493, 4.965866, 4.965929, 4.966646, 4.968236, 
    4.969983, 4.972405, 4.971874, 4.97155, 4.971457, 4.971603, 4.971999, 
    4.97266, 4.973596, 4.97482, 4.976341, 4.978161, 4.980283, 4.982701, 
    4.985398, 4.98835, 4.991515, 4.994833, 4.998222, 5.001579, 5.004774,
  // momentumX(29,29, 0-49)
    4.986812, 4.986425, 4.986062, 4.985725, 4.98542, 4.985151, 4.984928, 
    4.984759, 4.984652, 4.984617, 4.984658, 4.984773, 4.984951, 4.985173, 
    4.985413, 0, 4.968573, 4.969682, 4.971219, 4.972744, 4.974048, 4.972317, 
    4.970768, 4.968982, 4.967752, 4.967, 4.966858, 4.967312, 4.968576, 
    4.969975, 4.971971, 4.971394, 4.971013, 4.970857, 4.970938, 4.971271, 
    4.971876, 4.97277, 4.97397, 4.975489, 4.977334, 4.979512, 4.982013, 
    4.984826, 4.987921, 4.991253, 4.994759, 4.998352, 5.001921, 5.005327,
  // momentumX(29,30, 0-49)
    4.986113, 4.985028, 4.983992, 4.98301, 4.982088, 4.981229, 4.980436, 
    4.979713, 4.979061, 4.978491, 4.978013, 4.977649, 4.977439, 4.977439, 
    4.97774, 4.978108, 4.970986, 4.972597, 4.974332, 4.975877, 4.977121, 
    4.975759, 4.974507, 4.972983, 4.97189, 4.971142, 4.970854, 4.971008, 
    4.971807, 4.972627, 4.973881, 4.972935, 4.972168, 4.971625, 4.971332, 
    4.971322, 4.971624, 4.972265, 4.973269, 4.974652, 4.976425, 4.978588, 
    4.981136, 4.984048, 4.987289, 4.990808, 4.994532, 4.998365, 5.002188, 
    5.005852,
  // momentumX(29,31, 0-49)
    4.986139, 4.985011, 4.983933, 4.982914, 4.981956, 4.981061, 4.980238, 
    4.979491, 4.978826, 4.978252, 4.977779, 4.977426, 4.97722, 4.9772, 
    4.977429, 4.977726, 4.970573, 4.971944, 4.973413, 4.974692, 4.97569, 
    4.974526, 4.973392, 4.971966, 4.970906, 4.970163, 4.969861, 4.969983, 
    4.970693, 4.971382, 4.972375, 4.971571, 4.970947, 4.970544, 4.970392, 
    4.970518, 4.970953, 4.971724, 4.972854, 4.974358, 4.976247, 4.978524, 
    4.98118, 4.984198, 4.987542, 4.991161, 4.99498, 4.998902, 5.002809, 
    5.006545,
  // momentumX(29,32, 0-49)
    4.98621, 4.985024, 4.983895, 4.982825, 4.981821, 4.980885, 4.980024, 
    4.979245, 4.978554, 4.977959, 4.97747, 4.977098, 4.97686, 4.97678, 
    4.976899, 4.977179, 4.970335, 4.971414, 4.972563, 4.973532, 4.974247, 
    4.973269, 4.972249, 4.970926, 4.969913, 4.969187, 4.968878, 4.968968, 
    4.969584, 4.97014, 4.970872, 4.970227, 4.969762, 4.969515, 4.969513, 
    4.969784, 4.970358, 4.971261, 4.972516, 4.974138, 4.976139, 4.978522, 
    4.98128, 4.984394, 4.98783, 4.991536, 4.99544, 4.999442, 5.00342, 5.007222,
  // momentumX(29,33, 0-49)
    4.986322, 4.985071, 4.98388, 4.982752, 4.981695, 4.980709, 4.979803, 
    4.978983, 4.978255, 4.977623, 4.977099, 4.976686, 4.976392, 4.976228, 
    4.976206, 4.976455, 4.97019, 4.970946, 4.971748, 4.972381, 4.972796, 
    4.971999, 4.971097, 4.969897, 4.968946, 4.968251, 4.967942, 4.968001, 
    4.96851, 4.968925, 4.969399, 4.968927, 4.968636, 4.968554, 4.968711, 
    4.969135, 4.969853, 4.970891, 4.972271, 4.97401, 4.976117, 4.978599, 
    4.981448, 4.984647, 4.988163, 4.991945, 4.995917, 4.999985, 5.00402, 
    5.007871,
  // momentumX(29,34, 0-49)
    4.986467, 4.98515, 4.983893, 4.982704, 4.981585, 4.980543, 4.979585, 
    4.978714, 4.977937, 4.977258, 4.976682, 4.976209, 4.97584, 4.975573, 
    4.9754, 4.975558, 4.97007, 4.970491, 4.970932, 4.971223, 4.971337, 
    4.970714, 4.969939, 4.968884, 4.968016, 4.967366, 4.967063, 4.967083, 
    4.967473, 4.967741, 4.967969, 4.967685, 4.967576, 4.96767, 4.967996, 
    4.96858, 4.969448, 4.970625, 4.972131, 4.973985, 4.976196, 4.978769, 
    4.981701, 4.984973, 4.988553, 4.992392, 4.996415, 5.000526, 5.0046, 
    5.008479,
  // momentumX(29,35, 0-49)
    4.986632, 4.985251, 4.98393, 4.982677, 4.981496, 4.980392, 4.979373, 
    4.978443, 4.977607, 4.976867, 4.976226, 4.97568, 4.975222, 4.97484, 
    4.974514, 4.974512, 4.969934, 4.970024, 4.970108, 4.97006, 4.969883, 
    4.969428, 4.968791, 4.967904, 4.967138, 4.966548, 4.966253, 4.966227, 
    4.96648, 4.966601, 4.966601, 4.96651, 4.966591, 4.96687, 4.967371, 
    4.968122, 4.969146, 4.970466, 4.972102, 4.974071, 4.976381, 4.979041, 
    4.982045, 4.985377, 4.989005, 4.99288, 4.996932, 5.001062, 5.005144, 
    5.009022,
  // momentumX(29,36, 0-49)
    4.986797, 4.985363, 4.983984, 4.98267, 4.981424, 4.980255, 4.97917, 
    4.978174, 4.977268, 4.976458, 4.97574, 4.97511, 4.974553, 4.974052, 
    4.973577, 4.973351, 4.969756, 4.969531, 4.96927, 4.968902, 4.968448, 
    4.968158, 4.967667, 4.966969, 4.966328, 4.965811, 4.965522, 4.965443, 
    4.965545, 4.965516, 4.965311, 4.965418, 4.965693, 4.96616, 4.966842, 
    4.967765, 4.968948, 4.970416, 4.972183, 4.974266, 4.976675, 4.979414, 
    4.98248, 4.985857, 4.989515, 4.993406, 4.99746, 5.001577, 5.005634, 
    5.009474,
  // momentumX(29,37, 0-49)
    4.986938, 4.985464, 4.984036, 4.982665, 4.981359, 4.980126, 4.978973, 
    4.977904, 4.976924, 4.976033, 4.97523, 4.974505, 4.973844, 4.973222, 
    4.972605, 4.972109, 4.969525, 4.969004, 4.968421, 4.967756, 4.967048, 
    4.966916, 4.966578, 4.966092, 4.965594, 4.965162, 4.964882, 4.964739, 
    4.964676, 4.9645, 4.964114, 4.96442, 4.964892, 4.965548, 4.966413, 
    4.96751, 4.968857, 4.970472, 4.972372, 4.974567, 4.97707, 4.979882, 
    4.983001, 4.986409, 4.990077, 4.993959, 4.997983, 5.002053, 5.006046, 
    5.009804,
  // momentumX(29,38, 0-49)
    4.987028, 4.985529, 4.984065, 4.982647, 4.981288, 4.979993, 4.978771, 
    4.977629, 4.976569, 4.975593, 4.974696, 4.973871, 4.973101, 4.972361, 
    4.971611, 4.970821, 4.969233, 4.968444, 4.967564, 4.96663, 4.965697, 
    4.965714, 4.965539, 4.96528, 4.964942, 4.964607, 4.964337, 4.964119, 
    4.963884, 4.963566, 4.96303, 4.963531, 4.964195, 4.965038, 4.966087, 
    4.967357, 4.968866, 4.970628, 4.972659, 4.974966, 4.977559, 4.980438, 
    4.983595, 4.98702, 4.990678, 4.994521, 4.998483, 5.002466, 5.006349, 
    5.009973,
  // momentumX(29,39, 0-49)
    4.98703, 4.985528, 4.984045, 4.982595, 4.981189, 4.97984, 4.978554, 
    4.977337, 4.976196, 4.975132, 4.974139, 4.97321, 4.972332, 4.971474, 
    4.970599, 4.969515, 4.96888, 4.967854, 4.966705, 4.965531, 4.964404, 
    4.964564, 4.964558, 4.964538, 4.964377, 4.964149, 4.963889, 4.963593, 
    4.96318, 4.96273, 4.962073, 4.962762, 4.963613, 4.964639, 4.965863, 
    4.967302, 4.96897, 4.970879, 4.973037, 4.975451, 4.978129, 4.981064, 
    4.984251, 4.987672, 4.991296, 4.995074, 4.998935, 5.002787, 5.006506, 
    5.009941,
  // momentumX(29,40, 0-49)
    4.986917, 4.985433, 4.98395, 4.982483, 4.981046, 4.979649, 4.978304, 
    4.977018, 4.975799, 4.974646, 4.973557, 4.972527, 4.971539, 4.970568, 
    4.969579, 4.968217, 4.968469, 4.967233, 4.965849, 4.964469, 4.963177, 
    4.963475, 4.963636, 4.963868, 4.963894, 4.963784, 4.963535, 4.963162, 
    4.962571, 4.962003, 4.961255, 4.962122, 4.963151, 4.964351, 4.965744, 
    4.967346, 4.969165, 4.971212, 4.973492, 4.976008, 4.978761, 4.981743, 
    4.984945, 4.988344, 4.991908, 4.995585, 4.999307, 5.002978, 5.006479, 
    5.00966,
  // momentumX(29,41, 0-49)
    4.986656, 4.985214, 4.983752, 4.982286, 4.980833, 4.979402, 4.978008, 
    4.976662, 4.975368, 4.97413, 4.97295, 4.971819, 4.970726, 4.969647, 
    4.968551, 4.96694, 4.968, 4.966581, 4.964995, 4.963443, 4.96202, 
    4.962448, 4.962779, 4.963267, 4.963491, 4.963505, 4.963273, 4.962823, 
    4.962065, 4.961395, 4.960584, 4.96162, 4.962814, 4.964176, 4.965727, 
    4.967481, 4.969442, 4.971618, 4.974011, 4.976619, 4.979436, 4.98245, 
    4.98565, 4.989006, 4.992481, 4.996022, 4.99956, 5.002998, 5.00622, 5.00908,
  // momentumX(29,42, 0-49)
    4.986219, 4.984845, 4.983426, 4.981982, 4.980528, 4.979081, 4.977652, 
    4.976253, 4.974894, 4.973581, 4.972313, 4.971088, 4.969896, 4.968716, 
    4.96752, 4.965698, 4.967477, 4.965904, 4.964147, 4.962456, 4.960933, 
    4.961483, 4.961984, 4.962727, 4.963152, 4.963299, 4.96309, 4.962575, 
    4.961663, 4.96091, 4.960064, 4.961257, 4.962603, 4.964114, 4.96581, 
    4.967701, 4.969793, 4.972085, 4.974578, 4.977262, 4.980129, 4.98316, 
    4.986334, 4.989621, 4.992977, 4.996344, 4.99965, 5.0028, 5.00568, 5.00815,
  // momentumX(29,43, 0-49)
    4.985586, 4.984303, 4.982952, 4.981551, 4.980116, 4.978669, 4.977219, 
    4.975782, 4.97437, 4.97299, 4.971644, 4.970334, 4.969049, 4.967778, 
    4.966492, 4.964496, 4.966899, 4.965197, 4.963301, 4.961505, 4.959913, 
    4.960582, 4.961247, 4.96224, 4.962868, 4.963152, 4.962977, 4.962408, 
    4.961366, 4.960551, 4.959695, 4.961031, 4.962516, 4.964162, 4.965988, 
    4.968001, 4.970206, 4.972599, 4.975173, 4.977917, 4.980814, 4.983839, 
    4.986966, 4.990153, 4.993352, 4.996504, 4.999529, 5.002333, 5.004804, 
    5.006812,
  // momentumX(29,44, 0-49)
    4.984741, 4.983572, 4.98231, 4.980974, 4.979583, 4.978152, 4.9767, 
    4.975242, 4.973791, 4.972355, 4.970943, 4.969557, 4.968193, 4.966837, 
    4.96547, 4.96334, 4.966269, 4.964459, 4.962457, 4.960586, 4.958953, 
    4.959734, 4.960559, 4.961791, 4.962621, 4.963047, 4.962915, 4.962311, 
    4.961167, 4.960318, 4.959472, 4.96094, 4.96255, 4.964314, 4.966252, 
    4.968369, 4.970668, 4.973141, 4.975777, 4.978558, 4.981461, 4.984454, 
    4.987502, 4.990557, 4.993561, 4.996449, 4.999139, 5.001537, 5.003535, 
    5.00501,
  // momentumX(29,45, 0-49)
    4.983676, 4.982643, 4.981495, 4.980247, 4.978919, 4.977528, 4.976092, 
    4.974628, 4.973153, 4.971678, 4.970212, 4.968764, 4.967327, 4.965899, 
    4.964459, 4.962228, 4.965582, 4.963693, 4.96161, 4.959693, 4.958048, 
    4.958934, 4.95991, 4.961367, 4.962389, 4.962958, 4.962886, 4.962271, 
    4.961058, 4.960199, 4.959386, 4.960973, 4.962695, 4.964563, 4.966595, 
    4.968796, 4.971167, 4.973697, 4.976369, 4.979159, 4.982038, 4.984967, 
    4.987901, 4.990783, 4.99355, 4.996124, 4.998423, 5.000354, 5.001812, 
    5.002688,
  // momentumX(29,46, 0-49)
    4.982392, 4.981516, 4.980502, 4.979363, 4.978121, 4.976789, 4.97539, 
    4.973942, 4.972459, 4.970959, 4.969454, 4.967954, 4.96646, 4.964968, 
    4.963467, 4.961162, 4.96484, 4.962892, 4.96076, 4.958823, 4.957186, 
    4.958171, 4.959288, 4.960949, 4.962153, 4.962865, 4.962866, 4.962266, 
    4.961024, 4.960183, 4.959423, 4.961119, 4.962938, 4.964893, 4.967002, 
    4.969267, 4.971686, 4.974245, 4.976924, 4.979692, 4.982513, 4.985339, 
    4.988117, 4.990781, 4.993258, 4.995465, 4.997318, 4.998721, 4.999578, 
    4.999793,
  // momentumX(29,47, 0-49)
    4.980901, 4.9802, 4.979339, 4.97833, 4.977193, 4.975943, 4.9746, 
    4.973184, 4.971713, 4.970206, 4.968677, 4.967138, 4.965598, 4.964054, 
    4.962501, 4.960147, 4.964045, 4.96206, 4.959902, 4.957967, 4.956358, 
    4.957434, 4.958677, 4.960518, 4.961888, 4.96274, 4.962831, 4.962277, 
    4.961047, 4.960255, 4.959564, 4.961359, 4.963265, 4.965293, 4.967459, 
    4.969764, 4.972204, 4.974763, 4.977415, 4.980123, 4.982846, 4.985526, 
    4.988099, 4.990493, 4.992628, 4.994412, 4.995758, 4.996574, 4.996771, 
    4.996272,
  // momentumX(29,48, 0-49)
    4.979223, 4.978709, 4.978018, 4.977159, 4.976146, 4.974998, 4.973732, 
    4.972368, 4.970926, 4.969428, 4.967888, 4.966326, 4.96475, 4.963166, 
    4.961571, 4.959184, 4.963201, 4.961198, 4.959035, 4.957121, 4.955557, 
    4.956709, 4.958065, 4.960053, 4.961572, 4.96256, 4.962756, 4.96228, 
    4.961107, 4.960392, 4.959789, 4.961674, 4.963654, 4.965738, 4.967942, 
    4.970265, 4.972701, 4.975228, 4.977816, 4.980423, 4.983, 4.985481, 
    4.987796, 4.989864, 4.991597, 4.992898, 4.993679, 4.993851, 4.993337, 
    4.992082,
  // momentumX(29,49, 0-49)
    4.977364, 4.976999, 4.976442, 4.975697, 4.974771, 4.973678, 4.972433, 
    4.97105, 4.96955, 4.967954, 4.966277, 4.964537, 4.96275, 4.960918, 
    4.959042, 4.955583, 4.965085, 4.962095, 4.958641, 4.955575, 4.95313, 
    4.956073, 4.959288, 4.963607, 4.966753, 4.968592, 4.96859, 4.966987, 
    4.963706, 4.96112, 4.958558, 4.960826, 4.963123, 4.965455, 4.967843, 
    4.970289, 4.972789, 4.975318, 4.977843, 4.980316, 4.982681, 4.984867, 
    4.986794, 4.988374, 4.989514, 4.990113, 4.990091, 4.989372, 4.987904, 
    4.98567 ;

 momentumY =
  // momentumY(0,0, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumY(0,1, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumY(0,2, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumY(0,3, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumY(0,4, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumY(0,5, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumY(0,6, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumY(0,7, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumY(0,8, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumY(0,9, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumY(0,10, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumY(0,11, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumY(0,12, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumY(0,13, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumY(0,14, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumY(0,15, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumY(0,16, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumY(0,17, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumY(0,18, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumY(0,19, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumY(0,20, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 0, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumY(0,21, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 0, 5, 5, 5, 5, 5, 5, 5, 10, 
    10, 10, 10, 10, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5,
  // momentumY(0,22, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 0, 5, 5, 5, 5, 5, 5, 10, 10, 
    10, 10, 10, 10, 10, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5,
  // momentumY(0,23, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 0, 5, 5, 5, 5, 5, 10, 10, 
    10, 10, 10, 10, 10, 10, 10, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5,
  // momentumY(0,24, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 0, 5, 5, 5, 5, 5, 10, 10, 
    10, 10, 10, 10, 10, 10, 10, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5,
  // momentumY(0,25, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 0, 5, 5, 5, 5, 5, 10, 10, 
    10, 10, 10, 10, 10, 10, 10, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5,
  // momentumY(0,26, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 0, 5, 5, 5, 5, 5, 10, 10, 
    10, 10, 10, 10, 10, 10, 10, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5,
  // momentumY(0,27, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 0, 5, 5, 5, 5, 5, 10, 10, 
    10, 10, 10, 10, 10, 10, 10, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5,
  // momentumY(0,28, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 0, 5, 5, 5, 5, 5, 5, 10, 10, 
    10, 10, 10, 10, 10, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5,
  // momentumY(0,29, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 0, 5, 5, 5, 5, 5, 5, 5, 10, 
    10, 10, 10, 10, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5,
  // momentumY(0,30, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumY(0,31, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumY(0,32, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumY(0,33, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumY(0,34, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumY(0,35, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumY(0,36, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumY(0,37, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumY(0,38, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumY(0,39, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumY(0,40, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumY(0,41, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumY(0,42, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumY(0,43, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumY(0,44, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumY(0,45, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumY(0,46, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumY(0,47, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumY(0,48, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumY(0,49, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumY(1,0, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumY(1,1, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumY(1,2, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumY(1,3, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumY(1,4, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumY(1,5, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumY(1,6, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumY(1,7, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumY(1,8, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumY(1,9, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5.000001, 5.000003, 5.000003, 5.000003, 5.000003, 5.000003, 5.000001, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumY(1,10, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 
    5.00001, 5.000023, 5.000029, 5.00003, 5.000029, 5.000023, 5.00001, 
    5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumY(1,11, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000005, 
    5.000022, 5.000071, 5.000165, 5.000208, 5.000218, 5.000208, 5.000165, 
    5.000071, 5.000022, 5.000005, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5,
  // momentumY(1,12, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000009, 
    5.000041, 5.000161, 5.000472, 5.00103, 5.001293, 5.001361, 5.001293, 
    5.00103, 5.000472, 5.000161, 5.000041, 5.000009, 5.000001, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumY(1,13, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000013, 
    5.000065, 5.00028, 5.000989, 5.002667, 5.005479, 5.00688, 5.007271, 
    5.00688, 5.005479, 5.002667, 5.000989, 5.00028, 5.000065, 5.000013, 
    5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumY(1,14, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000016, 
    5.000087, 5.000412, 5.001609, 5.005196, 5.012874, 5.024823, 5.031068, 
    5.032917, 5.031068, 5.024823, 5.012874, 5.005196, 5.001609, 5.000412, 
    5.000087, 5.000016, 5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumY(1,15, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000018, 
    5.000104, 5.000527, 5.002232, 5.007843, 5.023126, 5.05233, 5.093832, 
    5.116333, 5.123362, 5.116333, 5.093832, 5.05233, 5.023126, 5.007843, 
    5.002232, 5.000527, 5.000104, 5.000018, 5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5,
  // momentumY(1,16, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000016, 5.000111, 
    5.000595, 5.002696, 5.010195, 5.032046, 5.08562, 5.174296, 5.284347, 
    5.345138, 5.365025, 5.345138, 5.284347, 5.174296, 5.08562, 5.032046, 
    5.010195, 5.002696, 5.000595, 5.00011, 5.000018, 5.000002, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5,
  // momentumY(1,17, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000013, 5.000091, 
    5.000609, 5.00287, 5.011568, 5.038834, 5.107607, 5.255316, 5.45458, 
    5.654781, 5.766831, 5.805127, 5.766831, 5.654781, 5.45458, 5.255316, 
    5.107607, 5.038834, 5.011568, 5.002866, 5.000595, 5.000104, 5.000016, 
    5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumY(1,18, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000008, 5.00006, 5.000425, 
    5.002811, 5.011596, 5.041329, 5.121252, 5.288161, 5.587032, 5.889495, 
    6.114048, 6.247925, 6.296353, 6.247925, 6.114048, 5.889495, 5.587032, 
    5.288161, 5.121252, 5.041325, 5.011568, 5.002696, 5.000527, 5.000087, 
    5.000013, 5.000001, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumY(1,19, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000003, 5.000028, 5.000218, 
    5.001533, 5.011003, 5.039038, 5.121291, 5.303221, 5.596775, 6.011393, 
    6.30257, 6.444544, 6.550306, 6.591668, 6.550305, 6.444544, 6.30257, 
    6.011393, 5.596775, 5.303215, 5.121252, 5.038834, 5.010195, 5.002232, 
    5.000412, 5.000065, 5.000009, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumY(1,20, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000014, 0, 5.039814, 
    5.109214, 5.288445, 5.596817, 5.95014, 6.326973, 6.498679, 6.541141, 
    6.600243, 6.624728, 6.600243, 6.541141, 6.498679, 6.326972, 5.950134, 
    5.596775, 5.288161, 5.107607, 5.032046, 5.007843, 5.001609, 5.00028, 
    5.000041, 5.000005, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumY(1,21, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 0, 5.108829, 
    5.260567, 5.588036, 6.011554, 6.326994, 6.546953, 6.566364, 6.535832, 
    6.558554, 6.576564, 6.558554, 6.535832, 6.566363, 6.546951, 6.326972, 
    6.011393, 5.587032, 5.255316, 5.08562, 5.023126, 5.005196, 5.000989, 
    5.000161, 5.000022, 5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumY(1,22, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 0, 5.226802, 5.467532, 
    5.892158, 6.303021, 6.498741, 6.56637, 6.621973, 6.765517, 6.920608, 
    6.987292, 6.920608, 6.765517, 6.621973, 6.566362, 6.498679, 6.30257, 
    5.889495, 5.45458, 5.174296, 5.05233, 5.012874, 5.002667, 5.000472, 
    5.000071, 5.00001, 5.000001, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumY(1,23, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 0, 5.378377, 5.679589, 
    6.119381, 6.445471, 6.541272, 6.535846, 6.765518, 7.138705, 7.442398, 
    7.559381, 7.442398, 7.138703, 6.765517, 6.535831, 6.541141, 6.444544, 
    6.114048, 5.654781, 5.284347, 5.093832, 5.024823, 5.005479, 5.00103, 
    5.000165, 5.000023, 5.000003, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumY(1,24, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 0, 5.461733, 5.797845, 
    6.254579, 6.551452, 6.600401, 6.558572, 6.920609, 7.442399, 7.841739, 
    7.990802, 7.841739, 7.442398, 6.920608, 6.558555, 6.600243, 6.550306, 
    6.247925, 5.766831, 5.345138, 5.116333, 5.031068, 5.00688, 5.001293, 
    5.000208, 5.000029, 5.000003, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumY(1,25, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 0, 5.488677, 5.83798, 
    6.303374, 6.592873, 6.624895, 6.576583, 6.987293, 7.559382, 7.990802, 
    8.150589, 7.990803, 7.559381, 6.987291, 6.576564, 6.624729, 6.591668, 
    6.296353, 5.805127, 5.365025, 5.123362, 5.032917, 5.007271, 5.001361, 
    5.000218, 5.00003, 5.000003, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumY(1,26, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 0, 5.461732, 5.797844, 
    6.254579, 6.551452, 6.600401, 6.558572, 6.920609, 7.442398, 7.841739, 
    7.990802, 7.841739, 7.442398, 6.920608, 6.558555, 6.600243, 6.550306, 
    6.247925, 5.766831, 5.345138, 5.116333, 5.031068, 5.00688, 5.001293, 
    5.000208, 5.000029, 5.000003, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumY(1,27, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 0, 5.378368, 
    5.679588, 6.119381, 6.445471, 6.541272, 6.535846, 6.765518, 7.138705, 
    7.442398, 7.55938, 7.442398, 7.138704, 6.765517, 6.535832, 6.541142, 
    6.444544, 6.114048, 5.654781, 5.284347, 5.093832, 5.024823, 5.005479, 
    5.00103, 5.000165, 5.000023, 5.000003, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumY(1,28, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000009, 0, 5.226734, 
    5.467518, 5.892155, 6.303021, 6.498741, 6.56637, 6.621974, 6.765516, 
    6.920608, 6.987291, 6.920608, 6.765516, 6.621973, 6.566363, 6.498679, 
    6.30257, 5.889495, 5.45458, 5.174296, 5.05233, 5.012874, 5.002667, 
    5.000472, 5.000071, 5.00001, 5.000001, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumY(1,29, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000013, 5.00007, 0, 
    5.108382, 5.260472, 5.588021, 6.011552, 6.326994, 6.546954, 6.566364, 
    6.535832, 6.558555, 6.576563, 6.558555, 6.535832, 6.566363, 6.546951, 
    6.326972, 6.011393, 5.587032, 5.255316, 5.08562, 5.023126, 5.005196, 
    5.000989, 5.000161, 5.000022, 5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumY(1,30, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000017, 5.000138, 5.000946, 
    5.005786, 5.03459, 5.108321, 5.288314, 5.5968, 5.950139, 6.326973, 
    6.49868, 6.541142, 6.600243, 6.624728, 6.600243, 6.541142, 6.498679, 
    6.326972, 5.950134, 5.596775, 5.288161, 5.107607, 5.032046, 5.007843, 
    5.001609, 5.00028, 5.000041, 5.000005, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumY(1,31, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000005, 5.000042, 5.000306, 
    5.001886, 5.010614, 5.038951, 5.121276, 5.303219, 5.596775, 6.011393, 
    6.30257, 6.444544, 6.550306, 6.591668, 6.550306, 6.444544, 6.30257, 
    6.011393, 5.596775, 5.303215, 5.121252, 5.038834, 5.010195, 5.002232, 
    5.000412, 5.000065, 5.000009, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumY(1,32, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000009, 5.000072, 5.000477, 
    5.002755, 5.011584, 5.041328, 5.121252, 5.288161, 5.587032, 5.889495, 
    6.114048, 6.247925, 6.296353, 6.247925, 6.114048, 5.889495, 5.587032, 
    5.288161, 5.121252, 5.041325, 5.011568, 5.002696, 5.000527, 5.000087, 
    5.000013, 5.000001, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumY(1,33, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000014, 5.000097, 
    5.000602, 5.002868, 5.011568, 5.038834, 5.107607, 5.255316, 5.45458, 
    5.654781, 5.766831, 5.805127, 5.766831, 5.654781, 5.45458, 5.255316, 
    5.107607, 5.038834, 5.011568, 5.002866, 5.000595, 5.000104, 5.000016, 
    5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumY(1,34, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000017, 5.00011, 
    5.000595, 5.002696, 5.010195, 5.032046, 5.08562, 5.174296, 5.284347, 
    5.345138, 5.365025, 5.345138, 5.284347, 5.174296, 5.08562, 5.032046, 
    5.010195, 5.002696, 5.000595, 5.00011, 5.000018, 5.000002, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5,
  // momentumY(1,35, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000018, 
    5.000104, 5.000527, 5.002232, 5.007843, 5.023126, 5.05233, 5.093832, 
    5.116333, 5.123362, 5.116333, 5.093832, 5.05233, 5.023126, 5.007843, 
    5.002232, 5.000527, 5.000104, 5.000018, 5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5,
  // momentumY(1,36, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000016, 
    5.000087, 5.000412, 5.001609, 5.005196, 5.012874, 5.024823, 5.031068, 
    5.032917, 5.031068, 5.024823, 5.012874, 5.005196, 5.001609, 5.000412, 
    5.000087, 5.000016, 5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumY(1,37, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000013, 
    5.000065, 5.00028, 5.000989, 5.002667, 5.005479, 5.00688, 5.007271, 
    5.00688, 5.005479, 5.002667, 5.000989, 5.00028, 5.000065, 5.000013, 
    5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumY(1,38, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000009, 
    5.000041, 5.000161, 5.000472, 5.00103, 5.001293, 5.001361, 5.001293, 
    5.00103, 5.000472, 5.000161, 5.000041, 5.000009, 5.000001, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumY(1,39, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000005, 
    5.000022, 5.000071, 5.000165, 5.000208, 5.000218, 5.000208, 5.000165, 
    5.000071, 5.000022, 5.000005, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5,
  // momentumY(1,40, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 
    5.00001, 5.000023, 5.000029, 5.00003, 5.000029, 5.000023, 5.00001, 
    5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumY(1,41, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5.000001, 5.000003, 5.000003, 5.000003, 5.000003, 5.000003, 5.000001, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumY(1,42, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumY(1,43, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumY(1,44, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumY(1,45, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumY(1,46, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumY(1,47, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumY(1,48, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumY(1,49, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumY(2,0, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumY(2,1, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumY(2,2, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumY(2,3, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5.000001, 5.000001, 5.000001, 5.000001, 5.000001, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumY(2,4, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 
    5.000003, 5.000006, 5.000008, 5.000009, 5.000008, 5.000006, 5.000003, 
    5.000001, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumY(2,5, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 
    5.000003, 5.000009, 5.000018, 5.00003, 5.000037, 5.000041, 5.000037, 
    5.00003, 5.000018, 5.000009, 5.000003, 5.000001, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumY(2,6, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000008, 
    5.00002, 5.000044, 5.000084, 5.000135, 5.000167, 5.000179, 5.000167, 
    5.000135, 5.000084, 5.000044, 5.00002, 5.000008, 5.000002, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumY(2,7, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000004, 5.000013, 
    5.000036, 5.000087, 5.000192, 5.000359, 5.000562, 5.000698, 5.000745, 
    5.000698, 5.000562, 5.000359, 5.000192, 5.000087, 5.000036, 5.000013, 
    5.000004, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumY(2,8, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000005, 
    5.000019, 5.000055, 5.000149, 5.000361, 5.000768, 5.001396, 5.002146, 
    5.002654, 5.002829, 5.002654, 5.002146, 5.001396, 5.000768, 5.000361, 
    5.000149, 5.000055, 5.000019, 5.000005, 5.000001, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5,
  // momentumY(2,9, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000007, 5.000025, 
    5.00008, 5.00023, 5.000596, 5.001375, 5.002819, 5.004971, 5.00749, 
    5.009201, 5.009799, 5.009201, 5.00749, 5.004971, 5.002819, 5.001375, 
    5.000596, 5.00023, 5.00008, 5.000025, 5.000007, 5.000001, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5,
  // momentumY(2,10, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000008, 5.000031, 
    5.000104, 5.000319, 5.000876, 5.002162, 5.004771, 5.009418, 5.016093, 
    5.023739, 5.028931, 5.030761, 5.028931, 5.023739, 5.016093, 5.009418, 
    5.004771, 5.002162, 5.000876, 5.000319, 5.000104, 5.000031, 5.000008, 
    5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumY(2,11, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.00001, 5.000034, 
    5.000126, 5.000408, 5.001172, 5.003046, 5.007127, 5.014987, 5.028435, 
    5.046975, 5.067611, 5.08152, 5.086449, 5.08152, 5.067611, 5.046975, 
    5.028435, 5.014987, 5.007127, 5.003045, 5.001171, 5.000405, 5.000127, 
    5.000036, 5.00001, 5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumY(2,12, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000009, 5.000036, 5.000136, 
    5.000466, 5.001442, 5.003905, 5.00958, 5.021203, 5.042273, 5.076715, 
    5.121716, 5.169673, 5.201324, 5.212531, 5.201324, 5.169673, 5.121716, 
    5.076715, 5.042273, 5.021201, 5.009576, 5.003897, 5.00143, 5.000474, 
    5.000143, 5.000039, 5.00001, 5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumY(2,13, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000008, 5.000033, 5.000133, 
    5.000481, 5.00157, 5.004634, 5.011772, 5.027131, 5.05641, 5.105655, 
    5.181499, 5.273223, 5.364344, 5.422204, 5.4425, 5.422204, 5.364344, 
    5.273223, 5.181498, 5.105653, 5.056403, 5.02711, 5.011728, 5.004572, 
    5.001609, 5.000513, 5.000149, 5.000039, 5.00001, 5.000002, 5, 5, 5, 5, 5, 
    5, 5, 5, 5,
  // momentumY(2,14, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000007, 5.000029, 5.000118, 5.000446, 
    5.001536, 5.004781, 5.013485, 5.031936, 5.068588, 5.132482, 5.229629, 
    5.367397, 5.516597, 5.650199, 5.73082, 5.75868, 5.73082, 5.650199, 
    5.516597, 5.367393, 5.229616, 5.132443, 5.068489, 5.031737, 5.013205, 
    5.004946, 5.001672, 5.000513, 5.000143, 5.000036, 5.000008, 5.000001, 5, 
    5, 5, 5, 5, 5, 5, 5,
  // momentumY(2,15, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000004, 5.000021, 5.000093, 5.000368, 
    5.001338, 5.004398, 5.013077, 5.035445, 5.07743, 5.152986, 5.270136, 
    5.425341, 5.623005, 5.808567, 5.954159, 6.038265, 6.066943, 6.038265, 
    5.954158, 5.808562, 5.622989, 5.425284, 5.269968, 5.152572, 5.076609, 
    5.034278, 5.01373, 5.004946, 5.001609, 5.000474, 5.000127, 5.000031, 
    5.000007, 5.000001, 5, 5, 5, 5, 5, 5, 5,
  // momentumY(2,16, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000014, 5.000063, 5.000268, 5.001024, 
    5.003561, 5.011195, 5.031907, 5.083897, 5.166404, 5.297246, 5.471339, 
    5.663941, 5.881144, 6.054009, 6.170801, 6.238191, 6.261086, 6.23819, 
    6.170798, 6.053992, 5.881079, 5.663725, 5.470706, 5.295689, 5.163324, 
    5.079466, 5.034278, 5.013205, 5.004572, 5.00143, 5.000405, 5.000104, 
    5.000025, 5.000005, 5, 5, 5, 5, 5, 5, 5,
  // momentumY(2,17, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000008, 5.000038, 5.000165, 5.00067, 
    5.002472, 5.008275, 5.024992, 5.068762, 5.178341, 5.314689, 5.498798, 
    5.701071, 5.878989, 6.057094, 6.174425, 6.241654, 6.28508, 6.300066, 
    6.285078, 6.24164, 6.174369, 6.056881, 5.878283, 5.699006, 5.493689, 
    5.304491, 5.163324, 5.076609, 5.031737, 5.011728, 5.003897, 5.001171, 
    5.000319, 5.00008, 5.000019, 5.000004, 5, 5, 5, 5, 5, 5,
  // momentumY(2,18, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5.000003, 5.000017, 5.000082, 5.000356, 5.001401, 
    5.005028, 5.016359, 5.047846, 5.129076, 5.339933, 5.523062, 5.725195, 
    5.900149, 6.010222, 6.107472, 6.153584, 6.174073, 6.196599, 6.204854, 
    6.196589, 6.174033, 6.153419, 6.106858, 6.008182, 5.894237, 5.710595, 
    5.493689, 5.295689, 5.152572, 5.068489, 5.02711, 5.009576, 5.003045, 
    5.000876, 5.00023, 5.000055, 5.000013, 5.000002, 5, 5, 5, 5, 5,
  // momentumY(2,19, 0-49)
    5, 5, 5, 5, 5, 5, 5.000001, 5.000007, 5.000029, 5.000135, 5.000575, 
    5.002245, 5.008015, 5.025926, 5.074886, 5.206708, 5.580922, 5.772137, 
    5.930871, 6.024444, 6.039964, 6.04226, 6.020387, 6.004436, 6.009708, 
    6.012484, 6.009684, 6.004327, 6.019951, 6.040654, 6.034697, 6.009424, 
    5.894236, 5.699005, 5.470706, 5.269968, 5.132443, 5.056403, 5.021201, 
    5.007127, 5.002162, 5.000596, 5.000149, 5.000036, 5.000008, 5.000001, 5, 
    5, 5, 5,
  // momentumY(2,20, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5.000001, 5.00001, 5.000042, 5.000171, 5.000613, 
    5.001966, 5.005518, 5.013143, 0, 6.070654, 6.10031, 6.109229, 6.073961, 
    5.989838, 5.897338, 5.812802, 5.764136, 5.750331, 5.746961, 5.750273, 
    5.763871, 5.811723, 5.893331, 5.976495, 6.034697, 6.008182, 5.878282, 
    5.663725, 5.425284, 5.229616, 5.105653, 5.042273, 5.014987, 5.004771, 
    5.001375, 5.000361, 5.000087, 5.00002, 5.000003, 5, 5, 5, 5,
  // momentumY(2,21, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5.000003, 5.000014, 5.000054, 5.000195, 5.00063, 
    5.001772, 5.004181, 0, 6.513035, 6.426273, 6.282675, 6.110457, 5.917133, 
    5.702082, 5.514227, 5.387189, 5.318944, 5.296926, 5.318848, 5.386738, 
    5.51234, 5.694969, 5.893331, 6.040654, 6.106857, 6.056882, 5.88108, 
    5.622988, 5.367393, 5.181498, 5.076715, 5.028435, 5.009418, 5.002819, 
    5.000768, 5.000192, 5.000044, 5.000009, 5.000001, 5, 5, 5,
  // momentumY(2,22, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000004, 5.000016, 5.000055, 5.000182, 
    5.000515, 5.001205, 0, 6.890601, 6.696692, 6.413081, 6.125101, 5.847679, 
    5.523096, 5.231614, 5.02129, 4.898302, 4.858558, 4.898164, 5.020628, 
    5.228783, 5.512339, 5.811723, 6.019951, 6.153419, 6.174369, 6.053992, 
    5.808561, 5.516597, 5.273223, 5.121716, 5.046975, 5.016093, 5.004971, 
    5.001396, 5.000359, 5.000084, 5.000018, 5.000003, 5, 5, 5,
  // momentumY(2,23, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000004, 5.000016, 5.000049, 5.000141, 
    5.000327, 0, 7.175317, 6.901651, 6.513165, 6.143483, 5.81144, 5.400992, 
    5.024344, 4.753988, 4.602839, 4.55656, 4.602668, 4.753143, 5.020628, 
    5.386737, 5.76387, 6.004326, 6.174033, 6.241639, 6.170797, 5.954158, 
    5.650199, 5.364344, 5.169673, 5.067611, 5.023739, 5.00749, 5.002146, 
    5.000562, 5.000135, 5.00003, 5.000006, 5.000001, 5, 5,
  // momentumY(2,24, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000006, 5.00002, 5.000057, 5.000128, 
    0, 7.33971, 7.028852, 6.586917, 6.171556, 5.805634, 5.335411, 4.902411, 
    4.603594, 4.448595, 4.40392, 4.448415, 4.602663, 4.89816, 5.318843, 
    5.750269, 6.009683, 6.196589, 6.285078, 6.23819, 6.038265, 5.73082, 
    5.422204, 5.201324, 5.08152, 5.028931, 5.009201, 5.002654, 5.000698, 
    5.000167, 5.000037, 5.000008, 5.000001, 5, 5,
  // momentumY(2,25, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000003, 5.000013, 5.000041, 5.000108, 
    5.000237, 0, 7.394997, 7.072412, 6.612961, 6.182293, 5.805012, 5.31426, 
    4.862948, 4.55748, 4.40407, 4.360934, 4.403889, 4.556526, 4.858529, 
    5.296904, 5.746947, 6.012478, 6.204852, 6.300065, 6.261086, 6.066943, 
    5.75868, 5.4425, 5.212531, 5.086449, 5.030761, 5.009799, 5.002829, 
    5.000745, 5.000179, 5.000041, 5.000009, 5.000001, 5, 5,
  // momentumY(2,26, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000003, 5.000014, 5.000048, 5.000146, 
    5.00039, 5.000851, 0, 7.33743, 7.027562, 6.586339, 6.171353, 5.805575, 
    5.335398, 4.902407, 4.603593, 4.448595, 4.403919, 4.448415, 4.602663, 
    4.898159, 5.318843, 5.750269, 6.009683, 6.196589, 6.285078, 6.23819, 
    6.038265, 5.73082, 5.422204, 5.201324, 5.08152, 5.028931, 5.009201, 
    5.002654, 5.000698, 5.000167, 5.000037, 5.000008, 5.000001, 5, 5,
  // momentumY(2,27, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5.000003, 5.000013, 5.000049, 5.000171, 5.000519, 
    5.001362, 5.002976, 0, 7.16783, 6.897426, 6.511255, 6.142797, 5.811236, 
    5.40094, 5.024333, 4.753986, 4.602839, 4.55656, 4.602669, 4.753144, 
    5.020627, 5.386737, 5.76387, 6.004327, 6.174033, 6.24164, 6.170797, 
    5.954158, 5.650199, 5.364344, 5.169673, 5.067611, 5.023739, 5.00749, 
    5.002146, 5.000562, 5.000135, 5.00003, 5.000006, 5.000001, 5, 5,
  // momentumY(2,28, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5.000002, 5.00001, 5.000044, 5.000165, 5.000557, 
    5.001666, 5.004333, 5.009483, 0, 6.869401, 6.684888, 6.407736, 6.123141, 
    5.847076, 5.522937, 5.231577, 5.021283, 4.898301, 4.858558, 4.898164, 
    5.020629, 5.228784, 5.51234, 5.811723, 6.019951, 6.153419, 6.174369, 
    6.053992, 5.808561, 5.516597, 5.273223, 5.121716, 5.046975, 5.016093, 
    5.004971, 5.001396, 5.000359, 5.000084, 5.000018, 5.000003, 5, 5, 5,
  // momentumY(2,29, 0-49)
    5, 5, 5, 5, 5, 5, 5.000001, 5.000007, 5.000031, 5.00013, 5.000485, 
    5.001624, 5.004813, 5.012438, 5.027185, 0, 6.458423, 6.39655, 6.269349, 
    6.105521, 5.915573, 5.701647, 5.514119, 5.387164, 5.318938, 5.296925, 
    5.318848, 5.386738, 5.51234, 5.694969, 5.893331, 6.040654, 6.106858, 
    6.056882, 5.88108, 5.622988, 5.367393, 5.181498, 5.076715, 5.028435, 
    5.009418, 5.002819, 5.000768, 5.000192, 5.000044, 5.000009, 5.000001, 5, 
    5, 5,
  // momentumY(2,30, 0-49)
    5, 5, 5, 5, 5, 5, 5.000004, 5.000019, 5.000091, 5.000392, 5.001544, 
    5.005568, 5.018255, 5.053765, 5.13902, 5.339774, 5.824156, 5.992731, 
    6.068674, 6.060568, 5.985876, 5.89627, 5.812539, 5.764076, 5.750317, 
    5.746958, 5.750272, 5.763871, 5.811723, 5.893331, 5.976495, 6.034697, 
    6.008182, 5.878283, 5.663725, 5.425284, 5.229616, 5.105653, 5.042273, 
    5.014987, 5.004771, 5.001375, 5.000361, 5.000087, 5.00002, 5.000003, 5, 
    5, 5, 5,
  // momentumY(2,31, 0-49)
    5, 5, 5, 5, 5, 5, 5.000002, 5.000012, 5.000059, 5.000257, 5.001028, 
    5.003737, 5.01235, 5.036781, 5.097425, 5.235366, 5.544514, 5.750298, 
    5.92068, 6.020491, 6.03864, 6.041875, 6.020286, 6.00441, 6.009703, 
    6.012483, 6.009684, 6.004327, 6.019951, 6.040655, 6.034697, 6.009424, 
    5.894237, 5.699006, 5.470706, 5.269968, 5.132443, 5.056403, 5.021201, 
    5.007127, 5.002162, 5.000596, 5.000149, 5.000036, 5.000008, 5.000001, 5, 
    5, 5, 5,
  // momentumY(2,32, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5.000005, 5.000028, 5.000126, 5.000518, 5.00194, 
    5.006609, 5.020349, 5.056161, 5.140028, 5.324083, 5.513662, 5.720868, 
    5.898491, 6.009674, 6.107315, 6.153543, 6.174064, 6.196596, 6.204853, 
    6.196589, 6.174033, 6.153419, 6.106858, 6.008182, 5.894237, 5.710595, 
    5.493689, 5.295689, 5.152572, 5.068489, 5.02711, 5.009576, 5.003045, 
    5.000876, 5.00023, 5.000055, 5.000013, 5.000002, 5, 5, 5, 5, 5,
  // momentumY(2,33, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000011, 5.000051, 5.000216, 5.000844, 
    5.002991, 5.009605, 5.02779, 5.072512, 5.172647, 5.311225, 5.497193, 
    5.700458, 5.878788, 6.057036, 6.17441, 6.241651, 6.28508, 6.300066, 
    6.285078, 6.241639, 6.174369, 6.056882, 5.878283, 5.699006, 5.493689, 
    5.304491, 5.163324, 5.076609, 5.031737, 5.011728, 5.003897, 5.001171, 
    5.000319, 5.00008, 5.000019, 5.000004, 5, 5, 5, 5, 5, 5,
  // momentumY(2,34, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5.000003, 5.000018, 5.000078, 5.000318, 5.001177, 
    5.003963, 5.012051, 5.033063, 5.082146, 5.165304, 5.29673, 5.471141, 
    5.663877, 5.881125, 6.054005, 6.170801, 6.238191, 6.261086, 6.238191, 
    6.170798, 6.053992, 5.88108, 5.663725, 5.470706, 5.295689, 5.163324, 
    5.079466, 5.034278, 5.013205, 5.004572, 5.00143, 5.000405, 5.000104, 
    5.000025, 5.000005, 5, 5, 5, 5, 5, 5, 5,
  // momentumY(2,35, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000006, 5.000025, 5.000106, 5.000411, 
    5.001449, 5.004638, 5.0134, 5.034968, 5.077124, 5.152843, 5.270081, 
    5.425323, 5.623, 5.808566, 5.954159, 6.038265, 6.066944, 6.038265, 
    5.954159, 5.808562, 5.622989, 5.425284, 5.269968, 5.152572, 5.076609, 
    5.034278, 5.01373, 5.004946, 5.001609, 5.000474, 5.000127, 5.000031, 
    5.000007, 5.000001, 5, 5, 5, 5, 5, 5, 5,
  // momentumY(2,36, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000007, 5.000031, 5.000127, 
    5.000473, 5.001596, 5.004863, 5.013367, 5.031859, 5.068552, 5.132469, 
    5.229624, 5.367395, 5.516597, 5.650199, 5.73082, 5.75868, 5.73082, 
    5.650199, 5.516597, 5.367393, 5.229616, 5.132443, 5.068489, 5.031737, 
    5.013205, 5.004946, 5.001672, 5.000513, 5.000143, 5.000036, 5.000008, 
    5.000001, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumY(2,37, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000009, 5.000036, 5.000139, 
    5.000494, 5.001589, 5.004607, 5.011755, 5.027123, 5.056408, 5.105654, 
    5.181498, 5.273223, 5.364344, 5.422204, 5.4425, 5.422204, 5.364344, 
    5.273223, 5.181498, 5.105653, 5.056403, 5.02711, 5.011728, 5.004572, 
    5.001609, 5.000513, 5.000149, 5.000039, 5.00001, 5.000002, 5, 5, 5, 5, 5, 
    5, 5, 5, 5,
  // momentumY(2,38, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.00001, 5.000037, 5.000138, 
    5.00047, 5.001437, 5.003901, 5.009578, 5.021202, 5.042273, 5.076715, 
    5.121716, 5.169673, 5.201324, 5.212531, 5.201324, 5.169673, 5.121716, 
    5.076715, 5.042273, 5.021201, 5.009576, 5.003897, 5.00143, 5.000474, 
    5.000143, 5.000039, 5.00001, 5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumY(2,39, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.00001, 5.000034, 
    5.000126, 5.000407, 5.001172, 5.003045, 5.007127, 5.014987, 5.028435, 
    5.046975, 5.067611, 5.08152, 5.086449, 5.08152, 5.067611, 5.046975, 
    5.028435, 5.014987, 5.007127, 5.003045, 5.001171, 5.000405, 5.000127, 
    5.000036, 5.00001, 5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumY(2,40, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000008, 5.000031, 
    5.000104, 5.000319, 5.000876, 5.002162, 5.004771, 5.009418, 5.016093, 
    5.023739, 5.028931, 5.030761, 5.028931, 5.023739, 5.016093, 5.009418, 
    5.004771, 5.002162, 5.000876, 5.000319, 5.000104, 5.000031, 5.000008, 
    5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumY(2,41, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000007, 5.000025, 
    5.00008, 5.00023, 5.000596, 5.001375, 5.002819, 5.004971, 5.00749, 
    5.009201, 5.009799, 5.009201, 5.00749, 5.004971, 5.002819, 5.001375, 
    5.000596, 5.00023, 5.00008, 5.000025, 5.000007, 5.000001, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5,
  // momentumY(2,42, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000005, 
    5.000019, 5.000055, 5.000149, 5.000361, 5.000768, 5.001396, 5.002146, 
    5.002654, 5.002829, 5.002654, 5.002146, 5.001396, 5.000768, 5.000361, 
    5.000149, 5.000055, 5.000019, 5.000005, 5.000001, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5,
  // momentumY(2,43, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000004, 5.000013, 
    5.000036, 5.000087, 5.000192, 5.000359, 5.000562, 5.000698, 5.000745, 
    5.000698, 5.000562, 5.000359, 5.000192, 5.000087, 5.000036, 5.000013, 
    5.000004, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumY(2,44, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000008, 
    5.00002, 5.000044, 5.000084, 5.000135, 5.000167, 5.000179, 5.000167, 
    5.000135, 5.000084, 5.000044, 5.00002, 5.000008, 5.000002, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumY(2,45, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 
    5.000003, 5.000009, 5.000018, 5.00003, 5.000037, 5.000041, 5.000037, 
    5.00003, 5.000018, 5.000009, 5.000003, 5.000001, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumY(2,46, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 
    5.000003, 5.000006, 5.000008, 5.000009, 5.000008, 5.000006, 5.000003, 
    5.000001, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumY(2,47, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5.000001, 5.000001, 5.000001, 5.000001, 5.000001, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumY(2,48, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumY(2,49, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5,
  // momentumY(3,0, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 
    5.000003, 5.000006, 5.00001, 5.000014, 5.000018, 5.000019, 5.000018, 
    5.000014, 5.00001, 5.000006, 5.000003, 5.000001, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumY(3,1, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000007, 
    5.000014, 5.000024, 5.000038, 5.000054, 5.000065, 5.000069, 5.000065, 
    5.000054, 5.000038, 5.000024, 5.000014, 5.000007, 5.000002, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumY(3,2, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000005, 
    5.000013, 5.000025, 5.000051, 5.000089, 5.000139, 5.000192, 5.00023, 
    5.000245, 5.00023, 5.000192, 5.000139, 5.000089, 5.000051, 5.000025, 
    5.000013, 5.000005, 5.000001, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumY(3,3, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000003, 5.000008, 5.00002, 
    5.000045, 5.000092, 5.000175, 5.000303, 5.000471, 5.000645, 5.000771, 
    5.000815, 5.000771, 5.000645, 5.000471, 5.000303, 5.000175, 5.000092, 
    5.000045, 5.00002, 5.000008, 5.000003, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5,
  // momentumY(3,4, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000004, 5.000012, 5.00003, 
    5.00007, 5.000153, 5.000309, 5.000576, 5.000975, 5.001488, 5.002019, 
    5.0024, 5.002537, 5.0024, 5.002019, 5.001488, 5.000975, 5.000576, 
    5.000309, 5.000153, 5.00007, 5.00003, 5.000012, 5.000004, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5,
  // momentumY(3,5, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000005, 5.000016, 
    5.000041, 5.000101, 5.000232, 5.000495, 5.000975, 5.001767, 5.002935, 
    5.004404, 5.005916, 5.006993, 5.007383, 5.006993, 5.005916, 5.004404, 
    5.002935, 5.001767, 5.000974, 5.000495, 5.000232, 5.000101, 5.000041, 
    5.000016, 5.000005, 5.000001, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumY(3,6, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000007, 5.00002, 5.000052, 
    5.000135, 5.000328, 5.000727, 5.001502, 5.002871, 5.005065, 5.008235, 
    5.012152, 5.016148, 5.018981, 5.020005, 5.018981, 5.016148, 5.012152, 
    5.008235, 5.005065, 5.00287, 5.001501, 5.000726, 5.000327, 5.000136, 
    5.000052, 5.00002, 5.000007, 5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumY(3,7, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000008, 5.000022, 5.000062, 
    5.000168, 5.000426, 5.000994, 5.002136, 5.004256, 5.007876, 5.013505, 
    5.021459, 5.0311, 5.040833, 5.047673, 5.050141, 5.047673, 5.040833, 
    5.0311, 5.021459, 5.013503, 5.007874, 5.004254, 5.00213, 5.000989, 
    5.000427, 5.000171, 5.000064, 5.000023, 5.000008, 5.000002, 5, 5, 5, 5, 
    5, 5, 5, 5, 5,
  // momentumY(3,8, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000008, 5.000023, 5.000071, 
    5.000197, 5.000516, 5.001256, 5.002826, 5.005837, 5.011214, 5.020035, 
    5.033278, 5.051542, 5.073155, 5.094623, 5.109491, 5.114835, 5.109491, 
    5.094623, 5.073154, 5.05154, 5.033274, 5.020027, 5.011199, 5.005819, 
    5.002808, 5.001259, 5.000525, 5.000204, 5.000074, 5.000025, 5.000008, 
    5.000002, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumY(3,9, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000008, 5.000024, 5.000072, 5.000215, 
    5.000583, 5.001472, 5.003447, 5.007477, 5.01482, 5.027332, 5.046957, 
    5.07516, 5.112832, 5.155911, 5.197577, 5.225729, 5.235758, 5.225728, 
    5.197576, 5.155908, 5.112823, 5.075142, 5.046923, 5.027278, 5.014745, 
    5.00741, 5.003462, 5.001504, 5.000608, 5.000228, 5.00008, 5.000026, 
    5.000009, 5.000002, 5, 5, 5, 5, 5, 5, 5,
  // momentumY(3,10, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000007, 5.000022, 5.000071, 5.000216, 
    5.00061, 5.001602, 5.003899, 5.008797, 5.018371, 5.034782, 5.061243, 
    5.100461, 5.15364, 5.221577, 5.295402, 5.36382, 5.408352, 5.423996, 
    5.408351, 5.363815, 5.29539, 5.221547, 5.153577, 5.100338, 5.061041, 
    5.034512, 5.018124, 5.008841, 5.004006, 5.001688, 5.000662, 5.000242, 
    5.000082, 5.000026, 5.000008, 5.000002, 5, 5, 5, 5, 5, 5,
  // momentumY(3,11, 0-49)
    5, 5, 5, 5, 5, 5, 5.000001, 5.000006, 5.000021, 5.000064, 5.000203, 
    5.000594, 5.001617, 5.004089, 5.009582, 5.020787, 5.04175, 5.075024, 
    5.125049, 5.193873, 5.280046, 5.383638, 5.488432, 5.579867, 5.636599, 
    5.656176, 5.636593, 5.57985, 5.488389, 5.383534, 5.279824, 5.193449, 
    5.124352, 5.074101, 5.040899, 5.020916, 5.009921, 5.004369, 5.001788, 
    5.000681, 5.000242, 5.00008, 5.000025, 5.000008, 5.000002, 5, 5, 5, 5, 5,
  // momentumY(3,12, 0-49)
    5, 5, 5, 5, 5, 5, 5.000005, 5.000017, 5.000055, 5.000177, 5.000535, 
    5.001513, 5.003968, 5.009657, 5.021753, 5.045288, 5.087358, 5.14761, 
    5.230261, 5.333305, 5.449304, 5.57871, 5.698251, 5.795069, 5.852182, 
    5.871558, 5.852166, 5.795019, 5.698119, 5.578391, 5.448622, 5.331985, 
    5.228084, 5.144711, 5.084641, 5.045663, 5.022761, 5.010503, 5.004496, 
    5.001788, 5.000662, 5.000228, 5.000074, 5.000023, 5.000007, 5.000001, 5, 
    5, 5, 5,
  // momentumY(3,13, 0-49)
    5, 5, 5, 5, 5, 5.000002, 5.000013, 5.000043, 5.000142, 5.000446, 
    5.001304, 5.003549, 5.008974, 5.021013, 5.045398, 5.090425, 5.167326, 
    5.262846, 5.378967, 5.506453, 5.631666, 5.760675, 5.867614, 5.947062, 
    5.992007, 6.007091, 5.991964, 5.946927, 5.867256, 5.75981, 5.629799, 
    5.502812, 5.372893, 5.25464, 5.159427, 5.091476, 5.048205, 5.023404, 
    5.010503, 5.004369, 5.001688, 5.000608, 5.000204, 5.000064, 5.00002, 
    5.000005, 5, 5, 5, 5,
  // momentumY(3,14, 0-49)
    5, 5, 5, 5, 5.000001, 5.000009, 5.000031, 5.000105, 5.00034, 5.001029, 
    5.002908, 5.007648, 5.018635, 5.041913, 5.086556, 5.164249, 5.291772, 
    5.421392, 5.55587, 5.681244, 5.783919, 5.882294, 5.952684, 5.99908, 
    6.024866, 6.03354, 6.024758, 5.998743, 5.951796, 5.880162, 5.77933, 
    5.672307, 5.540854, 5.400769, 5.271254, 5.167127, 5.093842, 5.048205, 
    5.022761, 5.009921, 5.004006, 5.001504, 5.000525, 5.000171, 5.000052, 
    5.000016, 5.000004, 5, 5, 5,
  // momentumY(3,15, 0-49)
    5, 5, 5, 5, 5.000005, 5.00002, 5.000069, 5.000233, 5.000735, 5.002163, 
    5.005921, 5.015044, 5.035314, 5.076136, 5.14962, 5.26931, 5.461556, 
    5.608839, 5.731626, 5.821412, 5.873544, 5.920516, 5.942305, 5.950413, 
    5.955587, 5.957473, 5.955333, 5.949632, 5.940266, 5.915689, 5.863268, 
    5.801664, 5.698636, 5.56323, 5.414839, 5.276899, 5.167127, 5.091476, 
    5.045663, 5.020916, 5.00884, 5.003462, 5.001259, 5.000427, 5.000136, 
    5.000041, 5.000012, 5.000003, 5, 5,
  // momentumY(3,16, 0-49)
    5, 5, 5, 5.000002, 5.000011, 5.000041, 5.000143, 5.000468, 5.001436, 
    5.004103, 5.010897, 5.026792, 5.060598, 5.124972, 5.232549, 5.396155, 
    5.662586, 5.799902, 5.878317, 5.906157, 5.892824, 5.879972, 5.850737, 
    5.821409, 5.806584, 5.801819, 5.806024, 5.819709, 5.846377, 5.869823, 
    5.871604, 5.866385, 5.813318, 5.711125, 5.5706, 5.414839, 5.271254, 
    5.159427, 5.084641, 5.040899, 5.018124, 5.00741, 5.002808, 5.000989, 
    5.000327, 5.000101, 5.00003, 5.000008, 5.000001, 5,
  // momentumY(3,17, 0-49)
    5, 5, 5.000001, 5.000005, 5.000021, 5.000075, 5.000259, 5.000828, 
    5.002479, 5.006911, 5.017881, 5.042683, 5.093165, 5.18362, 5.322259, 
    5.521502, 5.866402, 5.969814, 5.983183, 5.936786, 5.854723, 5.780489, 
    5.701207, 5.636169, 5.601222, 5.58957, 5.600065, 5.632699, 5.692458, 
    5.76054, 5.814003, 5.863031, 5.867137, 5.816883, 5.711125, 5.56323, 
    5.400769, 5.25464, 5.144711, 5.0741, 5.034512, 5.014745, 5.005819, 
    5.00213, 5.000726, 5.000232, 5.00007, 5.00002, 5.000005, 5,
  // momentumY(3,18, 0-49)
    5, 5, 5.000002, 5.000009, 5.000031, 5.000117, 5.000395, 5.001246, 
    5.003667, 5.010052, 5.025521, 5.059556, 5.126149, 5.238306, 5.394081, 
    5.615667, 6.035935, 6.101533, 6.04922, 5.929343, 5.78085, 5.644381, 
    5.515065, 5.414158, 5.357251, 5.337825, 5.354997, 5.407474, 5.498516, 
    5.607554, 5.707836, 5.802571, 5.86004, 5.867137, 5.813318, 5.698636, 
    5.540854, 5.372893, 5.228083, 5.124352, 5.061041, 5.027278, 5.011199, 
    5.004254, 5.001501, 5.000495, 5.000153, 5.000045, 5.000013, 5.000002,
  // momentumY(3,19, 0-49)
    5, 5, 5.000002, 5.000011, 5.000038, 5.00014, 5.000471, 5.001475, 
    5.004326, 5.011827, 5.029943, 5.069492, 5.145236, 5.266404, 5.417098, 
    5.657688, 6.133231, 6.183744, 6.085767, 5.90326, 5.691944, 5.490312, 
    5.308599, 5.169163, 5.086947, 5.058302, 5.082806, 5.156998, 5.279012, 
    5.426208, 5.569045, 5.70021, 5.80257, 5.863031, 5.866385, 5.801664, 
    5.672307, 5.502812, 5.331985, 5.193449, 5.100338, 5.046923, 5.020027, 
    5.007874, 5.00287, 5.000974, 5.000309, 5.000092, 5.000025, 5.000007,
  // momentumY(3,20, 0-49)
    5, 5, 5.000001, 5.000006, 5.000022, 5.000076, 5.000246, 5.000745, 
    5.002099, 5.005454, 5.012992, 5.028082, 5.054316, 5.092286, 5.134862, 0, 
    6.537839, 6.444597, 6.224334, 5.931908, 5.627497, 5.341224, 5.09673, 
    4.91181, 4.799217, 4.759322, 4.791854, 4.890079, 5.043821, 5.226887, 
    5.408791, 5.569041, 5.707834, 5.814003, 5.871604, 5.863268, 5.779329, 
    5.629799, 5.448622, 5.279824, 5.153577, 5.075142, 5.033274, 5.013503, 
    5.005065, 5.001767, 5.000576, 5.000175, 5.000051, 5.000014,
  // momentumY(3,21, 0-49)
    5, 5, 5, 5.000002, 5.000011, 5.000037, 5.000119, 5.000364, 5.001029, 
    5.002694, 5.006472, 5.01416, 5.027897, 5.048741, 5.073972, 0, 6.715348, 
    6.582877, 6.306049, 5.934135, 5.539999, 5.157746, 4.834559, 4.587932, 
    4.433352, 4.378251, 4.422956, 4.55676, 4.757838, 4.992012, 5.226871, 
    5.426194, 5.607547, 5.760535, 5.869822, 5.915688, 5.880161, 5.75981, 
    5.578391, 5.383534, 5.221547, 5.112823, 5.05154, 5.021459, 5.008235, 
    5.002935, 5.000975, 5.000303, 5.000089, 5.000024,
  // momentumY(3,22, 0-49)
    5, 5, 5, 5, 5.000004, 5.000016, 5.000052, 5.00016, 5.000462, 5.001224, 
    5.002986, 5.006641, 5.013321, 5.023751, 5.036767, 0, 6.819324, 6.665093, 
    6.350619, 5.917248, 5.445622, 4.973551, 4.571023, 4.255342, 4.050066, 
    3.976002, 4.036703, 4.214768, 4.470624, 4.757758, 5.043741, 5.278961, 
    5.498487, 5.692443, 5.846371, 5.940264, 5.951795, 5.867255, 5.69812, 
    5.488389, 5.29539, 5.155908, 5.073154, 5.0311, 5.012152, 5.004404, 
    5.001488, 5.000471, 5.000139, 5.000038,
  // momentumY(3,23, 0-49)
    5, 5, 5, 5, 5.000001, 5.000007, 5.000022, 5.00007, 5.000204, 5.000552, 
    5.001373, 5.003109, 5.006342, 5.011469, 5.017878, 0, 6.881858, 6.715767, 
    6.377157, 5.89924, 5.365091, 4.814788, 4.335211, 3.944315, 3.680533, 
    3.584269, 3.664799, 3.895799, 4.214448, 4.556406, 4.88979, 5.156824, 
    5.407378, 5.63265, 5.819686, 5.949622, 5.99874, 5.946925, 5.795018, 
    5.57985, 5.363815, 5.197576, 5.094623, 5.040833, 5.016148, 5.005916, 
    5.002019, 5.000645, 5.000192, 5.000054,
  // momentumY(3,24, 0-49)
    5, 5, 5, 5, 5, 5.000004, 5.000014, 5.000044, 5.000131, 5.000354, 
    5.000885, 5.002009, 5.004103, 5.00741, 5.011444, 0, 6.913795, 6.743283, 
    6.393038, 5.88919, 5.313772, 4.708361, 4.169513, 3.717096, 3.405324, 
    3.291309, 3.388295, 3.663615, 4.035308, 4.421719, 4.790909, 5.082253, 
    5.354696, 5.599913, 5.805953, 5.955301, 6.024744, 5.991959, 5.852164, 
    5.636593, 5.40835, 5.225728, 5.109491, 5.047673, 5.018981, 5.006993, 
    5.0024, 5.000771, 5.00023, 5.000065,
  // momentumY(3,25, 0-49)
    5, 5, 5, 5, 5.000001, 5.000007, 5.000023, 5.000068, 5.000196, 5.000519, 
    5.001256, 5.00277, 5.005505, 5.009689, 5.014659, 0, 6.917509, 6.746934, 
    6.394336, 5.883124, 5.294426, 4.670211, 4.109842, 3.634244, 3.304592, 
    3.184185, 3.287201, 3.579186, 3.97121, 4.374317, 4.756428, 5.056643, 
    5.336924, 5.589113, 5.801601, 5.957374, 6.033497, 6.007074, 5.871552, 
    5.656174, 5.423996, 5.235758, 5.114835, 5.050141, 5.020005, 5.007383, 
    5.002537, 5.000815, 5.000245, 5.000069,
  // momentumY(3,26, 0-49)
    5, 5, 5, 5, 5.000005, 5.000018, 5.000054, 5.000162, 5.000451, 5.001157, 
    5.00272, 5.005827, 5.011258, 5.019319, 5.028754, 0, 6.889607, 6.723534, 
    6.378369, 5.879577, 5.308405, 4.705863, 4.168527, 3.716762, 3.405225, 
    3.291283, 3.388287, 3.663613, 4.035307, 4.421719, 4.790908, 5.082252, 
    5.354695, 5.599913, 5.805953, 5.955301, 6.024744, 5.991959, 5.852164, 
    5.636593, 5.40835, 5.225728, 5.109491, 5.047673, 5.018981, 5.006993, 
    5.0024, 5.000771, 5.00023, 5.000065,
  // momentumY(3,27, 0-49)
    5, 5, 5, 5.000003, 5.000013, 5.000042, 5.000131, 5.000385, 5.001048, 
    5.002628, 5.006048, 5.012661, 5.02387, 5.039977, 5.058367, 0, 6.826754, 
    6.670672, 6.343395, 5.876875, 5.352436, 4.808751, 4.332749, 3.943442, 
    3.680258, 3.58419, 3.664778, 3.895793, 4.214446, 4.556406, 4.889789, 
    5.156823, 5.407378, 5.63265, 5.819686, 5.949621, 5.99874, 5.946925, 
    5.795018, 5.57985, 5.363815, 5.197576, 5.094623, 5.040833, 5.016148, 
    5.005916, 5.002019, 5.000645, 5.000192, 5.000054,
  // momentumY(3,28, 0-49)
    5, 5, 5.000001, 5.000009, 5.000028, 5.000093, 5.000291, 5.000842, 
    5.002254, 5.005562, 5.012565, 5.025754, 5.047345, 5.076943, 5.108829, 0, 
    6.720564, 6.584433, 6.289873, 5.876649, 5.422355, 4.96215, 4.566208, 
    4.253551, 4.049467, 3.975818, 4.036649, 4.214753, 4.470621, 4.757757, 
    5.04374, 5.27896, 5.498487, 5.692443, 5.846371, 5.940264, 5.951794, 
    5.867256, 5.69812, 5.488389, 5.29539, 5.155908, 5.073154, 5.0311, 
    5.012152, 5.004404, 5.001488, 5.000471, 5.000139, 5.000038,
  // momentumY(3,29, 0-49)
    5, 5, 5.000004, 5.000016, 5.000057, 5.000186, 5.000579, 5.001659, 
    5.004405, 5.010764, 5.024003, 5.048273, 5.086257, 5.134563, 5.180684, 0, 
    6.556565, 6.454806, 6.209808, 5.869759, 5.502885, 5.139183, 4.826483, 
    4.584808, 4.432256, 4.377896, 4.422847, 4.556728, 4.757828, 4.99201, 
    5.226871, 5.426193, 5.607547, 5.760535, 5.869822, 5.915688, 5.880161, 
    5.75981, 5.578391, 5.383534, 5.221547, 5.112823, 5.05154, 5.021459, 
    5.008235, 5.002935, 5.000975, 5.000303, 5.000089, 5.000024,
  // momentumY(3,30, 0-49)
    5, 5.000002, 5.000008, 5.000027, 5.0001, 5.000338, 5.001072, 5.003178, 
    5.008781, 5.022519, 5.053143, 5.113769, 5.216212, 5.355342, 5.494076, 
    5.709598, 6.125762, 6.156536, 6.034242, 5.81732, 5.566053, 5.311934, 
    5.084235, 4.906974, 4.7975, 4.758753, 4.791675, 4.890025, 5.043805, 
    5.226883, 5.40879, 5.569041, 5.707834, 5.814003, 5.871604, 5.863268, 
    5.779329, 5.629799, 5.448622, 5.279824, 5.153577, 5.075142, 5.033274, 
    5.013503, 5.005065, 5.001767, 5.000576, 5.000175, 5.000051, 5.000014,
  // momentumY(3,31, 0-49)
    5, 5.000001, 5.000006, 5.000023, 5.000086, 5.000294, 5.000936, 5.002785, 
    5.007725, 5.019886, 5.047167, 5.101953, 5.197631, 5.337241, 5.499212, 
    5.707389, 6.101362, 6.130861, 6.032712, 5.862597, 5.666519, 5.477023, 
    5.3025, 5.166655, 5.086007, 5.057975, 5.082697, 5.156963, 5.279002, 
    5.426205, 5.569045, 5.70021, 5.80257, 5.863031, 5.866385, 5.801664, 
    5.672307, 5.502812, 5.331985, 5.193449, 5.100338, 5.046923, 5.020027, 
    5.007874, 5.00287, 5.000974, 5.000309, 5.000092, 5.000025, 5.000007,
  // momentumY(3,32, 0-49)
    5, 5, 5.000003, 5.000016, 5.000057, 5.000198, 5.000641, 5.001941, 
    5.005484, 5.014384, 5.034873, 5.077482, 5.155878, 5.27987, 5.442998, 
    5.649105, 5.993998, 6.054826, 6.009722, 5.902009, 5.764829, 5.636314, 
    5.511456, 5.412694, 5.356704, 5.337633, 5.354934, 5.407454, 5.49851, 
    5.607553, 5.707836, 5.802571, 5.86004, 5.867137, 5.813318, 5.698636, 
    5.540854, 5.372893, 5.228083, 5.124352, 5.061041, 5.027278, 5.011199, 
    5.004254, 5.001501, 5.000495, 5.000153, 5.000045, 5.000013, 5.000002,
  // momentumY(3,33, 0-49)
    5, 5, 5.000001, 5.000009, 5.000031, 5.000113, 5.000374, 5.00116, 
    5.003356, 5.009038, 5.022561, 5.051877, 5.108922, 5.206487, 5.349631, 
    5.540675, 5.829793, 5.934906, 5.95664, 5.919773, 5.845279, 5.775891, 
    5.699202, 5.635369, 5.600927, 5.589468, 5.600031, 5.632689, 5.692454, 
    5.760539, 5.814003, 5.863031, 5.867137, 5.816883, 5.711125, 5.563231, 
    5.400769, 5.25464, 5.144711, 5.0741, 5.034512, 5.014745, 5.005819, 
    5.00213, 5.000726, 5.000232, 5.00007, 5.00002, 5.000005, 5,
  // momentumY(3,34, 0-49)
    5, 5, 5, 5.000003, 5.000016, 5.000058, 5.000192, 5.000611, 5.001822, 
    5.00506, 5.013054, 5.031149, 5.068315, 5.13659, 5.246739, 5.405913, 
    5.637955, 5.777564, 5.862308, 5.896429, 5.887648, 5.877523, 5.849693, 
    5.821001, 5.806437, 5.801769, 5.806009, 5.819705, 5.846376, 5.869823, 
    5.871605, 5.866385, 5.813318, 5.711125, 5.5706, 5.414839, 5.271254, 
    5.159427, 5.084641, 5.040899, 5.018124, 5.00741, 5.002808, 5.000989, 
    5.000327, 5.000101, 5.00003, 5.000008, 5.000001, 5,
  // momentumY(3,35, 0-49)
    5, 5, 5, 5.000001, 5.000007, 5.000026, 5.000089, 5.00029, 5.000893, 
    5.002561, 5.006839, 5.016948, 5.038792, 5.081545, 5.156356, 5.273779, 
    5.448004, 5.596495, 5.722991, 5.816328, 5.870923, 5.919303, 5.941797, 
    5.950219, 5.955517, 5.957448, 5.955325, 5.949628, 5.940266, 5.915689, 
    5.863268, 5.801664, 5.698636, 5.56323, 5.414839, 5.276899, 5.167127, 
    5.091476, 5.045663, 5.020916, 5.00884, 5.003462, 5.001259, 5.000427, 
    5.000136, 5.000041, 5.000012, 5.000003, 5, 5,
  // momentumY(3,36, 0-49)
    5, 5, 5, 5, 5.000002, 5.000011, 5.000038, 5.000125, 5.000399, 5.001182, 
    5.00327, 5.008418, 5.020082, 5.044224, 5.089479, 5.166116, 5.285483, 
    5.41548, 5.55173, 5.678836, 5.782701, 5.881738, 5.952456, 5.998994, 
    6.024836, 6.033529, 6.024755, 5.998743, 5.951795, 5.880162, 5.77933, 
    5.672307, 5.540854, 5.400769, 5.271254, 5.167127, 5.093842, 5.048205, 
    5.022761, 5.009921, 5.004006, 5.001504, 5.000525, 5.000171, 5.000052, 
    5.000016, 5.000004, 5, 5, 5,
  // momentumY(3,37, 0-49)
    5, 5, 5, 5, 5, 5.000004, 5.000015, 5.000051, 5.000163, 5.000501, 
    5.001435, 5.003837, 5.00953, 5.021924, 5.046564, 5.091146, 5.164802, 
    5.260377, 5.377213, 5.50543, 5.631152, 5.760442, 5.867519, 5.947026, 
    5.991995, 6.007086, 5.991962, 5.946927, 5.867255, 5.75981, 5.629799, 
    5.502812, 5.372893, 5.25464, 5.159427, 5.091476, 5.048205, 5.023404, 
    5.010503, 5.004369, 5.001688, 5.000608, 5.000204, 5.000064, 5.00002, 
    5.000005, 5, 5, 5, 5,
  // momentumY(3,38, 0-49)
    5, 5, 5, 5, 5, 5, 5.000005, 5.00002, 5.000062, 5.000195, 5.00058, 
    5.001613, 5.004166, 5.009988, 5.022183, 5.045549, 5.086459, 5.146701, 
    5.229607, 5.33292, 5.449109, 5.578621, 5.698215, 5.795055, 5.852177, 
    5.871556, 5.852166, 5.79502, 5.69812, 5.578392, 5.448622, 5.331985, 
    5.228083, 5.144711, 5.084641, 5.045663, 5.022761, 5.010503, 5.004496, 
    5.001788, 5.000662, 5.000228, 5.000074, 5.000023, 5.000007, 5.000001, 5, 
    5, 5, 5,
  // momentumY(3,39, 0-49)
    5, 5, 5, 5, 5, 5, 5.000001, 5.000007, 5.000022, 5.000071, 5.000218, 
    5.000627, 5.001684, 5.004201, 5.00973, 5.020876, 5.04146, 5.074723, 
    5.124831, 5.193744, 5.27998, 5.383608, 5.48842, 5.579863, 5.636596, 
    5.656175, 5.636593, 5.57985, 5.488389, 5.383535, 5.279824, 5.193449, 
    5.124352, 5.0741, 5.040899, 5.020916, 5.009921, 5.004369, 5.001788, 
    5.000681, 5.000242, 5.00008, 5.000025, 5.000008, 5.000002, 5, 5, 5, 5, 5,
  // momentumY(3,40, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000008, 5.000024, 5.000075, 5.000226, 
    5.00063, 5.001637, 5.003948, 5.008826, 5.018284, 5.034691, 5.061178, 
    5.100423, 5.153621, 5.221567, 5.295398, 5.363819, 5.408352, 5.423996, 
    5.408351, 5.363815, 5.29539, 5.221547, 5.153577, 5.100338, 5.061041, 
    5.034512, 5.018124, 5.00884, 5.004006, 5.001688, 5.000662, 5.000242, 
    5.000082, 5.000026, 5.000008, 5.000002, 5, 5, 5, 5, 5, 5,
  // momentumY(3,41, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000008, 5.000024, 5.000076, 5.00022, 
    5.000594, 5.001486, 5.003456, 5.007452, 5.014793, 5.027314, 5.046945, 
    5.075154, 5.112829, 5.15591, 5.197577, 5.225729, 5.235758, 5.225728, 
    5.197576, 5.155908, 5.112823, 5.075142, 5.046923, 5.027278, 5.014745, 
    5.00741, 5.003462, 5.001504, 5.000608, 5.000228, 5.00008, 5.000026, 
    5.000009, 5.000002, 5, 5, 5, 5, 5, 5, 5,
  // momentumY(3,42, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000008, 5.000024, 5.000072, 
    5.0002, 5.000521, 5.001258, 5.002819, 5.00583, 5.011209, 5.020034, 
    5.033277, 5.051541, 5.073155, 5.094623, 5.109491, 5.114835, 5.109491, 
    5.094623, 5.073154, 5.05154, 5.033274, 5.020027, 5.011199, 5.005819, 
    5.002808, 5.001259, 5.000525, 5.000204, 5.000074, 5.000025, 5.000008, 
    5.000002, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumY(3,43, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000008, 5.000023, 5.000063, 
    5.00017, 5.000428, 5.000993, 5.002134, 5.004256, 5.007876, 5.013503, 
    5.021459, 5.0311, 5.040833, 5.047673, 5.050141, 5.047673, 5.040833, 
    5.0311, 5.021459, 5.013503, 5.007874, 5.004254, 5.00213, 5.000989, 
    5.000427, 5.000171, 5.000064, 5.000023, 5.000008, 5.000002, 5, 5, 5, 5, 
    5, 5, 5, 5, 5,
  // momentumY(3,44, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000007, 5.00002, 5.000052, 
    5.000136, 5.000328, 5.000727, 5.001502, 5.002871, 5.005065, 5.008235, 
    5.012152, 5.016148, 5.018981, 5.020005, 5.018981, 5.016148, 5.012152, 
    5.008235, 5.005065, 5.00287, 5.001501, 5.000726, 5.000327, 5.000136, 
    5.000052, 5.00002, 5.000007, 5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumY(3,45, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000005, 5.000016, 
    5.000041, 5.000101, 5.000232, 5.000495, 5.000975, 5.001767, 5.002935, 
    5.004404, 5.005916, 5.006993, 5.007383, 5.006993, 5.005916, 5.004404, 
    5.002935, 5.001767, 5.000974, 5.000495, 5.000232, 5.000101, 5.000041, 
    5.000016, 5.000005, 5.000001, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumY(3,46, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000004, 5.000012, 5.00003, 
    5.00007, 5.000153, 5.000309, 5.000576, 5.000975, 5.001488, 5.002019, 
    5.0024, 5.002537, 5.0024, 5.002019, 5.001488, 5.000975, 5.000576, 
    5.000309, 5.000153, 5.00007, 5.00003, 5.000012, 5.000004, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5,
  // momentumY(3,47, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000003, 5.000008, 5.00002, 
    5.000045, 5.000092, 5.000175, 5.000303, 5.000471, 5.000645, 5.000771, 
    5.000815, 5.000771, 5.000645, 5.000471, 5.000303, 5.000175, 5.000092, 
    5.000045, 5.00002, 5.000008, 5.000003, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5,
  // momentumY(3,48, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000005, 
    5.000013, 5.000025, 5.000051, 5.000089, 5.000139, 5.000192, 5.000231, 
    5.000245, 5.000231, 5.000192, 5.000139, 5.000089, 5.000051, 5.000025, 
    5.000013, 5.000005, 5.000001, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumY(3,49, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000006, 
    5.000012, 5.000023, 5.000038, 5.000055, 5.000067, 5.000071, 5.000067, 
    5.000055, 5.000038, 5.000023, 5.000012, 5.000006, 5.000002, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumY(4,0, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000006, 5.000013, 
    5.000028, 5.000057, 5.000112, 5.000206, 5.000354, 5.000569, 5.00085, 
    5.001171, 5.001479, 5.001697, 5.001776, 5.001697, 5.001479, 5.001171, 
    5.00085, 5.000569, 5.000354, 5.000206, 5.000112, 5.000057, 5.000028, 
    5.000013, 5.000006, 5.000001, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumY(4,1, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000003, 5.000008, 5.000018, 5.000039, 
    5.000082, 5.000166, 5.000319, 5.000575, 5.000974, 5.001544, 5.002285, 
    5.003127, 5.003933, 5.004504, 5.00471, 5.004504, 5.003933, 5.003127, 
    5.002285, 5.001544, 5.000974, 5.000575, 5.000319, 5.000166, 5.000082, 
    5.000038, 5.000018, 5.000008, 5.000003, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumY(4,2, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000004, 5.00001, 5.000022, 5.00005, 
    5.000111, 5.000235, 5.000467, 5.000876, 5.001545, 5.002564, 5.003994, 
    5.005826, 5.00789, 5.009855, 5.011244, 5.011746, 5.011244, 5.009855, 
    5.00789, 5.005825, 5.003993, 5.002563, 5.001543, 5.000874, 5.000466, 
    5.000235, 5.000111, 5.00005, 5.000022, 5.00001, 5.000004, 5, 5, 5, 5, 5, 
    5, 5, 5, 5,
  // momentumY(4,3, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000005, 5.000011, 5.000026, 5.000062, 
    5.000142, 5.000312, 5.000645, 5.001252, 5.002286, 5.003933, 5.006382, 
    5.00975, 5.014007, 5.018755, 5.023253, 5.026416, 5.027557, 5.026416, 
    5.023252, 5.018755, 5.014006, 5.009748, 5.006378, 5.003928, 5.002279, 
    5.001247, 5.000645, 5.000314, 5.000144, 5.000063, 5.000027, 5.000011, 
    5.000005, 5.000001, 5, 5, 5, 5, 5, 5, 5,
  // momentumY(4,4, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000005, 5.000012, 5.00003, 5.000073, 
    5.000174, 5.000391, 5.000835, 5.001678, 5.003172, 5.005635, 5.009448, 
    5.014966, 5.022386, 5.031617, 5.041789, 5.051358, 5.058033, 5.060435, 
    5.058033, 5.051356, 5.041786, 5.031611, 5.022377, 5.014951, 5.009429, 
    5.005613, 5.003155, 5.001675, 5.00084, 5.000397, 5.000178, 5.000076, 
    5.000031, 5.000013, 5.000005, 5.000001, 5, 5, 5, 5, 5, 5,
  // momentumY(4,5, 0-49)
    5, 5, 5, 5, 5, 5, 5.000002, 5.000006, 5.000013, 5.000031, 5.000082, 
    5.0002, 5.000464, 5.00102, 5.002115, 5.004128, 5.00759, 5.013093, 
    5.021336, 5.032907, 5.048047, 5.066521, 5.086531, 5.105149, 5.117974, 
    5.122565, 5.117973, 5.105145, 5.086521, 5.066501, 5.048014, 5.032856, 
    5.021269, 5.01302, 5.007533, 5.004119, 5.002128, 5.001039, 5.00048, 
    5.00021, 5.000087, 5.000034, 5.000014, 5.000006, 5.000002, 5, 5, 5, 5, 5,
  // momentumY(4,6, 0-49)
    5, 5, 5, 5, 5, 5.000001, 5.000006, 5.000013, 5.000033, 5.000086, 
    5.000218, 5.00052, 5.001176, 5.002513, 5.005054, 5.009583, 5.017104, 
    5.028571, 5.04509, 5.06742, 5.095617, 5.129127, 5.164507, 5.196824, 
    5.218638, 5.226384, 5.218632, 5.196807, 5.164472, 5.12906, 5.095507, 
    5.067253, 5.04487, 5.028332, 5.016919, 5.009551, 5.005095, 5.002568, 
    5.001224, 5.00055, 5.000236, 5.000094, 5.000036, 5.000015, 5.000007, 
    5.000002, 5, 5, 5, 5,
  // momentumY(4,7, 0-49)
    5, 5, 5, 5, 5, 5.000005, 5.000013, 5.000032, 5.000086, 5.000224, 
    5.000552, 5.001284, 5.002817, 5.005834, 5.011383, 5.020915, 5.036179, 
    5.058282, 5.0886, 5.12762, 5.174555, 5.228317, 5.28298, 5.331494, 
    5.363276, 5.374424, 5.363256, 5.331442, 5.282871, 5.228115, 5.174216, 
    5.12711, 5.08793, 5.057558, 5.035612, 5.020813, 5.011489, 5.00599, 
    5.002948, 5.001372, 5.000603, 5.00025, 5.000099, 5.000037, 5.000015, 
    5.000006, 5.000001, 5, 5, 5,
  // momentumY(4,8, 0-49)
    5, 5, 5, 5, 5.000004, 5.000011, 5.00003, 5.000083, 5.000219, 5.000553, 
    5.001321, 5.002983, 5.00635, 5.012745, 5.024074, 5.042771, 5.071508, 
    5.110453, 5.160557, 5.220954, 5.288945, 5.363122, 5.434719, 5.495795, 
    5.534249, 5.547521, 5.534192, 5.49565, 5.434417, 5.36256, 5.288007, 
    5.219527, 5.158675, 5.108407, 5.069887, 5.04248, 5.024346, 5.013159, 
    5.006711, 5.003231, 5.001469, 5.000631, 5.000257, 5.000099, 5.000036, 
    5.000014, 5.000005, 5.000001, 5, 5,
  // momentumY(4,9, 0-49)
    5, 5, 5, 5.000003, 5.00001, 5.000027, 5.000073, 5.000201, 5.000522, 
    5.001283, 5.002978, 5.006522, 5.013456, 5.026117, 5.047627, 5.081541, 
    5.131313, 5.193063, 5.26604, 5.346703, 5.429886, 5.515448, 5.592755, 
    5.65555, 5.693194, 5.705945, 5.693052, 5.655185, 5.592003, 5.51405, 
    5.427536, 5.343099, 5.261235, 5.187773, 5.12704, 5.0808, 5.048308, 
    5.027168, 5.014386, 5.00718, 5.00338, 5.001504, 5.000631, 5.00025, 
    5.000094, 5.000034, 5.000013, 5.000005, 5, 5,
  // momentumY(4,10, 0-49)
    5, 5, 5.000001, 5.000008, 5.000023, 5.000062, 5.000174, 5.000464, 
    5.001174, 5.002803, 5.006311, 5.01339, 5.026711, 5.050013, 5.087704, 
    5.143996, 5.222599, 5.309128, 5.400571, 5.490787, 5.573659, 5.653591, 
    5.720015, 5.770827, 5.799431, 5.808886, 5.799106, 5.770001, 5.718316, 
    5.65044, 5.568353, 5.482604, 5.389545, 5.296785, 5.212377, 5.142366, 
    5.089346, 5.052536, 5.028989, 5.015037, 5.007341, 5.00338, 5.001469, 
    5.000603, 5.000236, 5.000087, 5.000031, 5.000011, 5.000004, 5,
  // momentumY(4,11, 0-49)
    5, 5.000001, 5.000006, 5.000018, 5.000051, 5.000142, 5.000389, 5.00101, 
    5.002481, 5.005745, 5.012537, 5.025723, 5.049498, 5.089058, 5.149407, 
    5.233919, 5.346392, 5.451672, 5.547588, 5.628493, 5.690985, 5.747229, 
    5.788034, 5.816257, 5.830287, 5.834641, 5.829595, 5.814518, 5.784492, 
    5.740716, 5.680092, 5.611754, 5.524933, 5.425946, 5.324495, 5.230956, 
    5.153233, 5.094786, 5.05476, 5.029618, 5.015037, 5.00718, 5.003231, 
    5.001372, 5.00055, 5.00021, 5.000076, 5.000027, 5.00001, 5.000003,
  // momentumY(4,12, 0-49)
    5, 5.000003, 5.000013, 5.000038, 5.000109, 5.000305, 5.000814, 5.002055, 
    5.004901, 5.011015, 5.023273, 5.046094, 5.08526, 5.146695, 5.233996, 
    5.347453, 5.493467, 5.603019, 5.683767, 5.735504, 5.761001, 5.781113, 
    5.78789, 5.788424, 5.785759, 5.784305, 5.784378, 5.784986, 5.780982, 
    5.768596, 5.740397, 5.704315, 5.641876, 5.555245, 5.451858, 5.343374, 
    5.242486, 5.158862, 5.096653, 5.05476, 5.028989, 5.014386, 5.006711, 
    5.002948, 5.001224, 5.00048, 5.000178, 5.000063, 5.000022, 5.000008,
  // momentumY(4,13, 0-49)
    5.000001, 5.000009, 5.000026, 5.000077, 5.000224, 5.000611, 5.001587, 
    5.003901, 5.009038, 5.019696, 5.040237, 5.07673, 5.135884, 5.222372, 
    5.33526, 5.470407, 5.644621, 5.740721, 5.789155, 5.798397, 5.778439, 
    5.757261, 5.727443, 5.699325, 5.679906, 5.672492, 5.677281, 5.692876, 
    5.71471, 5.734662, 5.742108, 5.744841, 5.718772, 5.661288, 5.574646, 
    5.467301, 5.352917, 5.246391, 5.158862, 5.094786, 5.052536, 5.027167, 
    5.013159, 5.00599, 5.002568, 5.001039, 5.000397, 5.000144, 5.00005, 
    5.000018,
  // momentumY(4,14, 0-49)
    5.000004, 5.000016, 5.000051, 5.00015, 5.000423, 5.001134, 5.002876, 
    5.006879, 5.015491, 5.032723, 5.064547, 5.118182, 5.199555, 5.309104, 
    5.438466, 5.581018, 5.776528, 5.845946, 5.853991, 5.817026, 5.75099, 
    5.688416, 5.622475, 5.56643, 5.530651, 5.517122, 5.525881, 5.554883, 
    5.600159, 5.649828, 5.690797, 5.731436, 5.745387, 5.726641, 5.672071, 
    5.58408, 5.472425, 5.352917, 5.242486, 5.153233, 5.089346, 5.048308, 
    5.024346, 5.011489, 5.005095, 5.002128, 5.00084, 5.000314, 5.000111, 
    5.000039,
  // momentumY(4,15, 0-49)
    5.000009, 5.00003, 5.000093, 5.000268, 5.000741, 5.001943, 5.004808, 
    5.011213, 5.02456, 5.050291, 5.095673, 5.167803, 5.269303, 5.393564, 
    5.523967, 5.657652, 5.868953, 5.907986, 5.878179, 5.799743, 5.692262, 
    5.590435, 5.489555, 5.406311, 5.354075, 5.333925, 5.345757, 5.386508, 
    5.452232, 5.527853, 5.598085, 5.67159, 5.722934, 5.744675, 5.730055, 
    5.67552, 5.58408, 5.467301, 5.343374, 5.230956, 5.142365, 5.080799, 
    5.04248, 5.020813, 5.009551, 5.004119, 5.001675, 5.000645, 5.000236, 
    5.000084,
  // momentumY(4,16, 0-49)
    5.000016, 5.000051, 5.000154, 5.000436, 5.001185, 5.003041, 5.007361, 
    5.016769, 5.035784, 5.071095, 5.130445, 5.218989, 5.333667, 5.459665, 
    5.573878, 5.686548, 5.908281, 5.92311, 5.866307, 5.756901, 5.615705, 
    5.477578, 5.342819, 5.232497, 5.162915, 5.135132, 5.148944, 5.199866, 
    5.28306, 5.380913, 5.476108, 5.57633, 5.659531, 5.718256, 5.744269, 
    5.730054, 5.672071, 5.574646, 5.451857, 5.324495, 5.212377, 5.12704, 
    5.069887, 5.035612, 5.016918, 5.007533, 5.003155, 5.001247, 5.000467, 
    5.000169,
  // momentumY(4,17, 0-49)
    5.000024, 5.000076, 5.000226, 5.000637, 5.0017, 5.004287, 5.01019, 
    5.022752, 5.047452, 5.091729, 5.162721, 5.26203, 5.379788, 5.493896, 
    5.577772, 5.66574, 5.886785, 5.890759, 5.822771, 5.696401, 5.531397, 
    5.360797, 5.193435, 5.055688, 4.967145, 4.93014, 4.944488, 5.003893, 
    5.101617, 5.218238, 5.334838, 5.456188, 5.56532, 5.655404, 5.718253, 
    5.744672, 5.726639, 5.661288, 5.555245, 5.425946, 5.296785, 5.187774, 
    5.108407, 5.057558, 5.028332, 5.01302, 5.005613, 5.00228, 5.000876, 
    5.000325,
  // momentumY(4,18, 0-49)
    5.000031, 5.000098, 5.00029, 5.000809, 5.002132, 5.005311, 5.012467, 
    5.027443, 5.05629, 5.106589, 5.184099, 5.286392, 5.397364, 5.489583, 
    5.535452, 5.605662, 5.800894, 5.810308, 5.749249, 5.622153, 5.445377, 
    5.247847, 5.050285, 4.884759, 4.775092, 4.726635, 4.739514, 4.805339, 
    4.914531, 5.046517, 5.181646, 5.319603, 5.449533, 5.565309, 5.659521, 
    5.722928, 5.745382, 5.718771, 5.641876, 5.524933, 5.389545, 5.261234, 
    5.158674, 5.08793, 5.04487, 5.021269, 5.009429, 5.003929, 5.001545, 
    5.000584,
  // momentumY(4,19, 0-49)
    5.000033, 5.000104, 5.000303, 5.000842, 5.002212, 5.00549, 5.012845, 
    5.02818, 5.057574, 5.108389, 5.185361, 5.283393, 5.381967, 5.449668, 
    5.45941, 5.528225, 5.651516, 5.679839, 5.644249, 5.534561, 5.360603, 
    5.14432, 4.920958, 4.727758, 4.594412, 4.531527, 4.540184, 4.609795, 
    4.727152, 4.870959, 5.022038, 5.172999, 5.319552, 5.45614, 5.576295, 
    5.67157, 5.731426, 5.744835, 5.704313, 5.611754, 5.482604, 5.343098, 
    5.219526, 5.12711, 5.067253, 5.032856, 5.014951, 5.00638, 5.002567, 
    5.000986,
  // momentumY(4,20, 0-49)
    5.000022, 5.000071, 5.000206, 5.000566, 5.001461, 5.003547, 5.008075, 
    5.017149, 5.033758, 5.061057, 5.100434, 5.148736, 5.196876, 5.232886, 
    5.249486, 0, 5.72522, 5.722096, 5.663104, 5.536474, 5.342846, 5.092929, 
    4.832631, 4.601823, 4.436234, 4.352537, 4.352442, 4.422397, 4.544476, 
    4.696456, 4.860911, 5.021814, 5.181428, 5.334681, 5.476007, 5.598027, 
    5.690766, 5.742093, 5.74039, 5.680089, 5.568351, 5.427535, 5.288007, 
    5.174216, 5.095507, 5.048014, 5.022378, 5.00975, 5.003997, 5.001556,
  // momentumY(4,21, 0-49)
    5.000014, 5.000044, 5.000126, 5.000348, 5.000903, 5.002204, 5.005051, 
    5.010816, 5.021541, 5.039646, 5.06693, 5.102845, 5.142964, 5.179457, 
    5.204838, 0, 5.693264, 5.683771, 5.624491, 5.49779, 5.296422, 5.020554, 
    4.725423, 4.45422, 4.252345, 4.146114, 4.139155, 4.214416, 4.347202, 
    4.512626, 4.695527, 4.870046, 5.045835, 5.217789, 5.380641, 5.527698, 
    5.649745, 5.734621, 5.768576, 5.740706, 5.650436, 5.514049, 5.36256, 
    5.228116, 5.12906, 5.066501, 5.031611, 5.014006, 5.005826, 5.002292,
  // momentumY(4,22, 0-49)
    5.000008, 5.000024, 5.000072, 5.000199, 5.000521, 5.00129, 5.002997, 
    5.006517, 5.013214, 5.024857, 5.043125, 5.068581, 5.099402, 5.130821, 
    5.156437, 0, 5.645344, 5.631002, 5.571152, 5.445369, 5.241158, 4.948497, 
    4.63036, 4.328893, 4.096667, 3.969621, 3.954431, 4.03174, 4.170502, 
    4.343932, 4.540859, 4.72441, 4.91267, 5.100444, 5.282361, 5.451836, 
    5.599946, 5.7146, 5.780928, 5.784469, 5.718306, 5.591999, 5.434416, 
    5.28287, 5.164471, 5.086521, 5.041785, 5.018754, 5.007888, 5.003124,
  // momentumY(4,23, 0-49)
    5.000003, 5.000014, 5.000041, 5.000118, 5.000312, 5.000783, 5.001848, 
    5.004087, 5.008446, 5.016229, 5.028857, 5.047226, 5.070715, 5.096325, 
    5.118713, 0, 5.596464, 5.578844, 5.518146, 5.392861, 5.187092, 4.88203, 
    4.546795, 4.220427, 3.96124, 3.815448, 3.794108, 3.875613, 4.021391, 
    4.202407, 4.412063, 4.602664, 4.800696, 5.001018, 5.198163, 5.385542, 
    5.554357, 5.692601, 5.784849, 5.814455, 5.769972, 5.655174, 5.495645, 
    5.33144, 5.196806, 5.105144, 5.051356, 5.023251, 5.009851, 5.003916,
  // momentumY(4,24, 0-49)
    5.000002, 5.000011, 5.000033, 5.000093, 5.000248, 5.000626, 5.001483, 
    5.003294, 5.006839, 5.01322, 5.023686, 5.039129, 5.059257, 5.081702, 
    5.101663, 0, 5.556334, 5.537187, 5.476232, 5.351586, 5.145324, 4.83245, 
    4.485684, 4.140932, 3.860631, 3.700632, 3.676901, 3.765053, 3.9187, 
    4.106887, 4.327, 4.52336, 4.728728, 4.937836, 5.14499, 5.343493, 
    5.524635, 5.676622, 5.784046, 5.829436, 5.799034, 5.693022, 5.534179, 
    5.363252, 5.21863, 5.117971, 5.058032, 5.026413, 5.011236, 5.004478,
  // momentumY(4,25, 0-49)
    5.000005, 5.000016, 5.000045, 5.000125, 5.000327, 5.000806, 5.00187, 
    5.004066, 5.00826, 5.015623, 5.027387, 5.044277, 5.06568, 5.088906, 
    5.109101, 0, 5.530094, 5.511153, 5.450953, 5.327627, 5.122614, 4.808633, 
    4.459426, 4.109352, 3.822037, 3.657288, 3.633398, 3.724782, 3.881723, 
    4.07268, 4.296721, 4.495244, 4.70334, 4.915673, 5.126443, 5.328887, 
    5.514308, 5.670983, 5.783531, 5.834264, 5.808712, 5.705871, 5.54749, 
    5.374413, 5.226382, 5.122564, 5.060434, 5.027554, 5.011736, 5.004682,
  // momentumY(4,26, 0-49)
    5.00001, 5.00003, 5.000083, 5.000225, 5.000573, 5.001377, 5.003111, 
    5.006579, 5.012978, 5.023774, 5.040254, 5.062696, 5.089457, 5.116624, 
    5.138906, 0, 5.520136, 5.503262, 5.445169, 5.324215, 5.122498, 4.814704, 
    4.473166, 4.133136, 3.856438, 3.698707, 3.676142, 3.764788, 3.918613, 
    4.10686, 4.326991, 4.523357, 4.728727, 4.937836, 5.144989, 5.343493, 
    5.524634, 5.676622, 5.784046, 5.829436, 5.799034, 5.693022, 5.534179, 
    5.363252, 5.21863, 5.117971, 5.058032, 5.026413, 5.011236, 5.004478,
  // momentumY(4,27, 0-49)
    5.000019, 5.000056, 5.000157, 5.000415, 5.001042, 5.002456, 5.005435, 
    5.011232, 5.021597, 5.038417, 5.062864, 5.094123, 5.128512, 5.160077, 
    5.183197, 0, 5.526995, 5.513671, 5.458173, 5.339542, 5.142099, 4.846486, 
    4.52138, 4.204391, 3.952483, 3.811342, 3.79244, 3.875007, 4.021184, 
    4.202338, 4.412041, 4.602656, 4.800694, 5.001017, 5.198163, 5.385541, 
    5.554357, 5.692601, 5.784849, 5.814455, 5.769972, 5.655174, 5.495645, 
    5.33144, 5.196806, 5.105144, 5.051356, 5.023251, 5.009851, 5.003916,
  // momentumY(4,28, 0-49)
    5.000035, 5.0001, 5.000277, 5.000724, 5.001793, 5.004173, 5.009095, 
    5.018476, 5.034788, 5.060286, 5.095444, 5.137174, 5.178433, 5.210751, 
    5.229156, 0, 5.549765, 5.540964, 5.487337, 5.369511, 5.17579, 4.895623, 
    4.591888, 4.304254, 4.082989, 3.963053, 3.951664, 4.030686, 4.170128, 
    4.343802, 4.540814, 4.724395, 4.912664, 5.100442, 5.28236, 5.451836, 
    5.599946, 5.7146, 5.780928, 5.784469, 5.718305, 5.591999, 5.434416, 
    5.28287, 5.164471, 5.086521, 5.041785, 5.018754, 5.007888, 5.003124,
  // momentumY(4,29, 0-49)
    5.000054, 5.000159, 5.000442, 5.001153, 5.00284, 5.006568, 5.014205, 
    5.028555, 5.05294, 5.08968, 5.137436, 5.189026, 5.232651, 5.257787, 
    5.262488, 0, 5.584862, 5.579939, 5.525392, 5.405305, 5.214372, 4.952533, 
    4.675216, 4.421723, 4.234072, 4.137152, 4.135252, 4.212865, 4.346626, 
    4.51242, 4.695455, 4.870021, 5.045825, 5.217786, 5.380639, 5.527698, 
    5.649745, 5.734621, 5.768576, 5.740706, 5.650436, 5.514049, 5.36256, 
    5.228116, 5.12906, 5.066501, 5.031611, 5.014006, 5.005826, 5.002292,
  // momentumY(4,30, 0-49)
    5.000076, 5.000227, 5.000637, 5.001688, 5.004233, 5.010009, 5.022226, 
    5.046075, 5.08837, 5.154881, 5.244466, 5.342824, 5.423133, 5.457164, 
    5.429102, 5.460217, 5.513269, 5.527208, 5.492916, 5.390181, 5.221525, 
    4.998848, 4.766492, 4.560466, 4.413423, 4.341393, 4.347546, 4.42042, 
    4.543725, 4.696185, 4.860814, 5.02178, 5.181416, 5.334677, 5.476006, 
    5.598026, 5.690766, 5.742093, 5.74039, 5.680089, 5.568351, 5.427535, 
    5.288007, 5.174216, 5.095507, 5.048014, 5.022378, 5.00975, 5.003997, 
    5.001556,
  // momentumY(4,31, 0-49)
    5.000073, 5.000221, 5.000621, 5.001653, 5.00416, 5.009876, 5.02202, 
    5.045835, 5.088351, 5.155962, 5.249051, 5.356033, 5.453192, 5.513427, 
    5.51753, 5.549628, 5.688647, 5.683352, 5.618227, 5.4899, 5.309708, 
    5.098572, 4.885837, 4.704521, 4.580997, 4.524658, 4.537004, 4.608436, 
    4.726605, 4.870749, 5.021959, 5.17297, 5.319542, 5.456137, 5.576294, 
    5.671569, 5.731426, 5.744835, 5.704313, 5.611754, 5.482604, 5.343098, 
    5.219526, 5.12711, 5.067253, 5.032856, 5.014951, 5.00638, 5.002567, 
    5.000986,
  // momentumY(4,32, 0-49)
    5.000058, 5.000175, 5.000499, 5.001343, 5.003422, 5.008226, 5.018595, 
    5.039321, 5.077241, 5.13961, 5.229686, 5.340741, 5.453701, 5.542929, 
    5.586711, 5.634364, 5.810377, 5.794869, 5.715106, 5.578702, 5.402011, 
    5.211908, 5.024439, 4.868459, 4.765963, 4.722025, 4.737376, 4.804413, 
    4.91415, 5.046367, 5.181589, 5.319583, 5.449525, 5.565306, 5.65952, 
    5.722928, 5.745382, 5.718771, 5.641876, 5.524932, 5.389545, 5.261234, 
    5.158674, 5.08793, 5.04487, 5.021269, 5.009429, 5.003929, 5.001545, 
    5.000584,
  // momentumY(4,33, 0-49)
    5.00004, 5.000121, 5.000348, 5.000955, 5.002475, 5.006059, 5.013967, 
    5.030193, 5.060858, 5.113483, 5.193935, 5.30105, 5.422253, 5.535433, 
    5.617548, 5.69124, 5.875936, 5.864213, 5.786301, 5.657351, 5.496267, 
    5.333714, 5.17509, 5.044634, 4.961142, 4.927159, 4.943112, 5.003295, 
    5.101369, 5.218139, 5.334802, 5.456174, 5.565315, 5.655402, 5.718253, 
    5.744672, 5.726639, 5.661288, 5.555245, 5.425946, 5.296785, 5.187774, 
    5.108407, 5.057558, 5.028332, 5.01302, 5.005613, 5.00228, 5.000876, 
    5.000325,
  // momentumY(4,34, 0-49)
    5.000024, 5.000075, 5.000218, 5.000609, 5.001614, 5.004035, 5.009521, 
    5.021117, 5.043819, 5.084566, 5.150602, 5.245469, 5.363938, 5.490148, 
    5.602442, 5.704795, 5.886364, 5.892461, 5.832005, 5.724312, 5.588806, 
    5.458125, 5.330325, 5.225271, 5.159105, 5.133275, 5.148096, 5.1995, 
    5.282907, 5.380851, 5.476084, 5.576321, 5.659528, 5.718254, 5.744268, 
    5.730054, 5.672071, 5.574646, 5.451857, 5.324495, 5.212377, 5.12704, 
    5.069887, 5.035612, 5.016918, 5.007533, 5.003155, 5.001247, 5.000467, 
    5.000169,
  // momentumY(4,35, 0-49)
    5.000014, 5.000041, 5.000124, 5.000355, 5.000961, 5.002462, 5.00596, 
    5.013583, 5.029061, 5.058093, 5.107836, 5.184575, 5.289448, 5.414499, 
    5.54309, 5.668658, 5.844255, 5.878744, 5.849082, 5.774486, 5.672875, 
    5.577171, 5.48142, 5.401774, 5.351748, 5.332812, 5.345255, 5.386293, 
    5.452143, 5.527818, 5.598071, 5.671585, 5.722932, 5.744674, 5.730054, 
    5.67552, 5.58408, 5.467301, 5.343374, 5.230956, 5.142365, 5.080799, 
    5.04248, 5.020813, 5.009551, 5.004119, 5.001675, 5.000645, 5.000236, 
    5.000084,
  // momentumY(4,36, 0-49)
    5.000007, 5.000022, 5.000065, 5.00019, 5.000528, 5.001387, 5.003449, 
    5.008088, 5.01785, 5.036942, 5.071377, 5.128031, 5.211954, 5.322424, 
    5.450345, 5.586574, 5.754741, 5.821698, 5.831575, 5.79887, 5.73787, 
    5.679853, 5.617424, 5.563701, 5.529284, 5.51648, 5.525597, 5.554762, 
    5.600111, 5.649807, 5.69079, 5.731433, 5.745385, 5.72664, 5.672071, 
    5.58408, 5.472425, 5.352917, 5.242486, 5.153233, 5.089346, 5.048308, 
    5.024346, 5.011489, 5.005095, 5.002128, 5.00084, 5.000314, 5.000111, 
    5.000039,
  // momentumY(4,37, 0-49)
    5.000002, 5.000011, 5.000032, 5.000094, 5.00027, 5.000727, 5.001855, 
    5.004479, 5.010196, 5.021828, 5.043808, 5.082083, 5.142909, 5.230166, 
    5.342067, 5.472644, 5.628459, 5.722989, 5.773468, 5.786318, 5.77012, 
    5.752038, 5.724462, 5.697757, 5.679138, 5.672138, 5.677126, 5.692811, 
    5.714684, 5.734652, 5.742105, 5.744839, 5.718772, 5.661288, 5.574646, 
    5.467301, 5.352917, 5.246391, 5.158862, 5.094786, 5.052536, 5.027167, 
    5.013159, 5.00599, 5.002568, 5.001039, 5.000397, 5.000144, 5.00005, 
    5.000018,
  // momentumY(4,38, 0-49)
    5, 5.000005, 5.000015, 5.000044, 5.000129, 5.000355, 5.000931, 5.002315, 
    5.005435, 5.012023, 5.025013, 5.048794, 5.088931, 5.150884, 5.237588, 
    5.348084, 5.483159, 5.591568, 5.673834, 5.728097, 5.756079, 5.778114, 
    5.786222, 5.787565, 5.785347, 5.784119, 5.784297, 5.784952, 5.780969, 
    5.768591, 5.740396, 5.704315, 5.641877, 5.555245, 5.451857, 5.343374, 
    5.242486, 5.158862, 5.096653, 5.05476, 5.028989, 5.014386, 5.006711, 
    5.002948, 5.001224, 5.00048, 5.000178, 5.000063, 5.000022, 5.000008,
  // momentumY(4,39, 0-49)
    5, 5.000001, 5.000007, 5.00002, 5.000057, 5.000163, 5.000438, 5.00112, 
    5.002711, 5.006193, 5.013331, 5.026992, 5.051274, 5.091135, 5.151162, 
    5.233976, 5.340683, 5.445152, 5.541938, 5.624341, 5.688284, 5.745618, 
    5.787155, 5.815814, 5.830077, 5.834549, 5.829556, 5.814503, 5.784487, 
    5.740712, 5.680091, 5.611754, 5.524933, 5.425946, 5.324495, 5.230956, 
    5.153233, 5.094786, 5.05476, 5.029618, 5.015037, 5.00718, 5.003231, 
    5.001372, 5.00055, 5.00021, 5.000076, 5.000027, 5.00001, 5.000003,
  // momentumY(4,40, 0-49)
    5, 5, 5.000002, 5.000009, 5.000025, 5.00007, 5.000193, 5.000509, 
    5.001269, 5.002991, 5.006652, 5.013947, 5.027512, 5.050968, 5.088504, 
    5.143935, 5.219826, 5.305856, 5.397701, 5.488678, 5.572298, 5.652788, 
    5.719582, 5.770612, 5.799332, 5.808841, 5.799087, 5.769994, 5.718313, 
    5.650439, 5.568352, 5.482605, 5.389545, 5.296785, 5.212377, 5.142365, 
    5.089346, 5.052536, 5.028989, 5.015037, 5.007341, 5.00338, 5.001469, 
    5.000603, 5.000236, 5.000087, 5.000031, 5.000011, 5.000004, 5,
  // momentumY(4,41, 0-49)
    5, 5, 5, 5.000003, 5.000011, 5.000029, 5.000081, 5.000217, 5.000558, 
    5.001357, 5.003117, 5.006752, 5.013795, 5.026531, 5.047973, 5.081492, 
    5.130116, 5.191607, 5.264742, 5.345742, 5.429265, 5.515083, 5.592558, 
    5.655453, 5.693151, 5.705927, 5.693044, 5.655183, 5.592001, 5.51405, 
    5.427535, 5.343099, 5.261235, 5.187774, 5.12704, 5.080799, 5.048308, 
    5.027167, 5.014386, 5.00718, 5.00338, 5.001504, 5.000631, 5.00025, 
    5.000094, 5.000034, 5.000013, 5.000005, 5, 5,
  // momentumY(4,42, 0-49)
    5, 5, 5, 5, 5.000005, 5.000012, 5.000032, 5.000088, 5.000232, 5.00058, 
    5.001373, 5.003073, 5.006487, 5.012912, 5.024214, 5.042749, 5.071041, 
    5.10987, 5.16003, 5.220561, 5.28869, 5.362971, 5.434639, 5.495757, 
    5.534231, 5.547513, 5.534188, 5.495649, 5.434417, 5.36256, 5.288007, 
    5.219526, 5.158674, 5.108407, 5.069887, 5.04248, 5.024346, 5.013159, 
    5.006711, 5.003231, 5.001469, 5.000631, 5.000257, 5.000099, 5.000036, 
    5.000014, 5.000005, 5.000001, 5, 5,
  // momentumY(4,43, 0-49)
    5, 5, 5, 5, 5.000001, 5.000005, 5.000013, 5.000034, 5.000092, 5.000234, 
    5.000571, 5.001317, 5.002868, 5.005898, 5.011437, 5.020907, 5.036011, 
    5.058069, 5.088407, 5.127475, 5.17446, 5.228262, 5.28295, 5.331479, 
    5.36327, 5.374421, 5.363255, 5.331441, 5.28287, 5.228115, 5.174216, 
    5.12711, 5.08793, 5.057558, 5.035612, 5.020813, 5.011489, 5.00599, 
    5.002948, 5.001372, 5.000603, 5.00025, 5.000099, 5.000037, 5.000015, 
    5.000006, 5.000001, 5, 5, 5,
  // momentumY(4,44, 0-49)
    5, 5, 5, 5, 5, 5.000001, 5.000006, 5.000014, 5.000034, 5.00009, 5.000225, 
    5.000533, 5.001195, 5.002535, 5.005076, 5.009581, 5.017048, 5.028498, 
    5.045024, 5.067372, 5.095585, 5.129107, 5.164498, 5.196819, 5.218636, 
    5.226383, 5.218631, 5.196807, 5.164472, 5.12906, 5.095506, 5.067253, 
    5.044869, 5.028332, 5.016918, 5.009551, 5.005095, 5.002568, 5.001224, 
    5.00055, 5.000236, 5.000094, 5.000036, 5.000015, 5.000007, 5.000002, 5, 
    5, 5, 5,
  // momentumY(4,45, 0-49)
    5, 5, 5, 5, 5, 5, 5.000002, 5.000006, 5.000013, 5.000032, 5.000083, 
    5.000204, 5.000471, 5.001028, 5.002122, 5.004128, 5.007573, 5.013069, 
    5.021315, 5.032892, 5.048037, 5.066514, 5.086528, 5.105148, 5.117975, 
    5.122566, 5.117973, 5.105145, 5.086521, 5.0665, 5.048013, 5.032856, 
    5.021268, 5.013019, 5.007533, 5.004119, 5.002128, 5.001039, 5.00048, 
    5.00021, 5.000087, 5.000034, 5.000014, 5.000006, 5.000002, 5, 5, 5, 5, 5,
  // momentumY(4,46, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000005, 5.000012, 5.00003, 5.000074, 
    5.000175, 5.000395, 5.000838, 5.001678, 5.003167, 5.005628, 5.009441, 
    5.01496, 5.022381, 5.031613, 5.041788, 5.051359, 5.058036, 5.060439, 
    5.058036, 5.051358, 5.041786, 5.03161, 5.022376, 5.014949, 5.009427, 
    5.005613, 5.003155, 5.001675, 5.00084, 5.000397, 5.000178, 5.000076, 
    5.000031, 5.000013, 5.000005, 5.000001, 5, 5, 5, 5, 5, 5,
  // momentumY(4,47, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5.000001, 5.000005, 5.000011, 5.000026, 5.000062, 
    5.000143, 5.000313, 5.000644, 5.001248, 5.002281, 5.003928, 5.006376, 
    5.009744, 5.014003, 5.018755, 5.023259, 5.026426, 5.027568, 5.026426, 
    5.023259, 5.018755, 5.014002, 5.009743, 5.006373, 5.003924, 5.002277, 
    5.001245, 5.000643, 5.000314, 5.000143, 5.000063, 5.000027, 5.000011, 
    5.000005, 5.000001, 5, 5, 5, 5, 5, 5, 5,
  // momentumY(4,48, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000004, 5.00001, 5.000022, 5.000049, 
    5.000109, 5.000232, 5.000462, 5.000867, 5.001534, 5.002549, 5.003979, 
    5.005815, 5.007891, 5.009873, 5.011274, 5.01178, 5.011274, 5.009873, 
    5.007891, 5.005815, 5.003978, 5.002548, 5.001532, 5.000866, 5.000462, 
    5.000232, 5.000109, 5.000049, 5.000022, 5.00001, 5.000004, 5, 5, 5, 5, 5, 
    5, 5, 5, 5,
  // momentumY(4,49, 0-49)
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5.000002, 5.000005, 5.000012, 5.00003, 
    5.000065, 5.000139, 5.000275, 5.000512, 5.000896, 5.001465, 5.002233, 
    5.00314, 5.004033, 5.004668, 5.004897, 5.004668, 5.004033, 5.00314, 
    5.002233, 5.001465, 5.000896, 5.000512, 5.000275, 5.000139, 5.000065, 
    5.00003, 5.000012, 5.000005, 5.000002, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5,
  // momentumY(5,0, 0-49)
    5, 5, 5, 5, 5, 5, 5.000002, 5.000006, 5.000013, 5.000028, 5.000061, 
    5.00013, 5.000265, 5.000516, 5.00096, 5.001699, 5.002862, 5.004584, 
    5.006996, 5.010178, 5.014109, 5.018611, 5.023259, 5.027408, 5.030265, 
    5.031285, 5.030264, 5.027405, 5.023253, 5.018603, 5.014096, 5.010162, 
    5.006977, 5.004565, 5.002849, 5.001694, 5.000961, 5.00052, 5.000268, 
    5.000132, 5.000062, 5.000028, 5.000013, 5.000006, 5.000002, 5, 5, 5, 5, 5,
  // momentumY(5,1, 0-49)
    5, 5, 5, 5, 5, 5.000004, 5.000008, 5.000015, 5.000031, 5.000068, 
    5.000149, 5.000312, 5.000626, 5.0012, 5.002189, 5.003802, 5.006291, 
    5.0099, 5.01486, 5.021302, 5.029162, 5.038113, 5.047316, 5.055529, 
    5.06116, 5.063167, 5.061155, 5.05552, 5.047298, 5.038086, 5.029122, 
    5.021251, 5.0148, 5.00984, 5.006246, 5.003785, 5.002189, 5.001209, 
    5.000637, 5.00032, 5.000154, 5.000071, 5.000032, 5.000015, 5.000008, 
    5.000004, 5, 5, 5, 5,
  // momentumY(5,2, 0-49)
    5, 5, 5, 5, 5.000005, 5.000009, 5.000016, 5.000033, 5.000074, 5.000168, 
    5.000363, 5.000746, 5.001466, 5.00274, 5.004883, 5.00829, 5.013408, 
    5.020618, 5.030261, 5.042474, 5.057049, 5.073393, 5.08998, 5.104668, 
    5.114639, 5.118178, 5.114626, 5.10464, 5.089929, 5.07331, 5.056931, 
    5.042319, 5.030082, 5.020443, 5.013276, 5.008237, 5.00488, 5.002761, 
    5.001492, 5.000769, 5.000379, 5.000178, 5.000082, 5.000035, 5.000017, 
    5.000009, 5.000005, 5.000001, 5, 5,
  // momentumY(5,3, 0-49)
    5, 5, 5, 5.000004, 5.000009, 5.000016, 5.000034, 5.000081, 5.000184, 
    5.000405, 5.000853, 5.001713, 5.00328, 5.005985, 5.010404, 5.017234, 
    5.027194, 5.040734, 5.058229, 5.079662, 5.104465, 5.131642, 5.158663, 
    5.182254, 5.198014, 5.203566, 5.197978, 5.182171, 5.158515, 5.131409, 
    5.104133, 5.079228, 5.057729, 5.040246, 5.026826, 5.017087, 5.010396, 
    5.006039, 5.00335, 5.001772, 5.000896, 5.000432, 5.000201, 5.000089, 
    5.000038, 5.000018, 5.00001, 5.000006, 5.000001, 5,
  // momentumY(5,4, 0-49)
    5, 5, 5.000002, 5.000008, 5.000016, 5.000034, 5.000082, 5.000193, 
    5.000432, 5.000931, 5.001913, 5.003746, 5.006992, 5.012434, 5.021055, 
    5.033954, 5.052146, 5.075799, 5.105033, 5.139303, 5.177319, 5.217662, 
    5.25659, 5.289864, 5.311574, 5.319134, 5.311477, 5.289647, 5.256206, 
    5.217056, 5.176451, 5.13817, 5.103726, 5.074522, 5.051179, 5.033571, 
    5.021023, 5.012565, 5.007167, 5.003901, 5.002026, 5.001004, 5.000476, 
    5.000216, 5.000093, 5.00004, 5.000018, 5.00001, 5.000005, 5,
  // momentumY(5,5, 0-49)
    5, 5.000001, 5.000006, 5.000015, 5.000033, 5.000081, 5.000193, 5.000442, 
    5.000971, 5.002039, 5.004083, 5.00779, 5.014157, 5.024488, 5.040304, 
    5.063102, 5.094024, 5.131987, 5.176251, 5.225178, 5.276432, 5.328592, 
    5.376917, 5.417064, 5.442416, 5.451099, 5.442188, 5.416547, 5.376002, 
    5.32715, 5.274362, 5.222458, 5.173093, 5.128881, 5.09165, 5.062176, 
    5.040218, 5.024799, 5.014578, 5.008171, 5.004367, 5.002228, 5.001084, 
    5.000504, 5.000224, 5.000095, 5.00004, 5.000018, 5.000009, 5.000004,
  // momentumY(5,6, 0-49)
    5.000001, 5.000005, 5.000013, 5.000031, 5.000074, 5.000183, 5.00043, 
    5.000967, 5.002075, 5.004246, 5.008282, 5.015374, 5.02715, 5.045572, 
    5.072659, 5.110019, 5.15846, 5.213607, 5.273174, 5.334088, 5.393208, 
    5.450352, 5.500582, 5.540859, 5.565177, 5.573293, 5.564681, 5.539737, 
    5.498604, 5.447233, 5.388718, 5.328151, 5.266213, 5.206674, 5.153087, 
    5.107989, 5.072482, 5.046282, 5.028121, 5.016266, 5.008961, 5.004705, 
    5.002356, 5.001125, 5.000514, 5.000224, 5.000093, 5.000038, 5.000018, 
    5.000008,
  // momentumY(5,7, 0-49)
    5.000004, 5.00001, 5.000028, 5.000067, 5.000166, 5.0004, 5.000918, 
    5.002015, 5.004214, 5.008401, 5.015932, 5.02872, 5.04916, 5.079797, 
    5.122718, 5.178854, 5.248075, 5.319426, 5.389174, 5.453479, 5.509659, 
    5.560696, 5.602446, 5.634424, 5.65239, 5.658066, 5.651396, 5.632189, 
    5.598525, 5.554535, 5.500804, 5.441733, 5.375283, 5.305392, 5.237004, 
    5.174875, 5.122472, 5.081369, 5.051301, 5.030718, 5.017484, 5.009469, 
    5.004883, 5.002399, 5.001125, 5.000504, 5.000216, 5.000089, 5.000036, 
    5.000016,
  // momentumY(5,8, 0-49)
    5.000009, 5.000022, 5.000058, 5.000145, 5.000354, 5.000831, 5.001863, 
    5.003988, 5.008126, 5.015749, 5.028997, 5.050632, 5.083705, 5.130813, 
    5.193053, 5.269456, 5.35902, 5.440007, 5.509358, 5.56441, 5.604834, 
    5.638444, 5.662354, 5.67907, 5.686673, 5.688493, 5.684813, 5.674917, 
    5.655134, 5.627209, 5.588828, 5.543271, 5.484299, 5.414421, 5.338465, 
    5.262632, 5.193025, 5.134175, 5.088205, 5.054886, 5.03237, 5.018123, 
    5.009644, 5.004883, 5.002356, 5.001084, 5.000476, 5.000201, 5.000082, 
    5.000034,
  // momentumY(5,9, 0-49)
    5.000019, 5.000048, 5.00012, 5.000298, 5.000716, 5.001643, 5.003593, 
    5.007489, 5.014842, 5.027926, 5.049793, 5.083932, 5.133445, 5.199761, 
    5.281408, 5.374544, 5.47942, 5.558947, 5.615193, 5.648915, 5.663444, 
    5.671911, 5.672351, 5.669973, 5.665254, 5.662431, 5.661954, 5.662679, 
    5.659845, 5.652761, 5.636622, 5.613993, 5.574114, 5.516903, 5.445178, 
    5.364569, 5.282547, 5.20661, 5.142382, 5.092508, 5.056751, 5.032938, 
    5.018123, 5.009469, 5.004705, 5.002228, 5.001004, 5.000433, 5.00018, 
    5.000075,
  // momentumY(5,10, 0-49)
    5.000036, 5.000093, 5.000239, 5.000585, 5.001373, 5.003076, 5.006561, 
    5.013308, 5.02562, 5.046711, 5.08042, 5.130344, 5.198357, 5.283011, 
    5.378876, 5.479668, 5.591911, 5.658225, 5.691349, 5.696425, 5.68037, 
    5.66087, 5.636159, 5.613672, 5.596256, 5.58842, 5.590661, 5.601462, 
    5.615591, 5.630049, 5.638243, 5.642887, 5.629557, 5.59555, 5.540604, 
    5.467718, 5.383308, 5.296116, 5.215004, 5.146606, 5.093976, 5.056751, 
    5.03237, 5.017484, 5.008961, 5.004367, 5.002027, 5.000896, 5.000381, 
    5.000162,
  // momentumY(5,11, 0-49)
    5.000071, 5.000181, 5.000453, 5.001088, 5.002494, 5.005449, 5.011323, 
    5.022336, 5.041712, 5.073508, 5.121789, 5.189017, 5.274099, 5.371275, 
    5.471056, 5.567159, 5.679311, 5.724144, 5.729917, 5.705225, 5.659316, 
    5.612999, 5.564149, 5.522204, 5.492456, 5.479336, 5.483345, 5.502607, 
    5.531834, 5.56584, 5.596796, 5.628322, 5.64375, 5.638568, 5.609673, 
    5.556548, 5.482425, 5.39456, 5.302978, 5.217842, 5.146606, 5.092508, 
    5.054886, 5.030718, 5.016266, 5.008171, 5.003901, 5.001774, 5.000774, 
    5.000335,
  // momentumY(5,12, 0-49)
    5.000131, 5.00033, 5.000812, 5.001908, 5.004274, 5.00911, 5.018438, 
    5.035336, 5.0639, 5.108568, 5.172517, 5.255433, 5.351807, 5.45142, 
    5.54234, 5.622025, 5.729712, 5.750149, 5.730207, 5.67971, 5.608513, 
    5.538956, 5.468381, 5.40834, 5.366759, 5.347938, 5.352461, 5.37809, 
    5.419709, 5.470071, 5.520361, 5.575464, 5.617815, 5.642097, 5.643387, 
    5.618141, 5.565696, 5.48967, 5.398307, 5.302978, 5.215004, 5.142382, 
    5.088205, 5.051301, 5.028121, 5.014579, 5.007169, 5.003353, 5.001502, 
    5.000663,
  // momentumY(5,13, 0-49)
    5.000229, 5.000569, 5.001369, 5.00315, 5.006894, 5.014339, 5.02826, 
    5.052577, 5.091915, 5.1502, 5.228284, 5.321659, 5.420121, 5.510469, 
    5.580884, 5.636158, 5.738116, 5.735927, 5.695858, 5.626519, 5.536742, 
    5.448798, 5.359662, 5.283228, 5.230228, 5.205044, 5.208557, 5.238231, 
    5.289241, 5.352497, 5.418259, 5.492509, 5.55786, 5.608896, 5.639956, 
    5.645646, 5.622089, 5.568675, 5.48967, 5.39456, 5.296116, 5.20661, 
    5.134175, 5.081369, 5.046282, 5.0248, 5.012568, 5.006046, 5.00278, 
    5.001256,
  // momentumY(5,14, 0-49)
    5.000374, 5.000917, 5.002163, 5.004873, 5.010436, 5.021191, 5.040668, 
    5.073408, 5.123923, 5.194474, 5.282308, 5.378265, 5.468612, 5.539557, 
    5.581494, 5.609149, 5.704862, 5.684734, 5.631863, 5.551764, 5.45104, 
    5.350298, 5.246478, 5.15581, 5.091814, 5.059381, 5.060057, 5.091223, 
    5.148467, 5.22124, 5.298869, 5.387869, 5.471773, 5.545377, 5.60301, 
    5.638582, 5.646293, 5.622088, 5.565695, 5.482424, 5.383307, 5.282547, 
    5.193025, 5.122472, 5.072483, 5.040219, 5.021027, 5.010407, 5.004912, 
    5.002266,
  // momentumY(5,15, 0-49)
    5.000567, 5.001374, 5.003187, 5.00704, 5.014763, 5.029299, 5.054786, 
    5.09597, 5.156433, 5.235746, 5.326997, 5.417121, 5.49086, 5.535902, 
    5.545708, 5.546775, 5.632914, 5.60088, 5.542744, 5.459904, 5.356049, 
    5.248635, 5.134977, 5.033073, 4.95883, 4.918158, 4.913803, 4.943549, 
    5.003622, 5.082602, 5.168946, 5.268797, 5.367137, 5.458964, 5.538911, 
    5.600954, 5.638575, 5.645641, 5.618137, 5.556546, 5.467716, 5.364568, 
    5.262632, 5.174875, 5.10799, 5.062179, 5.033578, 5.017106, 5.008286, 
    5.003901,
  // momentumY(5,16, 0-49)
    5.000793, 5.001904, 5.004345, 5.009432, 5.01941, 5.037717, 5.06884, 
    5.117216, 5.184804, 5.268004, 5.356136, 5.433732, 5.48586, 5.502688, 
    5.480472, 5.459173, 5.525829, 5.488203, 5.431913, 5.353796, 5.254422, 
    5.146871, 5.029435, 4.92056, 4.837578, 4.787774, 4.775797, 4.80067, 
    4.859735, 4.941498, 5.033751, 5.14112, 5.250391, 5.356567, 5.454606, 
    5.538887, 5.602984, 5.639937, 5.643376, 5.609665, 5.5406, 5.445177, 
    5.338465, 5.237003, 5.153089, 5.091654, 5.05119, 5.026856, 5.013346, 
    5.006411,
  // momentumY(5,17, 0-49)
    5.001009, 5.002405, 5.005424, 5.01161, 5.023516, 5.044888, 5.080247, 
    5.133332, 5.204224, 5.28643, 5.36658, 5.428285, 5.457914, 5.448078, 
    5.397178, 5.359798, 5.38727, 5.349489, 5.301646, 5.235264, 5.147697, 
    5.046798, 4.932895, 4.822896, 4.733915, 4.674499, 4.651908, 4.667727, 
    4.721311, 4.802092, 4.897588, 5.009571, 5.126815, 5.244068, 5.35647, 
    5.458864, 5.5453, 5.608845, 5.642067, 5.638551, 5.595541, 5.5169, 
    5.414419, 5.305392, 5.206675, 5.128885, 5.074537, 5.040285, 5.020535, 
    5.010053,
  // momentumY(5,18, 0-49)
    5.001149, 5.002726, 5.006095, 5.012916, 5.025878, 5.048788, 5.085967, 
    5.140407, 5.210714, 5.288495, 5.358942, 5.405567, 5.415976, 5.384698, 
    5.312162, 5.264491, 5.221843, 5.186554, 5.153127, 5.1055, 5.037116, 
    4.949855, 4.847899, 4.744311, 4.653742, 4.585035, 4.548517, 4.550172, 
    4.592954, 4.668444, 4.76445, 4.87837, 5.000965, 5.126472, 5.250022, 
    5.366846, 5.471569, 5.55773, 5.617738, 5.643708, 5.629535, 5.574101, 
    5.484294, 5.375281, 5.266214, 5.1731, 5.103745, 5.057774, 5.03019, 
    5.015046,
  // momentumY(5,19, 0-49)
    5.001132, 5.00268, 5.005971, 5.012604, 5.025155, 5.04725, 5.082956, 
    5.134978, 5.201641, 5.274235, 5.337543, 5.374701, 5.373543, 5.330182, 
    5.248117, 5.187968, 5.03577, 5.00039, 4.986063, 4.964749, 4.923753, 
    4.857672, 4.777114, 4.68915, 4.603427, 4.527005, 4.473067, 4.454343, 
    4.479911, 4.545097, 4.638662, 4.751842, 4.87722, 5.008308, 5.14009, 
    5.268059, 5.38738, 5.492204, 5.575282, 5.62822, 5.642832, 5.613966, 
    5.543258, 5.441728, 5.32815, 5.222465, 5.138189, 5.079276, 5.042429, 
    5.021496,
  // momentumY(5,20, 0-49)
    5.000885, 5.002056, 5.004517, 5.009397, 5.018436, 5.033949, 5.05833, 
    5.092862, 5.13604, 5.182454, 5.22361, 5.251111, 5.26051, 5.253445, 
    5.236856, 0, 4.882641, 4.890296, 4.897371, 4.893323, 4.87047, 4.819962, 
    4.758723, 4.686413, 4.605082, 4.517176, 4.437809, 4.388928, 4.388727, 
    4.437592, 4.525457, 4.634996, 4.760348, 4.894176, 5.031245, 5.167237, 
    5.297763, 5.417573, 5.519956, 5.596563, 5.638118, 5.636558, 5.588799, 
    5.500793, 5.388714, 5.274365, 5.176466, 5.104169, 5.057017, 5.029309,
  // momentumY(5,21, 0-49)
    5.000641, 5.001482, 5.003266, 5.006831, 5.013499, 5.025104, 5.043731, 
    5.070997, 5.106867, 5.148563, 5.190476, 5.225755, 5.249031, 5.258772, 
    5.257997, 0, 4.74108, 4.76133, 4.784954, 4.801523, 4.801844, 4.771854, 
    4.732392, 4.676557, 4.600542, 4.503641, 4.402691, 4.328095, 4.306149, 
    4.341571, 4.42612, 4.532413, 4.657756, 4.794104, 4.93592, 5.078889, 
    5.218863, 5.351027, 5.469194, 5.565336, 5.629769, 5.652613, 5.627135, 
    5.554501, 5.447219, 5.327146, 5.217059, 5.131421, 5.073335, 5.038131,
  // momentumY(5,22, 0-49)
    5.000444, 5.00103, 5.002293, 5.004852, 5.009718, 5.018359, 5.0326, 
    5.054197, 5.084013, 5.121048, 5.161894, 5.201262, 5.233709, 5.255754, 
    5.267343, 0, 4.627163, 4.653697, 4.689208, 4.723159, 4.745467, 4.737381, 
    4.725026, 4.694858, 4.635277, 4.538174, 4.417841, 4.312981, 4.261384, 
    4.275565, 4.351222, 4.44836, 4.569024, 4.704297, 4.848145, 4.995989, 
    5.143591, 5.286217, 5.41789, 5.530775, 5.614996, 5.659525, 5.65497, 
    5.598444, 5.498568, 5.375984, 5.256189, 5.158487, 5.089858, 5.047126,
  // momentumY(5,23, 0-49)
    5.000326, 5.000756, 5.0017, 5.003643, 5.007394, 5.014186, 5.025643, 
    5.043532, 5.069174, 5.102598, 5.141809, 5.182737, 5.220225, 5.249777, 
    5.26927, 0, 4.542715, 4.572813, 4.616893, 4.664588, 4.705509, 4.716725, 
    4.729808, 4.725214, 4.68426, 4.591591, 4.457345, 4.326142, 4.246144, 
    4.238336, 4.303779, 4.389193, 4.502711, 4.634574, 4.778222, 4.928749, 
    5.081713, 5.232281, 5.374473, 5.500473, 5.600245, 5.662012, 5.674566, 
    5.632014, 5.539653, 5.416502, 5.289604, 5.182093, 5.104459, 5.055098,
  // momentumY(5,24, 0-49)
    5.000295, 5.00068, 5.00153, 5.00328, 5.006674, 5.012842, 5.023315, 
    5.039814, 5.063758, 5.095514, 5.133634, 5.174624, 5.213623, 5.245886, 
    5.268474, 0, 4.488168, 4.520331, 4.569875, 4.626774, 4.680708, 4.705749, 
    4.737486, 4.751808, 4.725004, 4.637198, 4.495549, 4.347715, 4.248083, 
    4.223984, 4.28151, 4.357102, 4.464386, 4.592849, 4.73542, 4.886861, 
    5.042512, 5.19742, 5.345583, 5.479222, 5.588269, 5.660618, 5.684098, 
    5.651032, 5.564503, 5.442098, 5.311407, 5.19786, 5.114362, 5.060548,
  // momentumY(5,25, 0-49)
    5.000359, 5.000815, 5.001808, 5.003817, 5.007643, 5.014476, 5.025854, 
    5.043424, 5.068394, 5.100799, 5.138853, 5.178908, 5.216267, 5.246636, 
    5.267615, 0, 4.464517, 4.497284, 4.548565, 4.608568, 4.667108, 4.6971, 
    4.73595, 4.757792, 4.737058, 4.652288, 4.509429, 4.356791, 4.250607, 
    4.22062, 4.27515, 4.34684, 4.451613, 4.57867, 4.72073, 4.872409, 
    5.028946, 5.185324, 5.335518, 5.471749, 5.583937, 5.659878, 5.6871, 
    5.657343, 5.572935, 5.450924, 5.319024, 5.203423, 5.117879, 5.062491,
  // momentumY(5,26, 0-49)
    5.000526, 5.001181, 5.002566, 5.005302, 5.010374, 5.01916, 5.033297, 
    5.054275, 5.082738, 5.117734, 5.156352, 5.194211, 5.226768, 5.250868, 
    5.265858, 0, 4.47485, 4.506453, 4.555189, 4.611245, 4.664432, 4.688535, 
    4.720223, 4.735377, 4.710451, 4.625587, 4.487513, 4.343034, 4.245784, 
    4.222999, 4.281123, 4.356955, 4.46433, 4.592826, 4.735413, 4.886859, 
    5.042512, 5.19742, 5.345583, 5.479222, 5.588269, 5.660618, 5.684098, 
    5.651031, 5.564503, 5.442098, 5.311407, 5.19786, 5.114362, 5.060548,
  // momentumY(5,27, 0-49)
    5.000805, 5.001794, 5.003833, 5.007775, 5.014898, 5.026875, 5.045452, 
    5.071789, 5.105519, 5.144054, 5.182762, 5.21631, 5.240609, 5.254356, 
    5.259472, 0, 4.523546, 4.551486, 4.592946, 4.637959, 4.676403, 4.684864, 
    4.697034, 4.693454, 4.655822, 4.568797, 4.441556, 4.316923, 4.241585, 
    4.236356, 4.302987, 4.388885, 4.502593, 4.634529, 4.778204, 4.928742, 
    5.081711, 5.232281, 5.374472, 5.500473, 5.600244, 5.662012, 5.674566, 
    5.632014, 5.539653, 5.416502, 5.289604, 5.182093, 5.104459, 5.055098,
  // momentumY(5,28, 0-49)
    5.001189, 5.002643, 5.005589, 5.011191, 5.021119, 5.037401, 5.061837, 
    5.094956, 5.134828, 5.176611, 5.213614, 5.239749, 5.252041, 5.251792, 
    5.243953, 0, 4.61626, 4.63638, 4.665257, 4.692745, 4.709127, 4.695071, 
    4.679724, 4.649843, 4.594497, 4.505446, 4.395233, 4.299756, 4.254767, 
    4.27263, 4.350018, 4.447882, 4.568835, 4.704223, 4.848115, 4.995977, 
    5.143586, 5.286216, 5.417889, 5.530774, 5.614996, 5.659525, 5.65497, 
    5.598445, 5.498568, 5.375984, 5.256189, 5.158487, 5.089858, 5.047126,
  // momentumY(5,29, 0-49)
    5.001638, 5.003657, 5.007708, 5.01534, 5.02871, 5.05025, 5.081713, 
    5.122604, 5.168763, 5.212454, 5.244812, 5.259601, 5.255975, 5.238696, 
    5.215979, 0, 4.757369, 4.761571, 4.770969, 4.774717, 4.763777, 4.723468, 
    4.678093, 4.621346, 4.550265, 4.463518, 4.37518, 4.311992, 4.297986, 
    4.337866, 4.424553, 4.531772, 4.657499, 4.794, 4.935878, 5.078872, 
    5.218856, 5.351024, 5.469192, 5.565335, 5.629769, 5.652613, 5.627135, 
    5.554501, 5.447219, 5.327146, 5.217059, 5.131421, 5.073335, 5.038131,
  // momentumY(5,30, 0-49)
    5.002085, 5.004748, 5.010147, 5.020489, 5.03899, 5.069524, 5.115261, 
    5.176115, 5.24598, 5.31214, 5.358694, 5.372374, 5.346906, 5.283526, 
    5.188242, 5.105539, 4.913468, 4.864236, 4.846265, 4.829531, 4.79874, 
    4.743309, 4.680916, 4.612876, 4.541994, 4.469274, 4.40619, 4.370837, 
    4.379624, 4.433442, 4.523681, 4.634262, 4.760047, 4.894053, 5.031196, 
    5.167217, 5.297757, 5.417571, 5.519956, 5.596563, 5.638118, 5.636558, 
    5.588799, 5.500793, 5.388714, 5.274365, 5.176466, 5.104169, 5.057017, 
    5.029309,
  // momentumY(5,31, 0-49)
    5.002143, 5.004889, 5.010488, 5.021266, 5.040632, 5.072723, 5.12099, 
    5.185519, 5.260214, 5.332315, 5.385979, 5.407974, 5.391459, 5.335916, 
    5.244624, 5.177097, 5.096328, 5.048657, 5.011378, 4.966193, 4.904812, 
    4.824902, 4.735695, 4.645541, 4.563855, 4.495916, 4.451912, 4.441776, 
    4.473276, 4.541901, 4.637214, 4.751214, 4.876952, 5.008195, 5.140043, 
    5.268041, 5.387373, 5.492201, 5.575282, 5.62822, 5.642832, 5.613966, 
    5.543258, 5.441728, 5.328151, 5.222465, 5.138189, 5.079276, 5.042429, 
    5.021496,
  // momentumY(5,32, 0-49)
    5.001922, 5.004405, 5.009535, 5.019537, 5.037773, 5.068523, 5.115789, 
    5.180799, 5.258986, 5.338832, 5.40467, 5.442245, 5.443079, 5.405014, 
    5.329818, 5.271312, 5.264867, 5.214771, 5.161846, 5.095674, 5.012313, 
    4.915738, 4.80939, 4.706865, 4.621886, 4.561248, 4.53286, 4.540988, 
    4.588072, 4.666042, 4.76333, 4.877868, 5.000745, 5.126377, 5.249983, 
    5.366829, 5.471562, 5.557727, 5.617737, 5.643708, 5.629536, 5.574101, 
    5.484294, 5.375281, 5.266214, 5.1731, 5.103745, 5.057774, 5.03019, 
    5.015046,
  // momentumY(5,33, 0-49)
    5.00155, 5.003578, 5.007845, 5.01632, 5.032094, 5.059364, 5.102615, 
    5.16453, 5.242973, 5.328912, 5.40777, 5.464293, 5.487687, 5.473557, 
    5.422353, 5.376557, 5.412996, 5.361646, 5.298301, 5.217968, 5.119894, 
    5.013451, 4.898541, 4.791826, 4.709034, 4.656785, 4.640617, 4.661203, 
    4.717844, 4.800365, 4.89677, 5.009197, 5.126649, 5.243997, 5.35644, 
    5.458851, 5.545294, 5.608843, 5.642066, 5.638551, 5.595541, 5.5169, 
    5.414419, 5.305392, 5.206675, 5.128885, 5.074537, 5.040285, 5.020535, 
    5.010053,
  // momentumY(5,34, 0-49)
    5.001143, 5.002663, 5.005934, 5.012573, 5.025232, 5.04776, 5.084791, 
    5.14025, 5.21467, 5.302464, 5.391526, 5.466604, 5.514605, 5.528172, 
    5.505728, 5.478414, 5.53635, 5.487955, 5.419987, 5.331903, 5.225847, 
    5.115927, 5, 4.895658, 4.818719, 4.774924, 4.767848, 4.796153, 4.857343, 
    4.940302, 5.033179, 5.140856, 5.250273, 5.356515, 5.454584, 5.538877, 
    5.60298, 5.639935, 5.643376, 5.609665, 5.5406, 5.445177, 5.338465, 
    5.237003, 5.153089, 5.091654, 5.05119, 5.026856, 5.013346, 5.006411,
  // momentumY(5,35, 0-49)
    5.000779, 5.001836, 5.004165, 5.009008, 5.018488, 5.035882, 5.065555, 
    5.112102, 5.1783, 5.262308, 5.355819, 5.445318, 5.51646, 5.558745, 
    5.567586, 5.563785, 5.631766, 5.591699, 5.525231, 5.435889, 5.328604, 
    5.221323, 5.110783, 5.013813, 4.944966, 4.909076, 4.90834, 4.940494, 
    5.002017, 5.0818, 5.168562, 5.26862, 5.367057, 5.45893, 5.538898, 
    5.600948, 5.638573, 5.645639, 5.618137, 5.556546, 5.467717, 5.364568, 
    5.262632, 5.174875, 5.10799, 5.062179, 5.033578, 5.017106, 5.008286, 
    5.003901,
  // momentumY(5,36, 0-49)
    5.000493, 5.00118, 5.002732, 5.006036, 5.012685, 5.025267, 5.047535, 
    5.084073, 5.139023, 5.213765, 5.304395, 5.400975, 5.489923, 5.558537, 
    5.598734, 5.621789, 5.695973, 5.669862, 5.611474, 5.527821, 5.42626, 
    5.327377, 5.227425, 5.141449, 5.081936, 5.053137, 5.056394, 5.089209, 
    5.147419, 5.22072, 5.298621, 5.387753, 5.471721, 5.545353, 5.603, 
    5.638578, 5.646291, 5.622087, 5.565695, 5.482424, 5.383308, 5.282547, 
    5.193025, 5.122472, 5.072483, 5.040219, 5.021027, 5.010407, 5.004912, 
    5.002266,
  // momentumY(5,37, 0-49)
    5.000292, 5.00071, 5.00168, 5.003798, 5.008177, 5.016725, 5.032395, 
    5.059221, 5.101714, 5.163327, 5.244109, 5.338745, 5.436703, 5.525202, 
    5.5934, 5.644053, 5.725108, 5.718331, 5.675017, 5.604451, 5.51567, 
    5.430519, 5.345299, 5.272915, 5.223416, 5.200871, 5.206166, 5.236938, 
    5.288577, 5.352169, 5.418102, 5.492436, 5.557827, 5.608882, 5.639949, 
    5.645644, 5.622088, 5.568674, 5.489669, 5.39456, 5.296116, 5.20661, 
    5.134175, 5.081369, 5.046282, 5.0248, 5.012568, 5.006046, 5.00278, 
    5.001256,
  // momentumY(5,38, 0-49)
    5.000163, 5.000402, 5.000972, 5.002252, 5.004967, 5.01043, 5.02079, 
    5.039236, 5.069869, 5.116913, 5.18307, 5.267374, 5.363808, 5.462077, 
    5.550688, 5.62586, 5.715589, 5.73241, 5.710911, 5.660795, 5.591628, 
    5.525109, 5.458025, 5.401213, 5.362216, 5.345235, 5.350946, 5.377285, 
    5.419301, 5.469871, 5.520268, 5.57542, 5.617796, 5.642089, 5.643384, 
    5.61814, 5.565695, 5.489669, 5.398307, 5.302978, 5.215004, 5.142382, 
    5.088205, 5.051301, 5.028121, 5.014579, 5.007169, 5.003353, 5.001502, 
    5.000663,
  // momentumY(5,39, 0-49)
    5.000086, 5.000216, 5.000532, 5.00126, 5.002849, 5.006141, 5.012588, 
    5.024494, 5.045127, 5.078468, 5.128332, 5.196746, 5.282134, 5.37842, 
    5.476128, 5.568144, 5.666311, 5.708275, 5.713571, 5.690119, 5.646567, 
    5.603043, 5.557014, 5.517471, 5.489532, 5.477641, 5.482416, 5.502121, 
    5.53159, 5.565724, 5.596741, 5.628298, 5.64374, 5.638564, 5.60967, 
    5.556547, 5.482424, 5.39456, 5.302978, 5.217841, 5.146606, 5.092508, 
    5.054886, 5.030718, 5.016266, 5.008171, 5.003901, 5.001774, 5.000774, 
    5.000335,
  // momentumY(5,40, 0-49)
    5.000043, 5.00011, 5.000275, 5.000667, 5.001546, 5.00342, 5.007205, 
    5.014437, 5.02746, 5.049472, 5.084197, 5.134979, 5.203325, 5.287435, 
    5.381662, 5.479102, 5.581413, 5.64549, 5.67866, 5.685199, 5.671315, 
    5.65408, 5.631466, 5.610655, 5.594442, 5.587394, 5.59011, 5.601179, 
    5.615451, 5.629982, 5.638213, 5.642873, 5.629552, 5.595548, 5.540603, 
    5.467717, 5.383308, 5.296116, 5.215004, 5.146606, 5.093976, 5.056751, 
    5.03237, 5.017484, 5.008961, 5.004367, 5.002027, 5.000896, 5.000381, 
    5.000162,
  // momentumY(5,41, 0-49)
    5.000021, 5.000053, 5.000136, 5.000334, 5.000796, 5.001806, 5.003906, 
    5.008049, 5.015777, 5.029372, 5.051832, 5.086515, 5.136288, 5.202295, 
    5.282791, 5.373473, 5.471925, 5.54978, 5.606205, 5.641187, 5.657415, 
    5.667536, 5.669413, 5.668134, 5.664176, 5.661833, 5.66164, 5.662522, 
    5.65977, 5.652724, 5.636606, 5.613986, 5.57411, 5.516902, 5.445177, 
    5.364569, 5.282547, 5.20661, 5.142382, 5.092508, 5.056751, 5.032938, 
    5.018123, 5.009469, 5.004705, 5.002228, 5.001004, 5.000433, 5.00018, 
    5.000075,
  // momentumY(5,42, 0-49)
    5.00001, 5.000026, 5.000064, 5.00016, 5.000389, 5.000905, 5.002008, 
    5.004252, 5.008577, 5.016464, 5.030032, 5.051978, 5.08522, 5.132163, 
    5.193682, 5.268489, 5.354282, 5.43411, 5.503586, 5.559516, 5.601096, 
    5.635793, 5.660614, 5.678005, 5.686062, 5.688162, 5.684644, 5.674834, 
    5.655095, 5.62719, 5.588821, 5.543266, 5.484297, 5.41442, 5.338465, 
    5.262631, 5.193025, 5.134175, 5.088205, 5.054886, 5.03237, 5.018123, 
    5.009644, 5.004883, 5.002356, 5.001084, 5.000476, 5.000201, 5.000082, 
    5.000034,
  // momentumY(5,43, 0-49)
    5.000005, 5.000013, 5.00003, 5.000073, 5.000181, 5.000431, 5.000981, 
    5.002132, 5.00442, 5.008735, 5.016428, 5.029381, 5.049916, 5.080473, 
    5.122991, 5.178202, 5.245416, 5.316042, 5.385835, 5.450653, 5.507519, 
    5.559199, 5.60148, 5.633844, 5.652066, 5.657897, 5.651314, 5.632151, 
    5.598507, 5.554525, 5.500799, 5.441729, 5.37528, 5.30539, 5.237002, 
    5.174874, 5.122472, 5.081368, 5.051301, 5.030718, 5.017484, 5.009469, 
    5.004883, 5.002399, 5.001125, 5.000504, 5.000216, 5.000089, 5.000036, 
    5.000016,
  // momentumY(5,44, 0-49)
    5.000001, 5.000006, 5.000015, 5.000033, 5.000081, 5.000196, 5.000456, 
    5.001016, 5.002163, 5.004395, 5.008506, 5.01568, 5.027507, 5.045893, 
    5.072774, 5.109653, 5.157123, 5.211867, 5.271431, 5.332604, 5.392085, 
    5.449572, 5.500086, 5.540573, 5.56503, 5.573226, 5.564657, 5.539729, 
    5.498598, 5.447226, 5.38871, 5.328142, 5.266205, 5.206667, 5.153083, 
    5.107986, 5.07248, 5.046281, 5.028121, 5.016266, 5.008961, 5.004705, 
    5.002356, 5.001125, 5.000514, 5.000224, 5.000093, 5.000038, 5.000018, 
    5.000008,
  // momentumY(5,45, 0-49)
    5, 5.000002, 5.000007, 5.000016, 5.000035, 5.000085, 5.000203, 5.000461, 
    5.001007, 5.002101, 5.004179, 5.007924, 5.014315, 5.024631, 5.040349, 
    5.062917, 5.093406, 5.131166, 5.175416, 5.224458, 5.275883, 5.328215, 
    5.376691, 5.416956, 5.442389, 5.451115, 5.442218, 5.416569, 5.376009, 
    5.327141, 5.274342, 5.222435, 5.173072, 5.128863, 5.091638, 5.062168, 
    5.040212, 5.024796, 5.014577, 5.00817, 5.004367, 5.002228, 5.001084, 
    5.000504, 5.000224, 5.000095, 5.00004, 5.000018, 5.000009, 5.000004,
  // momentumY(5,46, 0-49)
    5, 5, 5.000003, 5.000008, 5.000017, 5.000037, 5.000086, 5.0002, 5.000446, 
    5.000955, 5.001951, 5.0038, 5.007055, 5.012488, 5.021063, 5.033856, 
    5.051858, 5.075415, 5.104631, 5.138946, 5.177042, 5.217485, 5.256517, 
    5.289888, 5.311668, 5.319259, 5.311596, 5.289727, 5.256232, 5.217037, 
    5.176403, 5.138111, 5.10367, 5.074477, 5.051146, 5.033548, 5.021009, 
    5.012557, 5.007162, 5.003898, 5.002025, 5.001004, 5.000476, 5.000216, 
    5.000093, 5.00004, 5.000018, 5.00001, 5.000005, 5,
  // momentumY(5,47, 0-49)
    5, 5, 5, 5.000004, 5.00001, 5.000017, 5.000035, 5.000082, 5.000188, 
    5.000413, 5.000865, 5.001729, 5.003295, 5.005988, 5.010376, 5.017145, 
    5.027009, 5.040486, 5.057955, 5.079401, 5.10426, 5.131539, 5.158699, 
    5.182441, 5.198313, 5.203908, 5.198285, 5.182379, 5.15859, 5.131369, 
    5.104017, 5.079085, 5.057591, 5.040131, 5.026741, 5.017027, 5.010357, 
    5.006016, 5.003337, 5.001766, 5.000893, 5.000431, 5.000199, 5.000088, 
    5.000038, 5.000018, 5.00001, 5.000006, 5.000001, 5,
  // momentumY(5,48, 0-49)
    5, 5, 5, 5, 5.000005, 5.000009, 5.000016, 5.000033, 5.000074, 5.000168, 
    5.00036, 5.000737, 5.001443, 5.002692, 5.004791, 5.008132, 5.013163, 
    5.020295, 5.029888, 5.0421, 5.056754, 5.073282, 5.09015, 5.105158, 
    5.115366, 5.118993, 5.115357, 5.105136, 5.090113, 5.073223, 5.056668, 
    5.041988, 5.029758, 5.020169, 5.013067, 5.00809, 5.004785, 5.002703, 
    5.001458, 5.00075, 5.000369, 5.000174, 5.000078, 5.000034, 5.000016, 
    5.000009, 5.000005, 5.000001, 5, 5,
  // momentumY(5,49, 0-49)
    5, 5, 5, 5, 5, 5.000002, 5.000004, 5.00001, 5.000021, 5.000049, 5.00011, 
    5.000237, 5.000488, 5.000957, 5.001791, 5.003193, 5.005428, 5.008776, 
    5.013537, 5.019944, 5.02806, 5.037715, 5.048037, 5.057581, 5.064183, 
    5.06655, 5.064181, 5.057576, 5.048025, 5.037696, 5.028031, 5.019907, 
    5.013492, 5.008731, 5.005393, 5.003181, 5.001791, 5.000962, 5.000493, 
    5.000242, 5.000113, 5.000051, 5.000022, 5.00001, 5.000005, 5.000002, 5, 
    5, 5, 5,
  // momentumY(6,0, 0-49)
    5.000001, 5.000006, 5.00001, 5.000018, 5.000034, 5.000072, 5.000154, 
    5.000316, 5.000631, 5.001208, 5.002222, 5.003925, 5.006657, 5.010836, 
    5.01693, 5.025394, 5.036568, 5.050474, 5.066961, 5.08557, 5.105506, 
    5.125745, 5.144631, 5.160282, 5.170508, 5.174044, 5.170405, 5.160065, 
    5.144283, 5.12525, 5.104868, 5.084815, 5.066161, 5.049734, 5.036002, 
    5.025083, 5.016811, 5.010836, 5.006715, 5.003999, 5.002289, 5.00126, 
    5.000666, 5.00034, 5.000166, 5.000079, 5.000038, 5.000019, 5.000011, 
    5.000007,
  // momentumY(6,1, 0-49)
    5.000005, 5.00001, 5.000018, 5.000033, 5.00007, 5.000151, 5.00032, 
    5.000653, 5.001278, 5.002406, 5.004348, 5.007544, 5.012561, 5.020073, 
    5.030783, 5.045307, 5.064008, 5.086517, 5.11232, 5.140503, 5.169809, 
    5.198979, 5.225753, 5.247741, 5.261885, 5.266718, 5.261647, 5.247239, 
    5.224946, 5.197832, 5.168324, 5.13874, 5.110439, 5.084771, 5.062673, 
    5.044592, 5.030516, 5.020079, 5.012699, 5.007718, 5.004508, 5.002532, 
    5.001365, 5.000708, 5.000353, 5.00017, 5.00008, 5.000038, 5.000021, 
    5.000012,
  // momentumY(6,2, 0-49)
    5.000009, 5.000016, 5.000031, 5.000069, 5.000152, 5.000327, 5.000679, 
    5.001356, 5.002598, 5.004784, 5.008452, 5.014331, 5.023312, 5.036367, 
    5.054408, 5.078065, 5.107471, 5.141197, 5.177971, 5.216177, 5.254053, 
    5.290477, 5.322897, 5.349, 5.365357, 5.37082, 5.364851, 5.347931, 
    5.321181, 5.288037, 5.250886, 5.212396, 5.173913, 5.137403, 5.104555, 
    5.076529, 5.053838, 5.036386, 5.023619, 5.014725, 5.008818, 5.005071, 
    5.002802, 5.001487, 5.000758, 5.000372, 5.000178, 5.000082, 5.000039, 
    5.000021,
  // momentumY(6,3, 0-49)
    5.000015, 5.000031, 5.000066, 5.000148, 5.000325, 5.000685, 5.001394, 
    5.002722, 5.005103, 5.009176, 5.015826, 5.026171, 5.041471, 5.06295, 
    5.091514, 5.127439, 5.170224, 5.216258, 5.26322, 5.308789, 5.351055, 
    5.389846, 5.422889, 5.44876, 5.464318, 5.469281, 5.463325, 5.446671, 
    5.41954, 5.385091, 5.344875, 5.301375, 5.2552, 5.208684, 5.164347, 
    5.124405, 5.090402, 5.063021, 5.042137, 5.027025, 5.016627, 5.009819, 
    5.005565, 5.003028, 5.001583, 5.000794, 5.000385, 5.00018, 5.000083, 
    5.00004,
  // momentumY(6,4, 0-49)
    5.000029, 5.000062, 5.00014, 5.00031, 5.000668, 5.001381, 5.002748, 
    5.005244, 5.009598, 5.016839, 5.0283, 5.045533, 5.070081, 5.103135, 
    5.145094, 5.195261, 5.252154, 5.308517, 5.361249, 5.407907, 5.447248, 
    5.481152, 5.508186, 5.528504, 5.5398, 5.542978, 5.537997, 5.524723, 
    5.502158, 5.472632, 5.436204, 5.394633, 5.346801, 5.294731, 5.241333, 
    5.189841, 5.143176, 5.103406, 5.07149, 5.047315, 5.029989, 5.018214, 
    5.010605, 5.005923, 5.003174, 5.001634, 5.000808, 5.000386, 5.00018, 
    5.000086,
  // momentumY(6,5, 0-49)
    5.000058, 5.000128, 5.000286, 5.000626, 5.001318, 5.002669, 5.005185, 
    5.009661, 5.017243, 5.029462, 5.048134, 5.075124, 5.1119, 5.158987, 
    5.215483, 5.279093, 5.347617, 5.408614, 5.459496, 5.498811, 5.526948, 
    5.548717, 5.563705, 5.573915, 5.578139, 5.578449, 5.57507, 5.567517, 
    5.553593, 5.534558, 5.508757, 5.477044, 5.435779, 5.385819, 5.329535, 
    5.270462, 5.212655, 5.159855, 5.114769, 5.078687, 5.051541, 5.032279, 
    5.019346, 5.011106, 5.006111, 5.003226, 5.001635, 5.000797, 5.000378, 
    5.000181,
  // momentumY(6,6, 0-49)
    5.000115, 5.000255, 5.000564, 5.001209, 5.002492, 5.00493, 5.009352, 
    5.016989, 5.029522, 5.049008, 5.077607, 5.11707, 5.168053, 5.229499, 
    5.298431, 5.370821, 5.445284, 5.502716, 5.543248, 5.567499, 5.578008, 
    5.582731, 5.581964, 5.579405, 5.574989, 5.571723, 5.570034, 5.569163, 
    5.56598, 5.56068, 5.55012, 5.534544, 5.507586, 5.468422, 5.417926, 
    5.358761, 5.295095, 5.231841, 5.173631, 5.123855, 5.084163, 5.05453, 
    5.033725, 5.019936, 5.011277, 5.006112, 5.003177, 5.001587, 5.000769, 
    5.000376,
  // momentumY(6,7, 0-49)
    5.000226, 5.000491, 5.001064, 5.002233, 5.004501, 5.008698, 5.016093, 
    5.028466, 5.048059, 5.0773, 5.118228, 5.171681, 5.236503, 5.309232, 
    5.384604, 5.457738, 5.530963, 5.576744, 5.600434, 5.605077, 5.595113, 
    5.581197, 5.563703, 5.547695, 5.534246, 5.527015, 5.526596, 5.532055, 
    5.539679, 5.548707, 5.554925, 5.558561, 5.5509, 5.529508, 5.493343, 
    5.443217, 5.382048, 5.31462, 5.246725, 5.183888, 5.130181, 5.087585, 
    5.056075, 5.034219, 5.019936, 5.011107, 5.005926, 5.003036, 5.001507, 
    5.000752,
  // momentumY(6,8, 0-49)
    5.000422, 5.000904, 5.001921, 5.003942, 5.007765, 5.014642, 5.026388, 
    5.045363, 5.074217, 5.115291, 5.169679, 5.236262, 5.311226, 5.388562, 
    5.461514, 5.526134, 5.591987, 5.620574, 5.624623, 5.609064, 5.579417, 
    5.548193, 5.515173, 5.486481, 5.46438, 5.452968, 5.453032, 5.463569, 
    5.480635, 5.502585, 5.524538, 5.547294, 5.560452, 5.560471, 5.544627, 
    5.511597, 5.462111, 5.399347, 5.328711, 5.256863, 5.190205, 5.133425, 
    5.088749, 5.056075, 5.033725, 5.019349, 5.010611, 5.00558, 5.002838, 
    5.001445,
  // momentumY(6,9, 0-49)
    5.000753, 5.001589, 5.003309, 5.006641, 5.012774, 5.023482, 5.041159, 
    5.068617, 5.108491, 5.162234, 5.228955, 5.304729, 5.382974, 5.456024, 
    5.5172, 5.565434, 5.620588, 5.629872, 5.615059, 5.581898, 5.535974, 
    5.490709, 5.444725, 5.404984, 5.375036, 5.359287, 5.358814, 5.372686, 
    5.397056, 5.429439, 5.464555, 5.504181, 5.536883, 5.558599, 5.565522, 
    5.554592, 5.52423, 5.475126, 5.410761, 5.337203, 5.261992, 5.192336, 
    5.133425, 5.087586, 5.054531, 5.032286, 5.018225, 5.009846, 5.005136, 
    5.00267,
  // momentumY(6,10, 0-49)
    5.001282, 5.002665, 5.005434, 5.010663, 5.020015, 5.035825, 5.060974, 
    5.098361, 5.149876, 5.215099, 5.290311, 5.368649, 5.441668, 5.501667, 
    5.54359, 5.570598, 5.614685, 5.605386, 5.574833, 5.52846, 5.471034, 
    5.416002, 5.360381, 5.31177, 5.275041, 5.254829, 5.25267, 5.267902, 
    5.297109, 5.337039, 5.382149, 5.435371, 5.484737, 5.526087, 5.55515, 
    5.567821, 5.560739, 5.532126, 5.482728, 5.416425, 5.34004, 5.261992, 
    5.190205, 5.130182, 5.084167, 5.051551, 5.03001, 5.016677, 5.008926, 
    5.004739,
  // momentumY(6,11, 0-49)
    5.002078, 5.004252, 5.008497, 5.016294, 5.029826, 5.051929, 5.085682, 
    5.133456, 5.195515, 5.268737, 5.346379, 5.41946, 5.479264, 5.519618, 
    5.53792, 5.542086, 5.576544, 5.550974, 5.508726, 5.454051, 5.390294, 
    5.330138, 5.268671, 5.213834, 5.171679, 5.146977, 5.141926, 5.156423, 
    5.187869, 5.232409, 5.284306, 5.34762, 5.410196, 5.467977, 5.516637, 
    5.551656, 5.568658, 5.564036, 5.535913, 5.485223, 5.416424, 5.337204, 
    5.256864, 5.183889, 5.12386, 5.078702, 5.04735, 5.027104, 5.014899, 
    5.008082,
  // momentumY(6,12, 0-49)
    5.003199, 5.006451, 5.012627, 5.023664, 5.042225, 5.071439, 5.11411, 
    5.171338, 5.240982, 5.31694, 5.390095, 5.450813, 5.491652, 5.508848, 
    5.502183, 5.484329, 5.5107, 5.471681, 5.42171, 5.363332, 5.298191, 
    5.237552, 5.174379, 5.116498, 5.070714, 5.04173, 5.032598, 5.044168, 
    5.075143, 5.121388, 5.177038, 5.247113, 5.3195, 5.390254, 5.455167, 
    5.509714, 5.549153, 5.568865, 5.565066, 5.535909, 5.482724, 5.41076, 
    5.328711, 5.246729, 5.17364, 5.114793, 5.071546, 5.042262, 5.023884, 
    5.013244,
  // momentumY(6,13, 0-49)
    5.004665, 5.00928, 5.017808, 5.032618, 5.056721, 5.093204, 5.144015, 
    5.208309, 5.2812, 5.354035, 5.416568, 5.459991, 5.479059, 5.472442, 
    5.441646, 5.404009, 5.422162, 5.372473, 5.318215, 5.260051, 5.197939, 
    5.141232, 5.080792, 5.023685, 4.976696, 4.944057, 4.92978, 4.936145, 
    4.963764, 5.008761, 5.065294, 5.139062, 5.21817, 5.298661, 5.376439, 
    5.447134, 5.506054, 5.548239, 5.568853, 5.564024, 5.532117, 5.475121, 
    5.399345, 5.314625, 5.231855, 5.159892, 5.10349, 5.063205, 5.036771, 
    5.020852,
  // momentumY(6,14, 0-49)
    5.006432, 5.012634, 5.023786, 5.042606, 5.072232, 5.115298, 5.172375, 
    5.240322, 5.311727, 5.376356, 5.424157, 5.448103, 5.445302, 5.416306, 
    5.363493, 5.308928, 5.315402, 5.257618, 5.201933, 5.147207, 5.091923, 
    5.043219, 4.99018, 4.938323, 4.893336, 4.858306, 4.838092, 4.836915, 
    4.85803, 4.898629, 4.953203, 5.027792, 5.110849, 5.19822, 5.285783, 
    5.369319, 5.444354, 5.506011, 5.549108, 5.568622, 5.560715, 5.524216, 
    5.462107, 5.382053, 5.295115, 5.212708, 5.143295, 5.09066, 5.054367, 
    5.031552,
  // momentumY(6,15, 0-49)
    5.008353, 5.01623, 5.03002, 5.052654, 5.087132, 5.135281, 5.196004, 
    5.263953, 5.329874, 5.383046, 5.414553, 5.419429, 5.396732, 5.348141, 
    5.276179, 5.207609, 5.194048, 5.130501, 5.075865, 5.027326, 4.982164, 
    4.945155, 4.904314, 4.862773, 4.823861, 4.788546, 4.762092, 4.751051, 
    4.762189, 4.794866, 4.844478, 4.917047, 5.001487, 5.09321, 5.187871, 
    5.281279, 5.369182, 5.446979, 5.509586, 5.551565, 5.567762, 5.554559, 
    5.511582, 5.443219, 5.358788, 5.270534, 5.190001, 5.124745, 5.077209, 
    5.045891,
  // momentumY(6,16, 0-49)
    5.010181, 5.019599, 5.035693, 5.061436, 5.099479, 5.150658, 5.212265, 
    5.277219, 5.335279, 5.376088, 5.392232, 5.380555, 5.341426, 5.277007, 
    5.189547, 5.10928, 5.061175, 4.993652, 4.942364, 4.902635, 4.870674, 
    4.848741, 4.82494, 4.799216, 4.771264, 4.738774, 4.706534, 4.683522, 
    4.680879, 4.701571, 4.742841, 4.810379, 4.893664, 4.987398, 5.086774, 
    5.187449, 5.285298, 5.376024, 5.45486, 5.516427, 5.555016, 5.565443, 
    5.544588, 5.493336, 5.417953, 5.329622, 5.241532, 5.164762, 5.10537, 
    5.064186,
  // momentumY(6,17, 0-49)
    5.011572, 5.022128, 5.039799, 5.067472, 5.107347, 5.159363, 5.219592, 
    5.279918, 5.329862, 5.35982, 5.363729, 5.339694, 5.288814, 5.213394, 
    5.115401, 5.023416, 4.91982, 4.848852, 4.803052, 4.775018, 4.75953, 
    4.755941, 4.754036, 4.749845, 4.738373, 4.712875, 4.676379, 4.639837, 
    4.619423, 4.623429, 4.652407, 4.711521, 4.790933, 4.884343, 4.986193, 
    5.091783, 5.19697, 5.297701, 5.389572, 5.46752, 5.525795, 5.558423, 
    5.560376, 5.529471, 5.46844, 5.385913, 5.294955, 5.209147, 5.138294, 
    5.086379,
  // momentumY(6,18, 0-49)
    5.012167, 5.023161, 5.04132, 5.069361, 5.109135, 5.160046, 5.217618, 
    5.273468, 5.317338, 5.340284, 5.337028, 5.306277, 5.249497, 5.169226, 
    5.067511, 4.957667, 4.773083, 4.697157, 4.658534, 4.645606, 4.650552, 
    4.668773, 4.693651, 4.71667, 4.727506, 4.714119, 4.676271, 4.625728, 
    4.583766, 4.56583, 4.577911, 4.624625, 4.69708, 4.787639, 4.889681, 
    4.997922, 5.108042, 5.21612, 5.318082, 5.409255, 5.484136, 5.536518, 
    5.560242, 5.550798, 5.507571, 5.435857, 5.34702, 5.255654, 5.174771, 
    5.111942,
  // momentumY(6,19, 0-49)
    5.011673, 5.022164, 5.039426, 5.06602, 5.103715, 5.152024, 5.206848, 
    5.260324, 5.302584, 5.324714, 5.321186, 5.290559, 5.234613, 5.15659, 
    5.058802, 4.913702, 4.622737, 4.538507, 4.507798, 4.513911, 4.544353, 
    4.588445, 4.64507, 4.700685, 4.73955, 4.744065, 4.709301, 4.645968, 
    4.579593, 4.53436, 4.524497, 4.554203, 4.616135, 4.700994, 4.800754, 
    4.909312, 5.022017, 5.134962, 5.244314, 5.345772, 5.434191, 5.503454, 
    5.546865, 5.558331, 5.534452, 5.477069, 5.394795, 5.301735, 5.213065, 
    5.139863,
  // momentumY(6,20, 0-49)
    5.009789, 5.018234, 5.032057, 5.053111, 5.08257, 5.119898, 5.161999, 
    5.20331, 5.237241, 5.258398, 5.264359, 5.256173, 5.237612, 5.213781, 
    5.189564, 0, 4.351584, 4.34895, 4.370693, 4.414233, 4.476791, 4.54938, 
    4.639208, 4.728305, 4.795688, 4.818511, 4.786697, 4.708689, 4.613272, 
    4.53438, 4.497091, 4.504663, 4.552106, 4.628093, 4.722847, 4.829231, 
    4.942132, 5.057541, 5.171772, 5.280826, 5.379914, 5.463161, 5.523698, 
    5.554443, 5.54987, 5.508664, 5.436234, 5.345024, 5.251167, 5.168735,
  // momentumY(6,21, 0-49)
    5.008009, 5.014865, 5.026288, 5.044007, 5.069425, 5.102808, 5.142482, 
    5.184568, 5.223716, 5.254673, 5.273949, 5.280734, 5.276828, 5.265878, 
    5.252289, 0, 4.170659, 4.190443, 4.237646, 4.309671, 4.403232, 4.505134, 
    4.625941, 4.743216, 4.833209, 4.872109, 4.84777, 4.765993, 4.654385, 
    4.551601, 4.492404, 4.478347, 4.510312, 4.576025, 4.664337, 4.767112, 
    4.878688, 4.994842, 5.111915, 5.226116, 5.33296, 5.426864, 5.501005, 
    5.547768, 5.560138, 5.534248, 5.47243, 5.384887, 5.287694, 5.197131,
  // momentumY(6,22, 0-49)
    5.006531, 5.012131, 5.021671, 5.036806, 5.059116, 5.089477, 5.127281, 
    5.16994, 5.2131, 5.25171, 5.281518, 5.300305, 5.308352, 5.308174, 
    5.303796, 0, 4.030805, 4.065196, 4.131796, 4.227709, 4.348972, 4.477757, 
    4.627515, 4.771355, 4.883232, 4.939029, 4.924598, 4.842271, 4.716929, 
    4.590865, 4.509266, 4.470721, 4.484496, 4.53761, 4.617585, 4.715239, 
    4.824254, 4.940064, 5.058887, 5.17696, 5.289956, 5.392478, 5.47778, 
    5.537942, 5.564931, 5.552924, 5.501613, 5.41886, 5.320036, 5.22286,
  // momentumY(6,23, 0-49)
    5.005608, 5.010423, 5.018781, 5.032283, 5.052613, 5.081013, 5.117546, 
    5.160475, 5.206153, 5.249742, 5.28655, 5.313443, 5.329684, 5.337036, 
    5.339309, 0, 3.936208, 3.979444, 4.05963, 4.173486, 4.31631, 4.465572, 
    4.636799, 4.799335, 4.926097, 4.994142, 4.988685, 4.909207, 4.776904, 
    4.635037, 4.536873, 4.476786, 4.473642, 4.514404, 4.585753, 4.677729, 
    4.783483, 4.898127, 5.017705, 5.138398, 5.255899, 5.364881, 5.458617, 
    5.528984, 5.567272, 5.566283, 5.52371, 5.445437, 5.345931, 5.243716,
  // momentumY(6,24, 0-49)
    5.005395, 5.009989, 5.017999, 5.030992, 5.050661, 5.078343, 5.114321, 
    5.157181, 5.203599, 5.248916, 5.288375, 5.318546, 5.338296, 5.349046, 
    5.354481, 0, 3.885182, 3.932935, 4.020948, 4.145664, 4.301788, 4.463101, 
    4.646461, 4.818689, 4.952569, 5.026831, 5.027077, 4.951261, 4.817554, 
    4.668488, 4.561754, 4.487683, 4.472909, 4.504726, 4.569493, 4.656837, 
    4.759587, 4.872656, 4.991975, 5.113683, 5.233487, 5.346098, 5.444815, 
    5.521412, 5.566805, 5.572984, 5.536391, 5.461555, 5.362166, 5.257078,
  // momentumY(6,25, 0-49)
    5.005977, 5.010957, 5.019516, 5.033198, 5.053604, 5.081876, 5.118042, 
    5.160445, 5.205666, 5.249183, 5.286569, 5.314772, 5.332943, 5.342594, 
    5.347287, 0, 3.875384, 3.92374, 4.013379, 4.140702, 4.30019, 4.464015, 
    4.64996, 4.823952, 4.9589, 5.034354, 5.036249, 4.962126, 4.829005, 
    4.67878, 4.570251, 4.491889, 4.473286, 4.501997, 4.564393, 4.650023, 
    4.75163, 4.864066, 4.983222, 5.105221, 5.225766, 5.339579, 5.439962, 
    5.518659, 5.566463, 5.575105, 5.5406, 5.46701, 5.367731, 5.261695,
  // momentumY(6,26, 0-49)
    5.007358, 5.013331, 5.023318, 5.038845, 5.061301, 5.09135, 5.128307, 
    5.169772, 5.211891, 5.250265, 5.281169, 5.302535, 5.31439, 5.318717, 
    5.319005, 0, 3.907399, 3.952108, 4.036621, 4.157588, 4.309739, 4.466147, 
    4.645107, 4.813356, 4.943969, 5.016002, 5.015329, 4.94009, 4.808348, 
    4.662022, 4.557912, 4.485681, 4.471959, 4.5043, 4.569307, 4.656758, 
    4.759554, 4.872642, 4.991968, 5.113681, 5.233484, 5.346098, 5.444815, 
    5.521413, 5.566805, 5.572984, 5.53639, 5.461555, 5.362166, 5.257078,
  // momentumY(6,27, 0-49)
    5.009464, 5.016989, 5.029191, 5.047569, 5.07317, 5.105905, 5.143998, 
    5.18394, 5.221245, 5.251712, 5.272612, 5.283283, 5.285047, 5.280668, 
    5.273688, 0, 3.984281, 4.020194, 4.092436, 4.198112, 4.332588, 4.472099, 
    4.634583, 4.789214, 4.909461, 4.973031, 4.965724, 4.887423, 4.759062, 
    4.622608, 4.529527, 4.472963, 4.471822, 4.513583, 4.585392, 4.677572, 
    4.783415, 4.898097, 5.017692, 5.138393, 5.255897, 5.36488, 5.458617, 
    5.528984, 5.567272, 5.566283, 5.52371, 5.445437, 5.345931, 5.243716,
  // momentumY(6,28, 0-49)
    5.012121, 5.021662, 5.036722, 5.058746, 5.08832, 5.12436, 5.163691, 
    5.201473, 5.232535, 5.253003, 5.261386, 5.258695, 5.247797, 5.232471, 
    5.216447, 0, 4.109945, 4.130611, 4.183319, 4.265604, 4.37358, 4.487952, 
    4.624791, 4.757003, 4.859302, 4.908553, 4.891548, 4.811182, 4.691791, 
    4.573579, 4.499115, 4.465442, 4.481968, 4.536459, 4.617074, 4.715014, 
    4.824155, 4.940021, 5.058867, 5.176952, 5.289953, 5.392476, 5.477779, 
    5.537941, 5.564931, 5.552924, 5.501613, 5.41886, 5.320036, 5.22286,
  // momentumY(6,29, 0-49)
    5.01504, 5.026921, 5.045306, 5.071594, 5.1058, 5.145628, 5.186234, 
    5.221255, 5.244844, 5.253647, 5.247667, 5.229831, 5.204763, 5.177385, 
    5.151611, 0, 4.284205, 4.28185, 4.307784, 4.359859, 4.434813, 4.518023, 
    4.622173, 4.724629, 4.802577, 4.8335, 4.806474, 4.727848, 4.624166, 
    4.531176, 4.480493, 4.472147, 4.507318, 4.574645, 4.663714, 4.766834, 
    4.878564, 4.994786, 5.11189, 5.226105, 5.332955, 5.426862, 5.501004, 
    5.547768, 5.560138, 5.534248, 5.47243, 5.384888, 5.287694, 5.197131,
  // momentumY(6,30, 0-49)
    5.01805, 5.03292, 5.056044, 5.089447, 5.133391, 5.184988, 5.237677, 
    5.28241, 5.310273, 5.315083, 5.294526, 5.249707, 5.183735, 5.100007, 
    5.000019, 4.8457, 4.545903, 4.460265, 4.430046, 4.441324, 4.48198, 
    4.537408, 4.612211, 4.688424, 4.746189, 4.764202, 4.733611, 4.662929, 
    4.579001, 4.51218, 4.48446, 4.498162, 4.54897, 4.626636, 4.722182, 
    4.82893, 4.941996, 5.057481, 5.171744, 5.280814, 5.379909, 5.463158, 
    5.523697, 5.554443, 5.54987, 5.508664, 5.436234, 5.345024, 5.251167, 
    5.168735,
  // momentumY(6,31, 0-49)
    5.019023, 5.03479, 5.059389, 5.094986, 5.141794, 5.196579, 5.252171, 
    5.298905, 5.32757, 5.332101, 5.310494, 5.263934, 5.195178, 5.107091, 
    5.00141, 4.883553, 4.684901, 4.605775, 4.566805, 4.557559, 4.570552, 
    4.598731, 4.639916, 4.681739, 4.709561, 4.707233, 4.671093, 4.611933, 
    4.553517, 4.517052, 4.514324, 4.54877, 4.613411, 4.699682, 4.800136, 
    4.909025, 5.021885, 5.134902, 5.244286, 5.345759, 5.434185, 5.503451, 
    5.546865, 5.558331, 5.534452, 5.477069, 5.394795, 5.301735, 5.213065, 
    5.139863,
  // momentumY(6,32, 0-49)
    5.018395, 5.033809, 5.058214, 5.094069, 5.14203, 5.199332, 5.259036, 
    5.311258, 5.346146, 5.356833, 5.340679, 5.298523, 5.232965, 5.146788, 
    5.041823, 4.942011, 4.822749, 4.747123, 4.69965, 4.673524, 4.664025, 
    4.668962, 4.681037, 4.693107, 4.696065, 4.679071, 4.64244, 4.597218, 
    4.562731, 4.552108, 4.569833, 4.620241, 4.694829, 4.786526, 4.889145, 
    4.997667, 5.107924, 5.216065, 5.318056, 5.409244, 5.484132, 5.536515, 
    5.560241, 5.550798, 5.507571, 5.435857, 5.34702, 5.255654, 5.174771, 
    5.111942,
  // momentumY(6,33, 0-49)
    5.016522, 5.030602, 5.0534, 5.087697, 5.134883, 5.193241, 5.256811, 
    5.316042, 5.360482, 5.382006, 5.376657, 5.344406, 5.287577, 5.209101, 
    5.111249, 5.021931, 4.958303, 4.88466, 4.830286, 4.790932, 4.763344, 
    4.748603, 4.736362, 4.723997, 4.707599, 4.681181, 4.647666, 4.616824, 
    4.603018, 4.612907, 4.64622, 4.708125, 4.789161, 4.883449, 4.985752, 
    5.091572, 5.196871, 5.297654, 5.389551, 5.46751, 5.525791, 5.558421, 
    5.560375, 5.529471, 5.46844, 5.385913, 5.294955, 5.209147, 5.138294, 
    5.086379,
  // momentumY(6,34, 0-49)
    5.013892, 5.025993, 5.046119, 5.077284, 5.121665, 5.178928, 5.244718, 
    5.310551, 5.365828, 5.401097, 5.410602, 5.392849, 5.349452, 5.283387, 
    5.197491, 5.117618, 5.088926, 5.017687, 4.958633, 4.909221, 4.867121, 
    4.835982, 4.804241, 4.772992, 4.742702, 4.71132, 4.683036, 4.66551, 
    4.668421, 4.693704, 4.738229, 4.807829, 4.892317, 4.98671, 5.086431, 
    5.187284, 5.285219, 5.375988, 5.454842, 5.516418, 5.555013, 5.565441, 
    5.544586, 5.493335, 5.417953, 5.329622, 5.241532, 5.164762, 5.10537, 
    5.064186,
  // momentumY(6,35, 0-49)
    5.010988, 5.020812, 5.037631, 5.064511, 5.10425, 5.157928, 5.223202, 
    5.293424, 5.358673, 5.408595, 5.435466, 5.43575, 5.409719, 5.359928, 
    5.289591, 5.220821, 5.212025, 5.144827, 5.083393, 5.026625, 4.973094, 
    4.928782, 4.882309, 4.837645, 4.798489, 4.765621, 4.743443, 4.737309, 
    4.752937, 4.789107, 4.841118, 4.915183, 5.000496, 5.092699, 5.187614, 
    5.281154, 5.369122, 5.446951, 5.509573, 5.55156, 5.56776, 5.554558, 
    5.511581, 5.443218, 5.358788, 5.270534, 5.190001, 5.124745, 5.077209, 
    5.045891,
  // momentumY(6,36, 0-49)
    5.008206, 5.015754, 5.029075, 5.051062, 5.084832, 5.132618, 5.194133, 
    5.265147, 5.33742, 5.400627, 5.445424, 5.465913, 5.46032, 5.430084, 
    5.378282, 5.323157, 5.325123, 5.264044, 5.202501, 5.140908, 5.078958, 
    5.024843, 4.968314, 4.915356, 4.871645, 4.839771, 4.823688, 4.826664, 
    4.851294, 4.894493, 4.950805, 5.026462, 5.110141, 5.197854, 5.285599, 
    5.369229, 5.444311, 5.505991, 5.549098, 5.568619, 5.560713, 5.524215, 
    5.462106, 5.382053, 5.295115, 5.212708, 5.143295, 5.09066, 5.054367, 
    5.031552,
  // momentumY(6,37, 0-49)
    5.005801, 5.011303, 5.021308, 5.038361, 5.065549, 5.105801, 5.160549, 
    5.228139, 5.302862, 5.375661, 5.436546, 5.477478, 5.494156, 5.486094, 
    5.455472, 5.416793, 5.425346, 5.372597, 5.313364, 5.249673, 5.182581, 
    5.122284, 5.060222, 5.003567, 4.958797, 4.929513, 4.918928, 4.928662, 
    4.958955, 5.005849, 5.063618, 5.138137, 5.217677, 5.298407, 5.37631, 
    5.447072, 5.506024, 5.548225, 5.568847, 5.564021, 5.532116, 5.475121, 
    5.399345, 5.314625, 5.231855, 5.159892, 5.10349, 5.063205, 5.036771, 
    5.020852,
  // momentumY(6,38, 0-49)
    5.003891, 5.007699, 5.014834, 5.027377, 5.048105, 5.080132, 5.126007, 
    5.186297, 5.258187, 5.335034, 5.407619, 5.466704, 5.505548, 5.521119, 
    5.513827, 5.494351, 5.508985, 5.466975, 5.412887, 5.350326, 5.281836, 
    5.219258, 5.155951, 5.099565, 5.056434, 5.03064, 5.024622, 5.038822, 
    5.071777, 5.119378, 5.175891, 5.246482, 5.319166, 5.390081, 5.455081, 
    5.509673, 5.549134, 5.568857, 5.565062, 5.535907, 5.482723, 5.41076, 
    5.32871, 5.246728, 5.17364, 5.114793, 5.071546, 5.042262, 5.023884, 
    5.013244,
  // momentumY(6,39, 0-49)
    5.002481, 5.004988, 5.009824, 5.01858, 5.03355, 5.057617, 5.093771, 
    5.144087, 5.20835, 5.282921, 5.360754, 5.432937, 5.491165, 5.529831, 
    5.546874, 5.548873, 5.571401, 5.542856, 5.497346, 5.439801, 5.37418, 
    5.313456, 5.252906, 5.200124, 5.160659, 5.138759, 5.136208, 5.152687, 
    5.185562, 5.231051, 5.283538, 5.347201, 5.409976, 5.467864, 5.516581, 
    5.55163, 5.568645, 5.56403, 5.53591, 5.485222, 5.416424, 5.337203, 
    5.256864, 5.183889, 5.12386, 5.078702, 5.04735, 5.027104, 5.014899, 
    5.008082,
  // momentumY(6,40, 0-49)
    5.001506, 5.003077, 5.006195, 5.012006, 5.022259, 5.039356, 5.066173, 
    5.105471, 5.158852, 5.225492, 5.301316, 5.379313, 5.451182, 5.50957, 
    5.549834, 5.574276, 5.607434, 5.595249, 5.56227, 5.514218, 5.45616, 
    5.401567, 5.34748, 5.301089, 5.266817, 5.248916, 5.24868, 5.265357, 
    5.295565, 5.336142, 5.381646, 5.435097, 5.484591, 5.526011, 5.555113, 
    5.567804, 5.56073, 5.532122, 5.482724, 5.416423, 5.340039, 5.261992, 
    5.190205, 5.130182, 5.084167, 5.051551, 5.03001, 5.016677, 5.008926, 
    5.004739,
  // momentumY(6,41, 0-49)
    5.000872, 5.001811, 5.003726, 5.007394, 5.014062, 5.025565, 5.044321, 
    5.073099, 5.114377, 5.169344, 5.236801, 5.312582, 5.390053, 5.461687, 
    5.521057, 5.566554, 5.612437, 5.619046, 5.602568, 5.568698, 5.523036, 
    5.478834, 5.434624, 5.396982, 5.369114, 5.355171, 5.356116, 5.371006, 
    5.396053, 5.428863, 5.464231, 5.504002, 5.536785, 5.558545, 5.565493, 
    5.554577, 5.524221, 5.475122, 5.410758, 5.337202, 5.261991, 5.192336, 
    5.133424, 5.087586, 5.054531, 5.032286, 5.018225, 5.009846, 5.005136, 
    5.00267,
  // momentumY(6,42, 0-49)
    5.000481, 5.001017, 5.00214, 5.004345, 5.008471, 5.015812, 5.028213, 
    5.048029, 5.077842, 5.119837, 5.174886, 5.241633, 5.316115, 5.392297, 
    5.463521, 5.525497, 5.583997, 5.61024, 5.613234, 5.597641, 5.568791, 
    5.538901, 5.507612, 5.480733, 5.460288, 5.450224, 5.451291, 5.462511, 
    5.480014, 5.502224, 5.524326, 5.547166, 5.560371, 5.560421, 5.544595, 
    5.511576, 5.462096, 5.399337, 5.328705, 5.25686, 5.190202, 5.133424, 
    5.088748, 5.056075, 5.033725, 5.019349, 5.010611, 5.00558, 5.002838, 
    5.001445,
  // momentumY(6,43, 0-49)
    5.000254, 5.000546, 5.001174, 5.002439, 5.00487, 5.009325, 5.017095, 
    5.029969, 5.050164, 5.080025, 5.121449, 5.175093, 5.239628, 5.311485, 
    5.385376, 5.456191, 5.523962, 5.567801, 5.590858, 5.595832, 5.586867, 
    5.574288, 5.558316, 5.543778, 5.53159, 5.525327, 5.525582, 5.531467, 
    5.539334, 5.548489, 5.55477, 5.558441, 5.550801, 5.52943, 5.493284, 
    5.443173, 5.382017, 5.3146, 5.246713, 5.18388, 5.130176, 5.087583, 
    5.056074, 5.034219, 5.019936, 5.011107, 5.005926, 5.003036, 5.001507, 
    5.000752,
  // momentumY(6,44, 0-49)
    5.000128, 5.000281, 5.000617, 5.00131, 5.002675, 5.005249, 5.009875, 
    5.017793, 5.030678, 5.050543, 5.079468, 5.119081, 5.169894, 5.230724, 
    5.298507, 5.369052, 5.439737, 5.495649, 5.53579, 5.560483, 5.571956, 
    5.577868, 5.578365, 5.576972, 5.573505, 5.570918, 5.569647, 5.568985, 
    5.565864, 5.560555, 5.549966, 5.534374, 5.507415, 5.468267, 5.417797, 
    5.358663, 5.295023, 5.231793, 5.1736, 5.123836, 5.084153, 5.054524, 
    5.033722, 5.019935, 5.011277, 5.006111, 5.003177, 5.001587, 5.000769, 
    5.000376,
  // momentumY(6,45, 0-49)
    5.000063, 5.000138, 5.000311, 5.000674, 5.001407, 5.002824, 5.005446, 
    5.010069, 5.017841, 5.03027, 5.049132, 5.07621, 5.112875, 5.159539, 
    5.21521, 5.277477, 5.343553, 5.403429, 5.454043, 5.493758, 5.522719, 
    5.545506, 5.561567, 5.57276, 5.57775, 5.578548, 5.575379, 5.567812, 
    5.55373, 5.5345, 5.508538, 5.476731, 5.435433, 5.385492, 5.329256, 
    5.270243, 5.212493, 5.159744, 5.114697, 5.078644, 5.051517, 5.032265, 
    5.019338, 5.011102, 5.00611, 5.003224, 5.001634, 5.000797, 5.000378, 
    5.000181,
  // momentumY(6,46, 0-49)
    5.000031, 5.000067, 5.00015, 5.000331, 5.000709, 5.001454, 5.002869, 
    5.005435, 5.009881, 5.017223, 5.02877, 5.046025, 5.070468, 5.103213, 
    5.144585, 5.193819, 5.249195, 5.304764, 5.3573, 5.404286, 5.444343, 
    5.479204, 5.507306, 5.528643, 5.540705, 5.544287, 5.539324, 5.525741, 
    5.502674, 5.472641, 5.435821, 5.39402, 5.3461, 5.29405, 5.24074, 
    5.189366, 5.142821, 5.103158, 5.071325, 5.047211, 5.029928, 5.018178, 
    5.010585, 5.005913, 5.00317, 5.001631, 5.000807, 5.000385, 5.000178, 
    5.000086,
  // momentumY(6,47, 0-49)
    5.000016, 5.000032, 5.000071, 5.000156, 5.000339, 5.000712, 5.00144, 
    5.002793, 5.0052, 5.009297, 5.015947, 5.026236, 5.041384, 5.062566, 
    5.090646, 5.125872, 5.167685, 5.213145, 5.259974, 5.305874, 5.348906, 
    5.388846, 5.423281, 5.450551, 5.467137, 5.472547, 5.466381, 5.448959, 
    5.420728, 5.385215, 5.34418, 5.300195, 5.253817, 5.207319, 5.163136, 
    5.123419, 5.089652, 5.062486, 5.041776, 5.026793, 5.016487, 5.009737, 
    5.005519, 5.003005, 5.001571, 5.000789, 5.000381, 5.000178, 5.000082, 
    5.00004,
  // momentumY(6,48, 0-49)
    5.00001, 5.000016, 5.000032, 5.00007, 5.000153, 5.000327, 5.000675, 
    5.00134, 5.002559, 5.004692, 5.008262, 5.013968, 5.022671, 5.035318, 
    5.052807, 5.075786, 5.104437, 5.137691, 5.174414, 5.213105, 5.252073, 
    5.290257, 5.324902, 5.35331, 5.371335, 5.377446, 5.370953, 5.352503, 
    5.323604, 5.288409, 5.249669, 5.210224, 5.171314, 5.134784, 5.102191, 
    5.074564, 5.052313, 5.035273, 5.022853, 5.014224, 5.008505, 5.004887, 
    5.002697, 5.001432, 5.000731, 5.000358, 5.00017, 5.000078, 5.000036, 
    5.000019,
  // momentumY(6,49, 0-49)
    5.000003, 5.000005, 5.00001, 5.000021, 5.000048, 5.000105, 5.000226, 
    5.000469, 5.000938, 5.001801, 5.003329, 5.005904, 5.010058, 5.016455, 
    5.025851, 5.039001, 5.056527, 5.078323, 5.104247, 5.133745, 5.165843, 
    5.199856, 5.232936, 5.261728, 5.280608, 5.287194, 5.280442, 5.261369, 
    5.232347, 5.199001, 5.164706, 5.132356, 5.102732, 5.076899, 5.055445, 
    5.038478, 5.025686, 5.016487, 5.010173, 5.006035, 5.00344, 5.001884, 
    5.000993, 5.000504, 5.000246, 5.000115, 5.000053, 5.000024, 5.000012, 
    5.000007,
  // momentumY(7,0, 0-49)
    5.000065, 5.000127, 5.000259, 5.000518, 5.001007, 5.001891, 5.003428, 
    5.005995, 5.010108, 5.016434, 5.025755, 5.038896, 5.056596, 5.079338, 
    5.107157, 5.139503, 5.175241, 5.211763, 5.247095, 5.279533, 5.307879, 
    5.331899, 5.350907, 5.364714, 5.372608, 5.374767, 5.371186, 5.361848, 
    5.346594, 5.326201, 5.300992, 5.271825, 5.239199, 5.204507, 5.169468, 
    5.135854, 5.105211, 5.078644, 5.05671, 5.039443, 5.026458, 5.017118, 
    5.010684, 5.006434, 5.003739, 5.002098, 5.001138, 5.000597, 5.000308, 
    5.000164,
  // momentumY(7,1, 0-49)
    5.000121, 5.000238, 5.00048, 5.000947, 5.001812, 5.003347, 5.005964, 
    5.010249, 5.016973, 5.027078, 5.041602, 5.061525, 5.087564, 5.119916, 
    5.158052, 5.20067, 5.245986, 5.289452, 5.328742, 5.362245, 5.389309, 
    5.411021, 5.42722, 5.438537, 5.444373, 5.445482, 5.441986, 5.433731, 
    5.419994, 5.40147, 5.377745, 5.349227, 5.315303, 5.277005, 5.236064, 
    5.194644, 5.154975, 5.118989, 5.08803, 5.062733, 5.043062, 5.028478, 
    5.018152, 5.011154, 5.00661, 5.003779, 5.002086, 5.001116, 5.000584, 
    5.000315,
  // momentumY(7,2, 0-49)
    5.000235, 5.000459, 5.00091, 5.001763, 5.003306, 5.005982, 5.010434, 
    5.017533, 5.028368, 5.04416, 5.066104, 5.095097, 5.131435, 5.174539, 
    5.222845, 5.274029, 5.325931, 5.371635, 5.409235, 5.437857, 5.457925, 
    5.47228, 5.481415, 5.48696, 5.488639, 5.487854, 5.484875, 5.479411, 
    5.470135, 5.457471, 5.440103, 5.41785, 5.388554, 5.352391, 5.310528, 
    5.264997, 5.218402, 5.17348, 5.132623, 5.097514, 5.068947, 5.046889, 
    5.030686, 5.019336, 5.011737, 5.006867, 5.003877, 5.00212, 5.001133, 
    5.000619,
  // momentumY(7,3, 0-49)
    5.000447, 5.000865, 5.001686, 5.003202, 5.005878, 5.010405, 5.017734, 
    5.029084, 5.045851, 5.069425, 5.100871, 5.14055, 5.18778, 5.240693, 
    5.296419, 5.351787, 5.405229, 5.447082, 5.476982, 5.495352, 5.503921, 
    5.507381, 5.506683, 5.504385, 5.500591, 5.497306, 5.494962, 5.493176, 
    5.490098, 5.485869, 5.478354, 5.466926, 5.447763, 5.419919, 5.383484, 
    5.339691, 5.290837, 5.239985, 5.190429, 5.145115, 5.106135, 5.074507, 
    5.050228, 5.032541, 5.020276, 5.012163, 5.007035, 5.003933, 5.00215, 
    5.001194,
  // momentumY(7,4, 0-49)
    5.00083, 5.001577, 5.003015, 5.005607, 5.010071, 5.01742, 5.028973, 
    5.046284, 5.070925, 5.104134, 5.146344, 5.196767, 5.253208, 5.312281, 
    5.370041, 5.423226, 5.472451, 5.504696, 5.522296, 5.52714, 5.522073, 
    5.513369, 5.501997, 5.491229, 5.481532, 5.475423, 5.473501, 5.47537, 
    5.478836, 5.483813, 5.487583, 5.489424, 5.484031, 5.469409, 5.444396, 
    5.408932, 5.364272, 5.312967, 5.258545, 5.204911, 5.155597, 5.11315, 
    5.078824, 5.052646, 5.033748, 5.020789, 5.012327, 5.007061, 5.003947, 
    5.002234,
  // momentumY(7,5, 0-49)
    5.00148, 5.002769, 5.005187, 5.009442, 5.016574, 5.027974, 5.045319, 
    5.070355, 5.104497, 5.148292, 5.200894, 5.259817, 5.321171, 5.380404, 
    5.433293, 5.477595, 5.517872, 5.536584, 5.539735, 5.53039, 5.512024, 
    5.492009, 5.470812, 5.452157, 5.436851, 5.427817, 5.425859, 5.430663, 
    5.439898, 5.453335, 5.467922, 5.483245, 5.492867, 5.494058, 5.484577, 
    5.462999, 5.429098, 5.384137, 5.330914, 5.273443, 5.216244, 5.163455, 
    5.118066, 5.081542, 5.053911, 5.034173, 5.020812, 5.012223, 5.006996, 
    5.004036,
  // momentumY(7,6, 0-49)
    5.002537, 5.004672, 5.008571, 5.015256, 5.026145, 5.042995, 5.067703, 
    5.101876, 5.146226, 5.199944, 5.260352, 5.323129, 5.38313, 5.435542, 
    5.476911, 5.507005, 5.535779, 5.539415, 5.528361, 5.50633, 5.476847, 
    5.447856, 5.418829, 5.393694, 5.373574, 5.361693, 5.35911, 5.365716, 
    5.379266, 5.39945, 5.423106, 5.450462, 5.474294, 5.491517, 5.499191, 
    5.494801, 5.476672, 5.444415, 5.399313, 5.344433, 5.284281, 5.224, 
    5.16831, 5.120595, 5.082476, 5.053929, 5.033796, 5.020385, 5.011956, 
    5.007038,
  // momentumY(7,7, 0-49)
    5.004174, 5.007567, 5.013592, 5.023635, 5.039485, 5.063149, 5.09643, 
    5.140269, 5.194015, 5.254954, 5.318458, 5.378851, 5.430717, 5.47008, 
    5.495052, 5.507923, 5.524962, 5.513952, 5.490565, 5.458614, 5.421184, 
    5.386325, 5.352101, 5.322395, 5.298602, 5.284111, 5.280297, 5.287394, 
    5.303493, 5.328266, 5.358603, 5.39561, 5.431551, 5.463284, 5.487547, 
    5.501169, 5.501382, 5.486283, 5.455358, 5.409954, 5.353441, 5.290848, 
    5.227934, 5.169954, 5.120609, 5.081582, 5.052734, 5.032722, 5.019694, 
    5.011834,
  // momentumY(7,8, 0-49)
    5.006591, 5.011756, 5.020663, 5.035065, 5.057024, 5.088521, 5.130782, 
    5.183451, 5.243975, 5.307598, 5.368227, 5.41984, 5.457864, 5.479952, 
    5.486041, 5.480951, 5.487695, 5.463608, 5.430469, 5.391768, 5.349826, 
    5.31244, 5.275925, 5.243874, 5.217835, 5.201171, 5.195599, 5.201853, 
    5.21865, 5.245731, 5.280169, 5.3241, 5.369467, 5.413232, 5.452092, 
    5.482594, 5.501349, 5.505374, 5.492573, 5.462371, 5.416243, 5.357937, 
    5.29305, 5.227945, 5.16834, 5.118135, 5.078969, 5.050519, 5.031245, 
    5.019186,
  // momentumY(7,9, 0-49)
    5.009975, 5.017505, 5.030089, 5.049776, 5.078679, 5.118333, 5.168806, 
    5.227921, 5.291047, 5.351834, 5.403693, 5.44137, 5.461924, 5.464885, 
    5.451752, 5.429615, 5.428216, 5.392973, 5.352669, 5.310205, 5.26699, 
    5.230297, 5.194464, 5.162518, 5.135951, 5.117805, 5.110119, 5.114284, 
    5.12995, 5.157085, 5.193079, 5.241197, 5.293196, 5.346199, 5.396987, 
    5.442087, 5.477869, 5.500757, 5.507577, 5.49611, 5.465787, 5.418324, 
    5.357944, 5.290869, 5.224051, 5.163567, 5.113378, 5.074952, 5.047724, 
    5.029982,
  // momentumY(7,10, 0-49)
    5.01446, 5.02496, 5.041936, 5.067563, 5.103665, 5.150827, 5.207461, 
    5.269351, 5.330144, 5.382782, 5.421267, 5.441902, 5.443639, 5.42762, 
    5.396376, 5.358976, 5.351389, 5.30677, 5.26151, 5.217797, 5.176116, 
    5.143035, 5.110799, 5.081596, 5.056532, 5.03793, 5.028039, 5.029017, 
    5.041786, 5.066779, 5.101882, 5.151564, 5.207518, 5.267011, 5.326935, 
    5.383892, 5.434252, 5.474237, 5.500106, 5.508534, 5.497243, 5.465786, 
    5.416254, 5.353475, 5.284362, 5.216415, 5.155936, 5.106784, 5.070136, 
    5.045145,
  // momentumY(7,11, 0-49)
    5.020058, 5.034059, 5.055914, 5.087668, 5.130448, 5.183438, 5.24315, 
    5.303562, 5.357356, 5.397788, 5.420244, 5.422883, 5.40632, 5.37279, 
    5.325267, 5.274648, 5.261842, 5.209301, 5.160816, 5.117825, 5.079991, 
    5.053068, 5.027225, 5.003541, 4.982328, 4.9647, 4.952865, 4.949788, 
    4.957981, 4.978666, 5.010483, 5.059205, 5.116598, 5.180028, 5.246441, 
    5.312511, 5.374698, 5.429252, 5.472255, 5.499822, 5.50852, 5.4961, 
    5.46238, 5.410001, 5.344549, 5.27369, 5.205394, 5.146018, 5.099126, 
    5.065478,
  // momentumY(7,12, 0-49)
    5.026608, 5.044453, 5.071303, 5.108771, 5.156913, 5.213257, 5.272523, 
    5.327488, 5.37078, 5.396759, 5.402548, 5.387994, 5.354888, 5.305989, 
    5.244225, 5.182299, 5.163545, 5.104256, 5.053853, 5.013101, 4.980991, 
    4.962399, 4.945583, 4.930279, 4.915555, 4.900771, 4.887709, 4.880032, 
    4.882082, 4.896287, 4.922391, 4.967634, 5.024047, 5.089039, 5.159525, 
    5.232173, 5.303509, 5.369896, 5.427476, 5.472199, 5.500046, 5.507537, 
    5.492572, 5.455415, 5.399471, 5.33125, 5.259198, 5.191624, 5.134699, 
    5.091459,
  // momentumY(7,13, 0-49)
    5.033735, 5.05548, 5.086987, 5.129162, 5.180753, 5.237656, 5.293234, 
    5.339825, 5.370763, 5.381915, 5.372065, 5.342326, 5.295123, 5.233254, 
    5.159248, 5.08756, 5.059693, 4.994692, 4.943421, 4.906126, 4.881305, 
    4.872905, 4.867583, 4.863523, 4.858131, 4.848498, 4.835467, 4.823103, 
    4.817653, 4.823181, 4.841021, 4.880143, 4.933115, 4.997382, 5.069714, 
    5.146647, 5.224686, 5.300283, 5.36973, 5.429057, 5.474072, 5.500647, 
    5.505333, 5.486337, 5.44461, 5.384568, 5.313798, 5.241476, 5.176003, 
    5.123024,
  // momentumY(7,14, 0-49)
    5.040861, 5.066214, 5.101596, 5.147029, 5.199935, 5.254867, 5.304424, 
    5.34119, 5.35965, 5.357197, 5.333939, 5.29176, 5.233256, 5.160916, 
    5.076638, 4.99614, 4.952772, 4.88308, 4.831912, 4.799187, 4.783082, 
    4.786512, 4.794985, 4.804932, 4.811784, 4.809976, 4.798848, 4.782353, 
    4.768427, 4.763132, 4.769983, 4.80008, 4.846959, 4.908147, 4.980169, 
    5.059281, 5.141819, 5.224236, 5.302959, 5.374205, 5.433871, 5.477612, 
    5.501223, 5.501401, 5.476885, 5.429611, 5.365265, 5.292587, 5.221282, 
    5.159416,
  // momentumY(7,15, 0-49)
    5.04727, 5.075588, 5.113734, 5.160819, 5.213135, 5.26433, 5.306828, 
    5.333897, 5.341276, 5.327645, 5.294003, 5.242578, 5.175807, 5.095669, 
    5.003297, 4.913842, 4.844732, 4.771318, 4.721283, 4.694343, 4.688432, 
    4.705205, 4.729593, 4.756072, 4.777933, 4.786829, 4.780121, 4.760928, 
    4.738266, 4.720271, 4.713288, 4.731091, 4.768864, 4.824393, 4.893883, 
    4.973128, 5.058129, 5.145205, 5.230836, 5.311429, 5.383089, 5.441543, 
    5.482284, 5.501088, 5.494987, 5.46355, 5.410028, 5.341596, 5.268045, 
    5.19916,
  // momentumY(7,16, 0-49)
    5.052221, 5.082582, 5.122238, 5.169528, 5.219952, 5.266737, 5.302544, 
    5.321485, 5.320392, 5.298859, 5.258375, 5.201202, 5.129457, 5.044556, 
    4.946846, 4.846074, 4.737124, 4.660678, 4.612901, 4.593229, 4.599227, 
    4.630776, 4.672967, 4.718068, 4.757268, 4.779699, 4.780499, 4.761142, 
    4.730637, 4.698801, 4.675304, 4.677201, 4.702387, 4.749299, 4.813816, 
    4.891094, 4.976588, 5.066315, 5.156695, 5.244262, 5.325356, 5.395911, 
    5.45143, 5.487248, 5.499257, 5.485078, 5.445483, 5.385374, 5.313462, 
    5.240213,
  // momentumY(7,17, 0-49)
    5.055084, 5.086399, 5.126359, 5.172816, 5.22089, 5.263784, 5.294598, 
    5.308188, 5.302143, 5.27656, 5.233084, 5.173849, 5.100662, 5.014484, 
    4.914962, 4.796424, 4.630887, 4.5516, 4.507199, 4.496636, 4.516641, 
    4.564325, 4.625845, 4.690973, 4.749099, 4.787496, 4.799221, 4.783396, 
    4.747558, 4.702156, 4.66026, 4.64256, 4.651261, 4.686162, 4.742951, 
    4.81599, 4.899972, 4.990417, 5.083542, 5.175914, 5.264064, 5.344178, 
    5.411934, 5.462564, 5.491307, 5.494365, 5.470315, 5.421548, 5.354854, 
    5.280277,
  // momentumY(7,18, 0-49)
    5.055455, 5.086561, 5.125804, 5.170914, 5.217056, 5.257705, 5.286389, 
    5.298403, 5.291608, 5.26616, 5.223593, 5.165879, 5.094666, 5.010685, 
    4.912883, 4.764289, 4.52522, 4.443193, 4.403152, 4.403866, 4.440429, 
    4.50552, 4.587378, 4.673081, 4.750764, 4.806866, 4.832855, 4.825094, 
    4.788147, 4.731499, 4.671028, 4.630623, 4.61889, 4.638094, 4.684124, 
    4.750472, 4.830854, 4.920098, 5.014065, 5.109241, 5.202271, 5.289577, 
    5.367074, 5.430085, 5.473558, 5.492756, 5.484509, 5.448822, 5.390132, 
    5.31718,
  // momentumY(7,19, 0-49)
    5.053221, 5.082938, 5.120615, 5.164308, 5.209677, 5.250699, 5.281166, 
    5.296271, 5.293453, 5.272348, 5.234126, 5.180676, 5.113756, 5.033909, 
    4.938658, 4.742922, 4.415196, 4.33217, 4.297563, 4.311978, 4.368104, 
    4.45188, 4.554541, 4.660558, 4.75763, 4.832474, 4.875569, 4.880461, 
    4.847667, 4.784114, 4.707324, 4.64267, 4.607326, 4.607371, 4.639596, 
    4.696743, 4.771411, 4.857562, 4.950556, 5.046688, 5.142635, 5.234991, 
    5.319911, 5.392896, 5.448824, 5.4824, 5.489161, 5.467055, 5.418115, 
    5.349228,
  // momentumY(7,20, 0-49)
    5.047519, 5.072911, 5.105344, 5.143125, 5.182673, 5.219129, 5.247638, 
    5.264693, 5.268921, 5.261077, 5.243481, 5.219299, 5.191885, 5.164235, 
    5.138397, 0, 4.114454, 4.114334, 4.146542, 4.211831, 4.306983, 4.4182, 
    4.544752, 4.671088, 4.786033, 4.877743, 4.936459, 4.953573, 4.925799, 
    4.857228, 4.766321, 4.677095, 4.616313, 4.594654, 4.610526, 4.65621, 
    4.723191, 4.804475, 4.894822, 4.990243, 5.087366, 5.182891, 5.273173, 
    5.353907, 5.420018, 5.465905, 5.486187, 5.477157, 5.438637, 5.375458,
  // momentumY(7,21, 0-49)
    5.042906, 5.065928, 5.096264, 5.132921, 5.173195, 5.212954, 5.247571, 
    5.273136, 5.287375, 5.289968, 5.282302, 5.266943, 5.247061, 5.225951, 
    5.206573, 0, 3.960332, 3.978011, 4.033281, 4.12433, 4.2451, 4.375662, 
    4.518851, 4.658369, 4.784651, 4.88853, 4.961393, 4.993842, 4.979385, 
    4.918301, 4.827318, 4.723927, 4.643672, 4.602317, 4.601614, 4.634759, 
    4.692778, 4.76789, 4.85425, 4.947518, 5.044199, 5.141039, 5.234534, 
    5.320562, 5.394155, 5.449563, 5.480793, 5.482881, 5.453789, 5.39637,
  // momentumY(7,22, 0-49)
    5.039219, 5.060489, 5.089365, 5.125412, 5.166588, 5.209273, 5.24895, 
    5.281309, 5.303318, 5.313817, 5.313527, 5.304658, 5.290368, 5.274252, 
    5.259961, 0, 3.835406, 3.868202, 3.942687, 4.05515, 4.197188, 4.343217, 
    4.499814, 4.650155, 4.786009, 4.900363, 4.985329, 5.030774, 5.027747, 
    4.973923, 4.885179, 4.770913, 4.6747, 4.616134, 4.600175, 4.62134, 
    4.670562, 4.739481, 4.821707, 4.912546, 5.008337, 5.105797, 5.201505, 
    5.291459, 5.370781, 5.433647, 5.473652, 5.484908, 5.46392, 5.41185,
  // momentumY(7,23, 0-49)
    5.037024, 5.057234, 5.085255, 5.120999, 5.162849, 5.207517, 5.250546, 
    5.287356, 5.314402, 5.329967, 5.334363, 5.329612, 5.318913, 5.30611, 
    5.295335, 0, 3.75083, 3.794178, 3.882296, 4.009888, 4.166729, 4.322514, 
    4.487185, 4.643687, 4.784962, 4.90581, 4.999001, 5.054017, 5.060269, 
    5.013733, 4.929824, 4.809685, 4.70313, 4.632049, 4.604081, 4.615284, 
    4.656912, 4.720334, 4.798786, 4.887294, 4.982037, 5.079676, 5.176805, 
    5.269478, 5.352865, 5.421083, 5.467453, 5.485446, 5.470525, 5.42257,
  // momentumY(7,24, 0-49)
    5.036716, 5.05663, 5.084397, 5.120026, 5.162042, 5.207297, 5.25141, 
    5.289758, 5.318656, 5.336201, 5.342546, 5.339622, 5.330624, 5.319474, 
    5.310493, 0, 3.710093, 3.758837, 3.854186, 3.98978, 4.154303, 4.314251, 
    4.482039, 4.640524, 4.783451, 4.906882, 5.004126, 5.064573, 5.076762, 
    5.03577, 4.956805, 4.834767, 4.72329, 4.645191, 4.609799, 4.614413, 
    4.65074, 4.710127, 4.785641, 4.872161, 4.96578, 5.063129, 5.160812, 
    5.254916, 5.340633, 5.41205, 5.462324, 5.484553, 5.473571, 5.428463,
  // momentumY(7,25, 0-49)
    5.038471, 5.058876, 5.086976, 5.122606, 5.164133, 5.208367, 5.251034, 
    5.287758, 5.315138, 5.33149, 5.337061, 5.33376, 5.324667, 5.313553, 
    5.304569, 0, 3.712392, 3.76137, 3.857336, 3.993675, 4.158824, 4.318006, 
    4.484923, 4.642324, 4.784227, 4.907133, 5.004549, 5.065886, 5.079467, 
    5.040195, 4.963305, 4.841302, 4.72898, 4.649186, 4.611698, 4.614275, 
    4.648862, 4.706868, 4.781345, 4.867144, 4.960334, 5.057543, 5.155376, 
    5.249931, 5.336409, 5.408885, 5.460465, 5.484119, 5.474478, 5.430358,
  // momentumY(7,26, 0-49)
    5.042217, 5.063863, 5.092844, 5.128556, 5.168951, 5.210625, 5.24946, 
    5.281579, 5.304241, 5.31635, 5.31849, 5.312615, 5.301614, 5.288908, 
    5.278151, 0, 3.755883, 3.80003, 3.890133, 4.020155, 4.179138, 4.333121, 
    4.495686, 4.649438, 4.788105, 4.907743, 5.001677, 5.059398, 5.069646, 
    5.02778, 4.949212, 4.828493, 4.718805, 4.642381, 4.608218, 4.613591, 
    4.650334, 4.709931, 4.785549, 4.872119, 4.96576, 5.06312, 5.160808, 
    5.254914, 5.340632, 5.412049, 5.462324, 5.484553, 5.473571, 5.428463,
  // momentumY(7,27, 0-49)
    5.047648, 5.071205, 5.101556, 5.137453, 5.176219, 5.214128, 5.247229, 
    5.272307, 5.287539, 5.292675, 5.288845, 5.278172, 5.26337, 5.247412, 
    5.233242, 0, 3.837907, 3.872372, 3.950503, 4.067498, 4.213774, 4.358329, 
    4.513062, 4.660518, 4.793601, 4.907108, 4.993864, 5.043576, 5.046104, 
    4.997985, 4.914999, 4.797587, 4.69459, 4.626752, 4.60112, 4.613746, 
    4.65615, 4.719967, 4.798612, 4.887213, 4.981999, 5.079659, 5.176796, 
    5.269475, 5.352864, 5.421082, 5.467452, 5.485446, 5.470524, 5.42257,
  // momentumY(7,28, 0-49)
    5.054279, 5.08032, 5.1125, 5.148775, 5.185695, 5.219107, 5.245215, 
    5.261521, 5.267226, 5.263089, 5.25097, 5.233331, 5.212831, 5.192018, 
    5.172996, 0, 3.95486, 3.975625, 4.036456, 4.134297, 4.261631, 4.392307, 
    4.535101, 4.672795, 4.797129, 4.90109, 4.976916, 5.014869, 5.006731, 
    4.951005, 4.863965, 4.753953, 4.662951, 4.608952, 4.596192, 4.619275, 
    4.669537, 4.738986, 4.821471, 4.912435, 5.008284, 5.105772, 5.201493, 
    5.291453, 5.370779, 5.433645, 5.473652, 5.484908, 5.46392, 5.41185,
  // momentumY(7,29, 0-49)
    5.061519, 5.090569, 5.125088, 5.162135, 5.197347, 5.22602, 5.244443, 
    5.250815, 5.245413, 5.230116, 5.207698, 5.181172, 5.153317, 5.126302, 
    5.101217, 0, 4.100039, 4.105047, 4.144559, 4.218102, 4.320959, 4.433148, 
    4.559563, 4.683653, 4.795854, 4.887011, 4.948723, 4.97219, 4.951942, 
    4.889277, 4.801144, 4.70358, 4.629909, 4.594042, 4.597061, 4.6324, 
    4.6916, 4.767314, 4.853972, 4.947385, 5.044137, 5.141009, 5.23452, 
    5.320555, 5.394152, 5.449561, 5.480793, 5.482881, 5.453789, 5.396369,
  // momentumY(7,30, 0-49)
    5.069942, 5.104444, 5.145037, 5.188226, 5.228665, 5.260446, 5.278681, 
    5.280539, 5.265384, 5.23421, 5.188872, 5.131349, 5.06307, 4.983942, 
    4.890614, 4.694397, 4.378685, 4.306954, 4.281877, 4.30549, 4.370964, 
    4.459809, 4.568273, 4.679267, 4.780853, 4.860884, 4.909776, 4.919673, 
    4.888474, 4.82117, 4.735869, 4.654694, 4.601761, 4.586124, 4.605887, 
    4.653808, 4.721985, 4.803879, 4.89453, 4.990101, 5.087297, 5.182858, 
    5.273158, 5.353899, 5.420014, 5.465903, 5.486187, 5.477157, 5.438637, 
    5.375458,
  // momentumY(7,31, 0-49)
    5.073872, 5.110393, 5.153061, 5.197888, 5.238931, 5.269813, 5.28551, 
    5.283435, 5.26344, 5.227028, 5.17638, 5.113566, 5.040033, 4.956133, 
    4.860312, 4.711382, 4.476999, 4.403505, 4.371749, 4.381316, 4.427418, 
    4.499416, 4.589086, 4.681817, 4.765648, 4.827684, 4.859194, 4.855018, 
    4.817186, 4.75356, 4.681082, 4.623222, 4.59458, 4.599795, 4.6354, 
    4.694525, 4.770272, 4.856986, 4.950268, 5.046546, 5.142564, 5.234956, 
    5.319895, 5.392888, 5.448821, 5.482398, 5.48916, 5.467055, 5.418115, 
    5.349227,
  // momentumY(7,32, 0-49)
    5.074563, 5.111968, 5.156186, 5.203183, 5.24673, 5.279979, 5.297396, 
    5.296023, 5.275575, 5.23764, 5.184599, 5.118748, 5.041742, 4.954269, 
    4.855663, 4.736937, 4.571723, 4.498174, 4.459996, 4.456672, 4.485158, 
    4.540483, 4.610906, 4.684608, 4.750361, 4.79529, 4.81181, 4.797491, 
    4.758013, 4.70317, 4.647774, 4.613843, 4.608014, 4.631615, 4.680494, 
    4.748522, 4.829835, 4.919573, 5.013799, 5.109106, 5.202204, 5.289543, 
    5.367058, 5.430077, 5.473555, 5.492754, 5.484507, 5.448821, 5.390131, 
    5.31718,
  // momentumY(7,33, 0-49)
    5.072055, 5.109157, 5.154137, 5.203316, 5.250513, 5.288494, 5.311002, 
    5.31429, 5.297483, 5.261912, 5.210007, 5.14432, 5.066876, 4.978845, 
    4.880323, 4.778907, 4.66792, 4.594558, 4.550687, 4.536237, 4.549191, 
    4.588276, 4.639575, 4.693966, 4.741624, 4.770691, 4.775239, 4.755387, 
    4.719284, 4.677091, 4.640542, 4.628673, 4.642346, 4.680838, 4.739939, 
    4.814349, 4.8991, 4.989961, 5.083307, 5.175795, 5.264003, 5.344147, 
    5.411918, 5.462556, 5.491303, 5.494362, 5.470314, 5.421547, 5.354854, 
    5.280277,
  // momentumY(7,34, 0-49)
    5.066685, 5.102252, 5.146866, 5.197575, 5.248649, 5.292713, 5.322759, 
    5.333969, 5.324487, 5.295034, 5.247876, 5.185752, 5.11112, 5.025746, 
    4.930516, 4.839296, 4.766814, 4.694075, 4.645786, 4.622183, 4.62171, 
    4.645421, 4.67846, 4.714131, 4.744484, 4.759594, 4.755527, 4.734432, 
    4.705405, 4.677551, 4.65919, 4.666082, 4.695303, 4.745059, 4.811397, 
    4.889759, 4.975869, 5.065935, 5.156497, 5.244161, 5.325305, 5.395886, 
    5.451417, 5.487242, 5.499254, 5.485077, 5.445483, 5.385374, 5.313462, 
    5.240213,
  // momentumY(7,35, 0-49)
    5.059091, 5.091941, 5.134801, 5.18574, 5.23992, 5.290249, 5.329171, 
    5.350695, 5.351656, 5.331776, 5.292833, 5.237574, 5.16882, 5.088939, 
    4.999584, 4.915709, 4.867932, 4.796804, 4.745568, 4.71463, 4.70265, 
    4.712214, 4.728501, 4.746943, 4.761694, 4.765309, 4.755863, 4.73676, 
    4.716686, 4.702873, 4.700494, 4.722412, 4.763369, 4.821098, 4.89199, 
    4.972076, 5.057559, 5.144899, 5.230677, 5.311346, 5.383048, 5.441524, 
    5.482273, 5.501082, 5.494984, 5.463549, 5.410028, 5.341596, 5.268045, 
    5.19916,
  // momentumY(7,36, 0-49)
    5.050116, 5.079262, 5.118917, 5.168323, 5.223925, 5.279467, 5.327296, 
    5.360398, 5.374112, 5.366771, 5.339256, 5.293997, 5.233984, 5.162076, 
    5.080613, 5.003589, 4.970191, 4.901921, 4.849092, 4.81234, 4.790542, 
    4.787408, 4.788884, 4.792263, 4.793777, 4.788606, 4.776517, 4.761394, 
    4.750595, 4.749277, 4.760054, 4.793442, 4.842779, 4.90564, 4.978724, 
    5.058472, 5.141376, 5.223999, 5.302834, 5.37414, 5.433838, 5.477597, 
    5.501214, 5.501397, 5.476884, 5.429609, 5.365265, 5.292587, 5.221282, 
    5.159416,
  // momentumY(7,37, 0-49)
    5.040674, 5.065457, 5.100637, 5.146596, 5.201307, 5.259878, 5.315217, 
    5.359754, 5.387404, 5.394824, 5.381534, 5.34921, 5.300679, 5.239072, 
    5.167283, 5.097776, 5.072126, 5.007897, 4.954634, 4.913358, 4.883272, 
    4.869039, 4.857895, 4.848771, 4.839742, 4.828416, 4.815767, 4.805543, 
    4.803319, 4.812391, 4.833456, 4.87515, 4.92999, 4.995509, 5.06863, 
    5.146039, 5.224351, 5.300103, 5.369635, 5.429007, 5.474048, 5.500636, 
    5.505328, 5.486333, 5.444608, 5.384567, 5.313798, 5.241476, 5.176003, 
    5.123024,
  // momentumY(7,38, 0-49)
    5.031587, 5.051754, 5.081593, 5.122414, 5.173713, 5.232343, 5.292474, 
    5.346719, 5.387997, 5.411265, 5.414304, 5.39752, 5.363111, 5.314147, 
    5.253855, 5.193147, 5.17178, 5.112633, 5.059998, 5.015416, 4.978568, 
    4.954986, 4.933573, 4.914676, 4.897844, 4.882706, 4.870935, 4.86574, 
    4.870833, 4.888049, 4.916724, 4.963934, 5.021742, 5.087658, 5.158724, 
    5.231721, 5.303259, 5.369761, 5.427405, 5.472163, 5.500027, 5.507529, 
    5.492567, 5.455412, 5.39947, 5.33125, 5.259198, 5.191624, 5.134699, 
    5.091459,
  // momentumY(7,39, 0-49)
    5.023478, 5.03917, 5.063326, 5.09785, 5.143517, 5.198998, 5.260269, 
    5.32098, 5.373845, 5.412485, 5.432821, 5.433532, 5.415639, 5.38168, 
    5.334877, 5.284673, 5.266556, 5.213517, 5.162659, 5.11611, 5.074186, 
    5.043216, 5.01401, 4.988095, 4.966056, 4.949053, 4.939028, 4.938462, 
    4.949347, 4.97249, 5.0063, 5.056495, 5.114914, 5.179015, 5.245848, 
    5.312171, 5.374506, 5.429146, 5.472199, 5.499791, 5.508503, 5.496091, 
    5.462376, 5.409999, 5.344549, 5.273689, 5.205394, 5.146018, 5.099126, 
    5.065478,
  // momentumY(7,40, 0-49)
    5.01671, 5.028383, 5.047037, 5.074806, 5.113331, 5.162851, 5.22134, 
    5.284199, 5.344914, 5.396571, 5.433529, 5.452536, 5.452931, 5.436152, 
    5.404949, 5.367265, 5.35313, 5.307418, 5.259766, 5.2129, 5.167883, 
    5.131764, 5.097353, 5.067103, 5.04221, 5.024868, 5.016986, 5.020291, 
    5.035318, 5.062237, 5.098837, 5.149593, 5.206281, 5.266251, 5.326477, 
    5.383618, 5.434089, 5.474142, 5.500051, 5.508503, 5.497226, 5.465776, 
    5.416249, 5.353471, 5.28436, 5.216414, 5.155935, 5.106784, 5.070136, 
    5.045145,
  // momentumY(7,41, 0-49)
    5.011393, 5.019699, 5.033443, 5.054687, 5.08547, 5.127131, 5.179427, 
    5.239829, 5.303455, 5.363914, 5.414792, 5.451157, 5.470404, 5.472347, 
    5.458686, 5.435668, 5.427438, 5.390626, 5.348041, 5.302955, 5.257243, 
    5.218533, 5.181604, 5.149585, 5.123898, 5.107349, 5.101637, 5.107809, 
    5.125257, 5.153823, 5.190883, 5.239744, 5.292246, 5.345578, 5.396583, 
    5.44182, 5.477694, 5.500643, 5.507504, 5.496064, 5.465759, 5.418307, 
    5.357935, 5.290864, 5.224049, 5.163566, 5.113376, 5.074951, 5.047723, 
    5.029982,
  // momentumY(7,42, 0-49)
    5.007448, 5.013103, 5.022773, 5.03824, 5.061559, 5.094617, 5.138445, 
    5.192428, 5.253744, 5.317492, 5.377594, 5.428209, 5.465016, 5.485915, 
    5.491031, 5.484582, 5.484806, 5.458848, 5.423669, 5.382972, 5.339408, 
    5.300989, 5.264325, 5.232959, 5.208259, 5.193301, 5.189502, 5.197357, 
    5.215441, 5.243477, 5.278582, 5.322964, 5.368637, 5.412613, 5.451626, 
    5.482244, 5.501094, 5.50519, 5.492446, 5.462286, 5.416188, 5.357902, 
    5.293029, 5.227933, 5.168333, 5.118133, 5.078968, 5.050518, 5.031245, 
    5.019185,
  // momentumY(7,43, 0-49)
    5.004671, 5.00836, 5.014862, 5.025596, 5.042367, 5.06715, 5.101645, 
    5.146619, 5.201205, 5.262506, 5.325803, 5.385471, 5.436242, 5.474329, 
    5.498009, 5.509168, 5.520347, 5.507353, 5.482279, 5.449014, 5.41083, 
    5.375861, 5.342307, 5.313881, 5.291713, 5.278893, 5.276544, 5.284764, 
    5.301612, 5.326838, 5.35743, 5.394591, 5.430645, 5.462481, 5.486856, 
    5.500595, 5.500926, 5.485937, 5.455106, 5.409778, 5.353324, 5.290773, 
    5.22789, 5.169929, 5.120594, 5.081575, 5.05273, 5.03272, 5.019693, 
    5.011834,
  // momentumY(7,44, 0-49)
    5.002813, 5.005119, 5.009302, 5.016413, 5.027887, 5.045482, 5.071043, 
    5.106079, 5.151144, 5.205262, 5.265625, 5.327862, 5.386883, 5.437991, 
    5.477863, 5.506032, 5.529777, 5.531497, 5.519186, 5.496544, 5.467158, 
    5.438933, 5.411334, 5.388013, 5.36974, 5.359428, 5.357933, 5.365097, 
    5.378753, 5.398783, 5.422194, 5.449341, 5.473051, 5.490255, 5.498004, 
    5.493757, 5.475805, 5.443734, 5.398806, 5.344073, 5.284039, 5.223843, 
    5.168211, 5.120537, 5.082442, 5.053911, 5.033787, 5.020379, 5.011954, 
    5.007036,
  // momentumY(7,45, 0-49)
    5.001627, 5.00301, 5.005588, 5.010087, 5.017568, 5.029425, 5.047313, 
    5.072919, 5.10756, 5.151648, 5.204203, 5.262649, 5.32308, 5.380993, 
    5.432267, 5.474555, 5.510695, 5.527712, 5.530097, 5.520863, 5.503451, 
    5.485116, 5.466168, 5.449955, 5.436787, 5.429237, 5.42793, 5.432586, 
    5.441073, 5.453529, 5.467171, 5.481771, 5.49093, 5.491922, 5.482465, 
    5.461075, 5.427461, 5.382823, 5.329916, 5.272722, 5.215748, 5.163129, 
    5.11786, 5.081418, 5.053839, 5.034134, 5.020792, 5.012212, 5.00699, 
    5.004033,
  // momentumY(7,46, 0-49)
    5.000904, 5.001698, 5.003219, 5.005941, 5.01059, 5.018181, 5.030026, 
    5.047634, 5.072513, 5.105799, 5.147814, 5.197673, 5.25313, 5.310821, 
    5.366889, 5.418075, 5.464053, 5.494967, 5.512374, 5.518117, 5.514961, 
    5.509031, 5.500986, 5.493574, 5.486524, 5.481907, 5.480128, 5.480912, 
    5.48242, 5.485212, 5.486995, 5.487328, 5.480935, 5.465807, 5.440713, 
    5.405491, 5.361278, 5.310514, 5.256648, 5.203514, 5.154617, 5.112494, 
    5.078404, 5.052387, 5.033595, 5.020703, 5.01228, 5.007036, 5.003934, 
    5.002227,
  // momentumY(7,47, 0-49)
    5.000479, 5.000916, 5.001769, 5.003335, 5.006079, 5.010685, 5.018091, 
    5.029477, 5.046185, 5.069523, 5.100471, 5.139313, 5.185328, 5.236683, 
    5.29062, 5.344086, 5.395159, 5.436237, 5.466683, 5.48693, 5.498612, 
    5.506318, 5.510494, 5.51297, 5.512695, 5.511067, 5.508265, 5.504123, 
    5.497348, 5.489172, 5.47811, 5.463986, 5.442956, 5.414068, 5.377319, 
    5.333785, 5.285583, 5.235593, 5.186958, 5.142507, 5.104268, 5.07323, 
    5.049392, 5.032015, 5.019961, 5.011981, 5.006932, 5.003879, 5.00212, 
    5.001179,
  // momentumY(7,48, 0-49)
    5.000237, 5.00046, 5.000906, 5.001745, 5.003255, 5.005858, 5.010167, 
    5.017009, 5.027408, 5.04252, 5.063472, 5.091123, 5.125785, 5.16698, 
    5.213346, 5.262811, 5.313305, 5.359091, 5.398305, 5.430139, 5.45493, 
    5.475578, 5.491802, 5.50423, 5.510761, 5.511994, 5.507837, 5.49834, 
    5.482945, 5.46386, 5.440705, 5.414022, 5.381519, 5.343398, 5.300726, 
    5.255343, 5.209594, 5.165942, 5.126526, 5.092831, 5.06552, 5.044494, 
    5.029083, 5.018308, 5.011105, 5.006493, 5.003665, 5.002002, 5.00107, 
    5.000583,
  // momentumY(7,49, 0-49)
    5.000078, 5.000158, 5.000323, 5.000648, 5.001265, 5.002378, 5.004317, 
    5.007565, 5.012781, 5.020815, 5.032668, 5.049388, 5.071904, 5.100811, 
    5.136148, 5.177304, 5.223419, 5.26947, 5.313471, 5.353898, 5.39002, 
    5.424407, 5.454918, 5.480593, 5.49589, 5.500593, 5.494115, 5.476953, 
    5.449314, 5.416775, 5.380487, 5.34278, 5.30167, 5.258408, 5.214767, 
    5.172745, 5.1342, 5.100561, 5.072627, 5.050539, 5.033884, 5.021892, 
    5.013636, 5.008191, 5.004746, 5.002652, 5.001432, 5.00075, 5.000383, 
    5.000201,
  // momentumY(8,0, 0-49)
    5.001369, 5.00236, 5.004135, 5.007111, 5.011874, 5.019187, 5.02997, 
    5.045208, 5.065813, 5.092411, 5.125103, 5.163265, 5.205472, 5.249606, 
    5.293155, 5.333694, 5.369721, 5.397316, 5.416229, 5.42692, 5.430637, 
    5.429839, 5.425939, 5.420931, 5.415915, 5.412307, 5.410614, 5.410615, 
    5.41119, 5.411488, 5.409767, 5.404738, 5.39423, 5.377171, 5.353137, 
    5.322467, 5.286308, 5.246513, 5.205389, 5.165338, 5.128472, 5.096318, 
    5.069674, 5.048647, 5.032804, 5.021383, 5.013495, 5.008281, 5.005001, 
    5.003084,
  // momentumY(8,1, 0-49)
    5.002229, 5.003803, 5.006566, 5.011106, 5.018226, 5.028921, 5.044301, 
    5.065442, 5.093146, 5.127659, 5.168413, 5.213895, 5.261753, 5.309123, 
    5.353121, 5.391528, 5.424201, 5.445468, 5.456513, 5.458668, 5.453891, 
    5.445782, 5.435674, 5.425931, 5.417472, 5.412071, 5.410341, 5.412109, 
    5.416037, 5.421542, 5.426564, 5.429821, 5.428074, 5.419613, 5.403261, 
    5.378569, 5.345982, 5.306887, 5.263489, 5.218513, 5.174774, 5.134702, 
    5.100015, 5.071559, 5.049369, 5.032875, 5.021171, 5.013241, 5.008139, 
    5.005085,
  // momentumY(8,2, 0-49)
    5.003713, 5.006243, 5.010573, 5.017516, 5.028118, 5.043579, 5.065092, 
    5.093582, 5.12938, 5.171907, 5.219525, 5.269629, 5.319023, 5.3645, 
    5.403409, 5.434417, 5.459604, 5.47129, 5.472511, 5.465329, 5.452096, 
    5.437172, 5.421472, 5.407487, 5.395916, 5.388781, 5.386798, 5.389922, 
    5.39677, 5.407083, 5.418703, 5.430604, 5.438771, 5.441057, 5.435635, 
    5.421216, 5.397282, 5.364281, 5.323711, 5.278013, 5.230247, 5.183597, 
    5.140839, 5.103923, 5.073798, 5.050491, 5.033351, 5.021364, 5.013425, 
    5.008539,
  // momentumY(8,3, 0-49)
    5.006076, 5.010056, 5.016683, 5.027022, 5.042336, 5.063916, 5.092799, 
    5.129389, 5.173098, 5.222139, 5.273632, 5.324032, 5.36979, 5.408006, 
    5.436888, 5.456504, 5.471837, 5.472431, 5.463517, 5.447612, 5.427128, 
    5.40682, 5.386859, 5.369648, 5.355633, 5.346969, 5.344492, 5.348353, 
    5.357283, 5.371386, 5.388593, 5.408371, 5.426187, 5.439701, 5.446662, 
    5.445097, 5.433551, 5.411355, 5.378881, 5.337667, 5.290347, 5.24031, 
    5.191145, 5.146004, 5.107107, 5.075537, 5.051323, 5.033752, 5.021726, 
    5.014085,
  // momentumY(8,4, 0-49)
    5.009637, 5.015692, 5.025481, 5.040294, 5.061502, 5.09025, 5.127049, 
    5.171336, 5.221224, 5.273581, 5.324505, 5.370071, 5.407087, 5.433594, 
    5.449055, 5.455122, 5.460109, 5.449643, 5.431532, 5.408463, 5.382619, 
    5.358882, 5.336395, 5.317299, 5.301744, 5.291907, 5.288743, 5.292657, 
    5.302639, 5.319189, 5.340461, 5.366611, 5.392787, 5.416655, 5.435787, 
    5.447778, 5.450466, 5.442185, 5.42209, 5.39045, 5.348847, 5.300132, 
    5.24806, 5.196651, 5.149448, 5.108942, 5.07633, 5.051642, 5.034104, 
    5.022564,
  // momentumY(8,5, 0-49)
    5.01475, 5.023616, 5.037497, 5.057807, 5.085801, 5.12212, 5.166306, 
    5.216456, 5.269265, 5.320505, 5.365861, 5.401783, 5.426079, 5.438101, 
    5.438597, 5.430701, 5.42629, 5.4058, 5.380095, 5.351824, 5.322756, 
    5.297715, 5.274599, 5.255134, 5.239125, 5.228632, 5.224696, 5.228026, 
    5.237998, 5.255537, 5.279135, 5.309788, 5.342454, 5.374955, 5.404862, 
    5.429592, 5.446565, 5.453413, 5.448264, 5.430104, 5.399138, 5.357038, 
    5.306925, 5.252957, 5.199602, 5.15078, 5.109215, 5.07619, 5.051716, 
    5.034968,
  // momentumY(8,6, 0-49)
    5.021751, 5.034218, 5.053062, 5.079626, 5.114713, 5.158042, 5.207815, 
    5.260664, 5.312117, 5.35747, 5.39277, 5.415498, 5.424806, 5.421356, 
    5.406937, 5.385913, 5.373868, 5.3448, 5.313278, 5.281764, 5.251529, 
    5.227237, 5.205383, 5.187147, 5.171925, 5.161469, 5.156841, 5.159067, 
    5.168033, 5.185125, 5.209272, 5.242446, 5.279513, 5.318528, 5.357177, 
    5.392874, 5.422873, 5.444416, 5.454944, 5.452408, 5.435674, 5.404944, 
    5.362053, 5.310448, 5.254735, 5.199829, 5.15, 5.108155, 5.075609, 5.052327,
  // momentumY(8,7, 0-49)
    5.03087, 5.047679, 5.07213, 5.105202, 5.146861, 5.19554, 5.247961, 
    5.299513, 5.345158, 5.38049, 5.402569, 5.410242, 5.403994, 5.385534, 
    5.357308, 5.324667, 5.306974, 5.270771, 5.235045, 5.202008, 5.172415, 
    5.150715, 5.131906, 5.116521, 5.103456, 5.093926, 5.088892, 5.089666, 
    5.096759, 5.112054, 5.135026, 5.168761, 5.208121, 5.251438, 5.296572, 
    5.341026, 5.38205, 5.416742, 5.442186, 5.45566, 5.454984, 5.438967, 
    5.407883, 5.363819, 5.310629, 5.253408, 5.197519, 5.147527, 5.106443, 
    5.075536,
  // momentumY(8,8, 0-49)
    5.042141, 5.063857, 5.094147, 5.13329, 5.180078, 5.231492, 5.282947, 
    5.329145, 5.365218, 5.387711, 5.395039, 5.387403, 5.366355, 5.334259, 
    5.293848, 5.251297, 5.229727, 5.187588, 5.148976, 5.115803, 5.088339, 
    5.070806, 5.056664, 5.045733, 5.036299, 5.028781, 5.023865, 5.023066, 
    5.027584, 5.039847, 5.060001, 5.092403, 5.132013, 5.177479, 5.226856, 
    5.277767, 5.32753, 5.373251, 5.411896, 5.440407, 5.455941, 5.456232, 
    5.440107, 5.408016, 5.362398, 5.307615, 5.249297, 5.193226, 5.14417, 
    5.105097,
  // momentumY(8,9, 0-49)
    5.055322, 5.08219, 5.118004, 5.162039, 5.21173, 5.262723, 5.309602, 
    5.347069, 5.371074, 5.379469, 5.372033, 5.35006, 5.315778, 5.271844, 
    5.22097, 5.170115, 5.145872, 5.098701, 5.058197, 5.025952, 5.0018, 
    4.989735, 4.981704, 4.976761, 4.972498, 4.968266, 4.964252, 4.962024, 
    4.963476, 4.971612, 4.987387, 5.016612, 5.05449, 5.100041, 5.151529, 
    5.206686, 5.262909, 5.317366, 5.367041, 5.408783, 5.439424, 5.456029, 
    5.456311, 5.439203, 5.405454, 5.357993, 5.301782, 5.243008, 5.187781, 
    5.140861,
  // momentumY(8,10, 0-49)
    5.069841, 5.101693, 5.142138, 5.189268, 5.239218, 5.286673, 5.326009, 
    5.352551, 5.363453, 5.357918, 5.336849, 5.30226, 5.256696, 5.202795, 
    5.143048, 5.085224, 5.058656, 5.007109, 4.965445, 4.934928, 4.915015, 
    4.909478, 4.908812, 4.911294, 4.913756, 4.914239, 4.912184, 4.908985, 
    4.907153, 4.910244, 4.920147, 4.944366, 4.97854, 5.022159, 5.07372, 
    5.131052, 5.191589, 5.252552, 5.310984, 5.363772, 5.407672, 5.439425, 
    5.456047, 5.4553, 5.436343, 5.400368, 5.35093, 5.293661, 5.235225, 
    5.181823,
  // momentumY(8,11, 0-49)
    5.084838, 5.121063, 5.164775, 5.212887, 5.260504, 5.301888, 5.331789, 
    5.346568, 5.34467, 5.326456, 5.293612, 5.248514, 5.193708, 5.13161, 
    5.064352, 5.000533, 4.970798, 4.915408, 4.873148, 4.844985, 4.83006, 
    4.831906, 4.839677, 4.850883, 4.861561, 4.868284, 4.869509, 4.866175, 
    4.861197, 4.858579, 4.861226, 4.878594, 4.907023, 4.946648, 4.996276, 
    5.053806, 5.116663, 5.182054, 5.247064, 5.308654, 5.363636, 5.408683, 
    5.44047, 5.45601, 5.453212, 5.431593, 5.392934, 5.341518, 5.283602, 
    5.226091,
  // momentumY(8,12, 0-49)
    5.099267, 5.138888, 5.184268, 5.231308, 5.274516, 5.308251, 5.328059, 
    5.331479, 5.318122, 5.289199, 5.246833, 5.19346, 5.131418, 5.062748, 
    4.989133, 4.919843, 4.884488, 4.825829, 4.783488, 4.758223, 4.748928, 
    4.758839, 4.775925, 4.796943, 4.817178, 4.831673, 4.837736, 4.835538, 
    4.828052, 4.819459, 4.813668, 4.822335, 4.842855, 4.876289, 4.92189, 
    4.977654, 5.040928, 5.108822, 5.178389, 5.246644, 5.310491, 5.366675, 
    5.411796, 5.442484, 5.455814, 5.449941, 5.424872, 5.383087, 5.32959, 
    5.271071,
  // momentumY(8,13, 0-49)
    5.112081, 5.153917, 5.199409, 5.243758, 5.281303, 5.306915, 5.317125, 
    5.310584, 5.287816, 5.250561, 5.201094, 5.141697, 5.07436, 5.000659, 
    4.921747, 4.846888, 4.801401, 4.740222, 4.698379, 4.676562, 4.673483, 
    4.691962, 4.719002, 4.750622, 4.781459, 4.80514, 4.817774, 4.818466, 
    4.809773, 4.795585, 4.780596, 4.77881, 4.789131, 4.813954, 4.853247, 
    4.905177, 4.966969, 5.035536, 5.107794, 5.180731, 5.25133, 5.316455, 
    5.372781, 5.41683, 5.445218, 5.455135, 5.445074, 5.415627, 5.37001, 
    5.313847,
  // momentumY(8,14, 0-49)
    5.122416, 5.165294, 5.209671, 5.250387, 5.28198, 5.300036, 5.302077, 
    5.287667, 5.25795, 5.214927, 5.160814, 5.097618, 5.026911, 4.949761, 
    4.8667, 4.785186, 4.722669, 4.659978, 4.619365, 4.601606, 4.605288, 
    4.632604, 4.669907, 4.712483, 4.754512, 4.788497, 4.809477, 4.815284, 
    4.807504, 4.789055, 4.764913, 4.75128, 4.749103, 4.762674, 4.793109, 
    4.838937, 4.897255, 4.964674, 5.037851, 5.11364, 5.18903, 5.260995, 
    5.326344, 5.381658, 5.423375, 5.448099, 5.453174, 5.437504, 5.402347, 
    5.351675,
  // momentumY(8,15, 0-49)
    5.129766, 5.172712, 5.215269, 5.252206, 5.278469, 5.290407, 5.286373, 
    5.266594, 5.232567, 5.18635, 5.129982, 5.065152, 4.993019, 4.914148, 
    4.828405, 4.73751, 4.64882, 4.585863, 4.547379, 4.534361, 4.545287, 
    4.581367, 4.628794, 4.682116, 4.735318, 4.780255, 4.811194, 4.824649, 
    4.820728, 4.800571, 4.768612, 4.74255, 4.725894, 4.725502, 4.744281, 
    4.781486, 4.83417, 4.898561, 4.970917, 5.047832, 5.126202, 5.203052, 
    5.275322, 5.339731, 5.392716, 5.430585, 5.449921, 5.448276, 5.425073, 
    5.382407,
  // momentumY(8,16, 0-49)
    5.134052, 5.176439, 5.217067, 5.250836, 5.273164, 5.281045, 5.27343, 
    5.250941, 5.215213, 5.16822, 5.111789, 5.047322, 4.975654, 4.896925, 
    4.81037, 4.704902, 4.579583, 4.517775, 4.48243, 4.474857, 4.49339, 
    4.537728, 4.59462, 4.65787, 4.721575, 4.777524, 4.819635, 4.843246, 
    4.846655, 4.828532, 4.791764, 4.754059, 4.721835, 4.705099, 4.70937, 
    4.735244, 4.779961, 4.839344, 4.909132, 4.985513, 5.065176, 5.145107, 
    5.222342, 5.293738, 5.355831, 5.404837, 5.436883, 5.448555, 5.437765, 
    5.404779,
  // momentumY(8,17, 0-49)
    5.13558, 5.177178, 5.216339, 5.248187, 5.268536, 5.274807, 5.266268, 
    5.243672, 5.208608, 5.162899, 5.108179, 5.045659, 4.975985, 4.899038, 
    4.813493, 4.685416, 4.513347, 4.454445, 4.423234, 4.421718, 4.448077, 
    4.499756, 4.565007, 4.636907, 4.70996, 4.776448, 4.830373, 4.866174, 
    4.880282, 4.868591, 4.831599, 4.784774, 4.737452, 4.702971, 4.690291, 
    4.702183, 4.736541, 4.78889, 4.854359, 4.928604, 5.007979, 5.08934, 
    5.169746, 5.246167, 5.315263, 5.37328, 5.416127, 5.43977, 5.440993, 
    5.418493,
  // momentumY(8,18, 0-49)
    5.134904, 5.175833, 5.214426, 5.246045, 5.266733, 5.274041, 5.267223, 
    5.246889, 5.214422, 5.171445, 5.119457, 5.059613, 4.99252, 4.917845, 
    4.833514, 4.673349, 4.446044, 4.392892, 4.366827, 4.371818, 4.406159, 
    4.46414, 4.53652, 4.615712, 4.696862, 4.773158, 4.838974, 4.888155, 
    4.915483, 4.914273, 4.88238, 4.830496, 4.7705, 4.718554, 4.687547, 
    4.683339, 4.705169, 4.748554, 4.808033, 4.878636, 4.956275, 5.037578, 
    5.119546, 5.199218, 5.273369, 5.338331, 5.389959, 5.423878, 5.43611, 
    5.42413,
  // momentumY(8,19, 0-49)
    5.132595, 5.173156, 5.21232, 5.245671, 5.269256, 5.280378, 5.277858, 
    5.261819, 5.23324, 5.193517, 5.144123, 5.086297, 5.020607, 4.946133, 
    4.858912, 4.659686, 4.369835, 4.327592, 4.308208, 4.320153, 4.362873, 
    4.426592, 4.505294, 4.590879, 4.679287, 4.764817, 4.84228, 4.905135, 
    4.946831, 4.958759, 4.936626, 4.884299, 4.815693, 4.74858, 4.699572, 
    4.678265, 4.686046, 4.71891, 4.770968, 4.836618, 4.91126, 4.991214, 
    5.073359, 5.154741, 5.232225, 5.30225, 5.360712, 5.4031, 5.424982, 
    5.422957,
  // momentumY(8,20, 0-49)
    5.126199, 5.16312, 5.199585, 5.231456, 5.255075, 5.268044, 5.269554, 
    5.260229, 5.241733, 5.216325, 5.186499, 5.154742, 5.123319, 5.093983, 
    5.067405, 0, 4.110707, 4.123703, 4.162252, 4.22343, 4.302578, 4.387699, 
    4.480834, 4.576489, 4.673163, 4.767192, 4.854263, 4.927924, 4.980938, 
    5.003913, 4.991771, 4.940973, 4.867107, 4.788014, 4.72289, 4.684924, 
    4.678152, 4.699588, 4.743227, 4.802933, 4.873587, 4.951164, 5.032368, 
    5.114204, 5.193589, 5.267064, 5.330619, 5.379736, 5.409759, 5.416706,
  // momentumY(8,21, 0-49)
    5.123293, 5.160292, 5.19839, 5.233569, 5.261959, 5.280674, 5.288291, 
    5.284894, 5.271763, 5.25098, 5.225037, 5.196559, 5.168098, 5.141923, 
    5.119676, 0, 4.030297, 4.047019, 4.093606, 4.164876, 4.254046, 4.343937, 
    4.441362, 4.540665, 4.641256, 4.74086, 4.835884, 4.920084, 4.985749, 
    5.023064, 5.026696, 4.98524, 4.915319, 4.832731, 4.757448, 4.705839, 
    4.685367, 4.695097, 4.729599, 4.782505, 4.848262, 4.922476, 5.001632, 
    5.082644, 5.162446, 5.237658, 5.304375, 5.358139, 5.394198, 5.408191,
  // momentumY(8,22, 0-49)
    5.121522, 5.158882, 5.19856, 5.236558, 5.268754, 5.291821, 5.30385, 
    5.304541, 5.29497, 5.277183, 5.253765, 5.227507, 5.201188, 5.177412, 
    5.158434, 0, 3.962537, 3.984438, 4.038232, 4.117738, 4.215069, 4.308348, 
    4.409274, 4.511858, 4.616008, 4.720365, 4.821665, 4.913651, 4.988194, 
    5.035557, 5.051208, 5.016985, 4.95165, 4.868662, 4.787441, 4.726087, 
    4.694775, 4.694649, 4.721154, 4.767963, 4.829233, 4.900268, 4.97734, 
    5.057264, 5.136958, 5.2131, 5.281876, 5.338915, 5.379454, 5.398909,
  // momentumY(8,23, 0-49)
    5.120916, 5.158588, 5.199337, 5.239162, 5.273767, 5.299524, 5.314222, 
    5.31733, 5.309831, 5.293787, 5.271873, 5.247006, 5.222109, 5.199984, 
    5.183231, 0, 3.917093, 3.943388, 4.002137, 4.086914, 4.189435, 4.283938, 
    4.386425, 4.49054, 4.59648, 4.703573, 4.808774, 4.905783, 4.986151, 
    5.040359, 5.064946, 5.036311, 4.975649, 4.894337, 4.810658, 4.743364, 
    4.704498, 4.696982, 4.71723, 4.759143, 4.816749, 4.885137, 4.960407, 
    5.039274, 5.118623, 5.195158, 5.265129, 5.324236, 5.367732, 5.390903,
  // momentumY(8,24, 0-49)
    5.121484, 5.15919, 5.200179, 5.240473, 5.275757, 5.302342, 5.317935, 
    5.321938, 5.315293, 5.30006, 5.278937, 5.254865, 5.230805, 5.209631, 
    5.194072, 0, 3.898081, 3.926662, 3.987599, 4.074533, 4.179204, 4.273223, 
    4.375597, 4.479658, 4.58575, 4.69365, 4.800478, 4.89992, 4.983319, 
    5.04135, 5.071414, 5.046269, 4.989053, 4.909707, 4.825484, 4.755218, 
    4.711973, 4.699844, 4.715989, 4.754571, 4.8096, 4.876063, 4.949962, 
    5.027952, 5.106898, 5.183519, 5.254107, 5.31441, 5.359709, 5.385231,
  // momentumY(8,25, 0-49)
    5.12319, 5.160546, 5.200797, 5.240048, 5.274151, 5.299625, 5.314344, 
    5.317798, 5.31093, 5.295742, 5.274842, 5.251086, 5.227356, 5.206459, 
    5.191058, 0, 3.905595, 3.934001, 3.99451, 4.080811, 4.184822, 4.277218, 
    4.378278, 4.481149, 4.586186, 4.693312, 4.799687, 4.89899, 4.982497, 
    5.040989, 5.072271, 5.047817, 4.991623, 4.913149, 4.829183, 4.758409, 
    4.714091, 4.70067, 4.715574, 4.753094, 4.807269, 4.873075, 4.946495, 
    5.024164, 5.102949, 5.179572, 5.250342, 5.311027, 5.356915, 5.383218,
  // momentumY(8,26, 0-49)
    5.125965, 5.16261, 5.201203, 5.237979, 5.269135, 5.291635, 5.303749, 
    5.305204, 5.296997, 5.28103, 5.259737, 5.235774, 5.211836, 5.190529, 
    5.174261, 0, 3.937386, 3.963501, 4.021425, 4.104737, 4.20558, 4.295581, 
    4.394385, 4.495152, 4.598157, 4.703125, 4.807133, 4.903847, 4.984638, 
    5.040278, 5.0684, 5.04177, 4.983876, 4.904703, 4.821317, 4.752176, 
    4.709991, 4.698662, 4.715331, 4.75422, 4.809419, 4.87597, 4.949917, 
    5.027929, 5.106887, 5.183514, 5.254105, 5.314409, 5.359708, 5.385231,
  // momentumY(8,27, 0-49)
    5.129717, 5.165435, 5.201689, 5.23486, 5.261594, 5.279465, 5.287314, 
    5.285252, 5.274403, 5.256595, 5.234052, 5.209174, 5.184377, 5.16194, 
    5.143804, 0, 3.989284, 4.01185, 4.065571, 4.143941, 4.239443, 4.326462, 
    4.422174, 4.519982, 4.619985, 4.72141, 4.821146, 4.912863, 4.98817, 
    5.037752, 5.058598, 5.027196, 4.965382, 4.884583, 4.802653, 4.737598, 
    4.700779, 4.694783, 4.716008, 4.758492, 4.81641, 4.884964, 4.96032, 
    5.03923, 5.118601, 5.195146, 5.265124, 5.324234, 5.36773, 5.390903,
  // momentumY(8,28, 0-49)
    5.134365, 5.169187, 5.202791, 5.231663, 5.252913, 5.264796, 5.266833, 
    5.25964, 5.244601, 5.223562, 5.198596, 5.171845, 5.145388, 5.121049, 
    5.100052, 0, 4.056873, 4.075941, 4.124346, 4.195992, 4.284093, 4.367258, 
    4.458745, 4.55243, 4.648153, 4.744445, 4.837958, 4.922404, 4.989758, 
    5.030591, 5.041007, 5.003144, 4.936561, 4.854705, 4.776264, 4.7182, 
    4.689766, 4.691714, 4.719532, 4.767098, 4.828782, 4.900036, 4.977222, 
    5.057204, 5.136929, 5.213084, 5.281867, 5.338911, 5.379453, 5.398908,
  // momentumY(8,29, 0-49)
    5.139871, 5.174164, 5.205247, 5.229603, 5.244735, 5.249564, 5.244349, 
    5.230343, 5.209353, 5.183419, 5.154596, 5.124834, 5.095839, 5.068839, 
    5.043989, 0, 4.134919, 4.152247, 4.194923, 4.258248, 4.336938, 4.414831, 
    4.500596, 4.588754, 4.67878, 4.768302, 4.853632, 4.928486, 4.985303, 
    5.014688, 5.012098, 4.966738, 4.896005, 4.815494, 4.744064, 4.696627, 
    4.679617, 4.691761, 4.727758, 4.781523, 4.847747, 4.922211, 5.001495, 
    5.082574, 5.16241, 5.23764, 5.304365, 5.358133, 5.394195, 5.408189,
  // momentumY(8,30, 0-49)
    5.149293, 5.187366, 5.220729, 5.245617, 5.259345, 5.260664, 5.249608, 
    5.227057, 5.194283, 5.152627, 5.103288, 5.047123, 4.984291, 4.913467, 
    4.830404, 4.635087, 4.366791, 4.33845, 4.330659, 4.350416, 4.397135, 
    4.457949, 4.533136, 4.614896, 4.700094, 4.78401, 4.861721, 4.926516, 
    4.971288, 4.987126, 4.969789, 4.916682, 4.843794, 4.76844, 4.708371, 
    4.675247, 4.67223, 4.696182, 4.74135, 4.801925, 4.873054, 4.950885, 
    5.032222, 5.114128, 5.19355, 5.267044, 5.330608, 5.37973, 5.409755, 
    5.416704,
  // momentumY(8,31, 0-49)
    5.154108, 5.192601, 5.225134, 5.247748, 5.25784, 5.254495, 5.238242, 
    5.21049, 5.172945, 5.127208, 5.074561, 5.015869, 4.951433, 4.880641, 
    4.801196, 4.644937, 4.432422, 4.392949, 4.379121, 4.393623, 4.43407, 
    4.491832, 4.56249, 4.638905, 4.717442, 4.792549, 4.859183, 4.911111, 
    4.942367, 4.945229, 4.916481, 4.861229, 4.793419, 4.729975, 4.685867, 
    4.669163, 4.680465, 4.715677, 4.769167, 4.835639, 4.910736, 4.990936, 
    5.073214, 5.154664, 5.232185, 5.30223, 5.360701, 5.403094, 5.424978, 
    5.422956,
  // momentumY(8,32, 0-49)
    5.157407, 5.197023, 5.230282, 5.252917, 5.262111, 5.256892, 5.237898, 
    5.206759, 5.165463, 5.115866, 5.059437, 4.997152, 4.929425, 4.855934, 
    4.775219, 4.651386, 4.489683, 4.443143, 4.423618, 4.431955, 4.465497, 
    4.519353, 4.584921, 4.655719, 4.727498, 4.793783, 4.849238, 4.888139, 
    4.905953, 4.896959, 4.860013, 4.806783, 4.748804, 4.70111, 4.675007, 
    4.67511, 4.700132, 4.745621, 4.806382, 4.877728, 4.955783, 5.037313, 
    5.119405, 5.199143, 5.273329, 5.33831, 5.389947, 5.423872, 5.436106, 
    5.424129,
  // momentumY(8,33, 0-49)
    5.158516, 5.199754, 5.23505, 5.259749, 5.270575, 5.266178, 5.24701, 
    5.214706, 5.171402, 5.119178, 5.05975, 4.994316, 4.923507, 4.847308, 
    4.764863, 4.663693, 4.545833, 4.494422, 4.469296, 4.470886, 4.496832, 
    4.54519, 4.604345, 4.668429, 4.732591, 4.78956, 4.833763, 4.860198, 
    4.866086, 4.848289, 4.808124, 4.76158, 4.717298, 4.687345, 4.679305, 
    4.695044, 4.732172, 4.786329, 4.852901, 4.927793, 5.007535, 5.089099, 
    5.169616, 5.246097, 5.315227, 5.37326, 5.416117, 5.439764, 5.44099, 
    5.418491,
  // momentumY(8,34, 0-49)
    5.156674, 5.199654, 5.237898, 5.26634, 5.281066, 5.280095, 5.263408, 
    5.232435, 5.189331, 5.136365, 5.075525, 5.008317, 4.935713, 4.858127, 
    4.77535, 4.688264, 4.605028, 4.550157, 4.519898, 4.514716, 4.532631, 
    4.573838, 4.625031, 4.68093, 4.736253, 4.78332, 4.816595, 4.832085, 
    4.828914, 4.806611, 4.768563, 4.732501, 4.703937, 4.691649, 4.700083, 
    4.72925, 4.776286, 4.837176, 4.907887, 4.984814, 5.064787, 5.144894, 
    5.222227, 5.293676, 5.355797, 5.404819, 5.436873, 5.448549, 5.437762, 
    5.404777,
  // momentumY(8,35, 0-49)
    5.151281, 5.195655, 5.237204, 5.270538, 5.291034, 5.29586, 5.284276, 
    5.257265, 5.216847, 5.165399, 5.10517, 5.038023, 4.965342, 4.888039, 
    4.806555, 4.727874, 4.66922, 4.612257, 4.577751, 4.566242, 4.576077, 
    4.608909, 4.650864, 4.69726, 4.742668, 4.779547, 4.802795, 4.809654, 
    4.800983, 4.778551, 4.746922, 4.72342, 4.710607, 4.714301, 4.736648, 
    4.776581, 4.831155, 4.89677, 4.969879, 5.047243, 5.125873, 5.202868, 
    5.275223, 5.339676, 5.392687, 5.430571, 5.449914, 5.448271, 5.425071, 
    5.382406,
  // momentumY(8,36, 0-49)
    5.142104, 5.187049, 5.231609, 5.270293, 5.297827, 5.310411, 5.306343, 
    5.285905, 5.250766, 5.203276, 5.145887, 5.080808, 5.009852, 4.934427, 
    4.85556, 4.782229, 4.739129, 4.681488, 4.643786, 4.626654, 4.628716, 
    4.652565, 4.684572, 4.720676, 4.75562, 4.782554, 4.797193, 4.798059, 
    4.787327, 4.768233, 4.745573, 4.734941, 4.736442, 4.753576, 4.786968, 
    4.834998, 4.894826, 4.963222, 5.037002, 5.113153, 5.188756, 5.260842, 
    5.326259, 5.381612, 5.423351, 5.448085, 5.453167, 5.4375, 5.402345, 
    5.351675,
  // momentumY(8,37, 0-49)
    5.129393, 5.173698, 5.220318, 5.263993, 5.299031, 5.320687, 5.326133, 
    5.314678, 5.287379, 5.246348, 5.194114, 5.133163, 5.065706, 4.993609, 
    4.918402, 4.849136, 4.814672, 4.757637, 4.717738, 4.695762, 4.690593, 
    4.705426, 4.727391, 4.753076, 4.777669, 4.795451, 4.803186, 4.800547, 
    4.790458, 4.776838, 4.763995, 4.765265, 4.778885, 4.806695, 4.848376, 
    4.902049, 4.965028, 5.034365, 5.107103, 5.18033, 5.251101, 5.316327, 
    5.372707, 5.41679, 5.445196, 5.455124, 5.445068, 5.415625, 5.370009, 
    5.313847,
  // momentumY(8,38, 0-49)
    5.113876, 5.156118, 5.203286, 5.250753, 5.292802, 5.323964, 5.340252, 
    5.339784, 5.322693, 5.290582, 5.245847, 5.191123, 5.128939, 5.06156, 
    4.990949, 4.92551, 4.895123, 4.839703, 4.798448, 4.772382, 4.760661, 
    4.766866, 4.779205, 4.794943, 4.809895, 4.819722, 4.822293, 4.81818, 
    4.810492, 4.803233, 4.799835, 4.811351, 4.83469, 4.870549, 4.918038, 
    4.975163, 5.039362, 5.107861, 5.17781, 5.2463, 5.31029, 5.36656, 
    5.411729, 5.442446, 5.455794, 5.449931, 5.424867, 5.383084, 5.329588, 
    5.27107,
  // momentumY(8,39, 0-49)
    5.096656, 5.135428, 5.181291, 5.230628, 5.278194, 5.318223, 5.345743, 
    5.35758, 5.352668, 5.331766, 5.29685, 5.250499, 5.195425, 5.134211, 
    5.069193, 5.00797, 4.979156, 4.926097, 4.884192, 4.854754, 4.837235, 
    4.835485, 4.838983, 4.845691, 4.852136, 4.855419, 4.85442, 4.850298, 
    4.845923, 4.844999, 4.849974, 4.869821, 4.900551, 4.94209, 4.99318, 
    5.051761, 5.115341, 5.181213, 5.246534, 5.308325, 5.363435, 5.408561, 
    5.440397, 5.455967, 5.453187, 5.43158, 5.392928, 5.341514, 5.283599, 
    5.22609,
  // momentumY(8,40, 0-49)
    5.079001, 5.113148, 5.155824, 5.20466, 5.255383, 5.302495, 5.340465, 
    5.364939, 5.373489, 5.365705, 5.342792, 5.306976, 5.260952, 5.2075, 
    5.149253, 5.093055, 5.064897, 5.0148, 4.972912, 4.940837, 4.918354, 
    4.909531, 4.905233, 4.904131, 4.903456, 4.901661, 4.898442, 4.895254, 
    4.894445, 4.899253, 4.911187, 4.93741, 4.973363, 5.018431, 5.071098, 
    5.129232, 5.190343, 5.251703, 5.310411, 5.363389, 5.407419, 5.439262, 
    5.455943, 5.455236, 5.436306, 5.400346, 5.350918, 5.293653, 5.235221, 
    5.181822,
  // momentumY(8,41, 0-49)
    5.062121, 5.090923, 5.128824, 5.174737, 5.225716, 5.277128, 5.323496, 
    5.359679, 5.381943, 5.388488, 5.379393, 5.356171, 5.321213, 5.27729, 
    5.227234, 5.177218, 5.149961, 5.103456, 5.062327, 5.028457, 5.001982, 
    4.98717, 4.976339, 4.968845, 4.962564, 4.957095, 4.952728, 4.950969, 
    4.953513, 4.963099, 4.980418, 5.011087, 5.050213, 5.096777, 5.149055, 
    5.204819, 5.261506, 5.316321, 5.366274, 5.40823, 5.439034, 5.455762, 
    5.456133, 5.439089, 5.405383, 5.35795, 5.301758, 5.242993, 5.187772, 
    5.140857,
  // momentumY(8,42, 0-49)
    5.046977, 5.07022, 5.102299, 5.143245, 5.191529, 5.243844, 5.29543, 
    5.341003, 5.375879, 5.396879, 5.402698, 5.393766, 5.371802, 5.339299, 
    5.299088, 5.256725, 5.231469, 5.189376, 5.149957, 5.115338, 5.086065, 
    5.066585, 5.050688, 5.038368, 5.028037, 5.02018, 5.015453, 5.015247, 
    5.020588, 5.033757, 5.054786, 5.087964, 5.128242, 5.174273, 5.224139, 
    5.275482, 5.32564, 5.371724, 5.410694, 5.439491, 5.455265, 5.455751, 
    5.439777, 5.407797, 5.36226, 5.307529, 5.249246, 5.193198, 5.144154, 
    5.105088,
  // momentumY(8,43, 0-49)
    5.034163, 5.052107, 5.077977, 5.1126, 5.155713, 5.205489, 5.25843, 
    5.309834, 5.354713, 5.388844, 5.409515, 5.415804, 5.408386, 5.389111, 
    5.360541, 5.327561, 5.306041, 5.269506, 5.233062, 5.199059, 5.168477, 
    5.145934, 5.126657, 5.111196, 5.098354, 5.089241, 5.084676, 5.085835, 
    5.093141, 5.108504, 5.131452, 5.165137, 5.204473, 5.247838, 5.293118, 
    5.337825, 5.379192, 5.41429, 5.440164, 5.454059, 5.453766, 5.438076, 
    5.407258, 5.363396, 5.310354, 5.253236, 5.197416, 5.147466, 5.106408, 
    5.075515,
  // momentumY(8,44, 0-49)
    5.023893, 5.037152, 5.057038, 5.08481, 5.121122, 5.165492, 5.215907, 
    5.268845, 5.319784, 5.364102, 5.398016, 5.419214, 5.427063, 5.422406, 
    5.407182, 5.385447, 5.369846, 5.3404, 5.308588, 5.276946, 5.246899, 
    5.223215, 5.202463, 5.185639, 5.171791, 5.162381, 5.15825, 5.160318, 
    5.168521, 5.184505, 5.207436, 5.239498, 5.275653, 5.314039, 5.352384, 
    5.388091, 5.418369, 5.440388, 5.451512, 5.449613, 5.433495, 5.403317, 
    5.360887, 5.309646, 5.254205, 5.199492, 5.149795, 5.108033, 5.075538, 
    5.052284,
  // momentumY(8,45, 0-49)
    5.016068, 5.025445, 5.040023, 5.06117, 5.090047, 5.127151, 5.171838, 
    5.22204, 5.274341, 5.324514, 5.368355, 5.402508, 5.425014, 5.435463, 
    5.434813, 5.426049, 5.418765, 5.398278, 5.373139, 5.345995, 5.318683, 
    5.296079, 5.275944, 5.259601, 5.246169, 5.237257, 5.233617, 5.23592, 
    5.243749, 5.258614, 5.279437, 5.307597, 5.338169, 5.369109, 5.398049, 
    5.4224, 5.439507, 5.446893, 5.442554, 5.425341, 5.395344, 5.354149, 
    5.304817, 5.251482, 5.198609, 5.150136, 5.108815, 5.075948, 5.051572, 
    5.034879,
  // momentumY(8,46, 0-49)
    5.010371, 5.016713, 5.026895, 5.042174, 5.063859, 5.092983, 5.129908, 
    5.173916, 5.222999, 5.273985, 5.323053, 5.366474, 5.401325, 5.425965, 
    5.440145, 5.44553, 5.448809, 5.439283, 5.423095, 5.402858, 5.380724, 
    5.361625, 5.344312, 5.33029, 5.318596, 5.310812, 5.307542, 5.309251, 
    5.315293, 5.327178, 5.343702, 5.365603, 5.388121, 5.409129, 5.4263, 
    5.437255, 5.439753, 5.431987, 5.41292, 5.382617, 5.342471, 5.295172, 
    5.244368, 5.194016, 5.147643, 5.107752, 5.075573, 5.051174, 5.03382, 
    5.022387,
  // momentumY(8,47, 0-49)
    5.006379, 5.010458, 5.017199, 5.027631, 5.042955, 5.064367, 5.092776, 
    5.128459, 5.170724, 5.217763, 5.2668, 5.314528, 5.357748, 5.393965, 
    5.421778, 5.441412, 5.456867, 5.46001, 5.454927, 5.44398, 5.429455, 
    5.416289, 5.403948, 5.393989, 5.385193, 5.379011, 5.375869, 5.37608, 
    5.378881, 5.385936, 5.396016, 5.409431, 5.421616, 5.430514, 5.434071, 
    5.430398, 5.418005, 5.396079, 5.364757, 5.325294, 5.280035, 5.23211, 
    5.184909, 5.141459, 5.10393, 5.073397, 5.049934, 5.032877, 5.021182, 
    5.013739,
  // momentumY(8,48, 0-49)
    5.003644, 5.006086, 5.010241, 5.016864, 5.02692, 5.041507, 5.061704, 
    5.088339, 5.121694, 5.161249, 5.20556, 5.252367, 5.298956, 5.342635, 
    5.381233, 5.413701, 5.441738, 5.458355, 5.465828, 5.466006, 5.46107, 
    5.455938, 5.450424, 5.446013, 5.441033, 5.436764, 5.433451, 5.431307, 
    5.42953, 5.430123, 5.431936, 5.435133, 5.435347, 5.430807, 5.42, 
    5.401847, 5.375895, 5.342507, 5.302944, 5.259302, 5.21424, 5.17055, 
    5.13068, 5.096348, 5.068379, 5.046762, 5.030877, 5.019772, 5.012416, 
    5.007883,
  // momentumY(8,49, 0-49)
    5.001472, 5.002565, 5.00451, 5.007768, 5.012981, 5.020984, 5.032765, 
    5.049376, 5.071753, 5.100489, 5.135601, 5.176348, 5.22122, 5.268123, 
    5.314735, 5.359285, 5.403051, 5.435205, 5.457379, 5.470873, 5.477746, 
    5.48514, 5.4914, 5.497845, 5.49962, 5.498258, 5.49363, 5.486034, 
    5.474223, 5.463232, 5.452115, 5.442515, 5.428285, 5.40822, 5.38172, 
    5.348891, 5.31062, 5.268536, 5.22482, 5.181884, 5.141978, 5.106841, 
    5.077487, 5.054176, 5.036537, 5.023789, 5.01498, 5.009157, 5.005493, 
    5.003342,
  // momentumY(9,0, 0-49)
    5.013042, 5.019694, 5.029954, 5.044734, 5.064919, 5.091146, 5.123545, 
    5.161498, 5.203522, 5.247341, 5.290179, 5.329203, 5.361989, 5.386886, 
    5.403194, 5.411325, 5.413615, 5.407965, 5.397056, 5.382667, 5.366389, 
    5.350346, 5.335258, 5.322433, 5.312547, 5.306667, 5.305348, 5.308775, 
    5.316498, 5.328191, 5.342663, 5.358954, 5.37482, 5.38847, 5.398046, 
    5.401766, 5.398109, 5.386037, 5.365193, 5.336077, 5.300086, 5.259408, 
    5.216734, 5.174833, 5.136135, 5.102393, 5.074556, 5.052821, 5.03683, 
    5.025922,
  // momentumY(9,1, 0-49)
    5.018539, 5.027684, 5.041417, 5.060682, 5.086233, 5.118349, 5.15655, 
    5.19942, 5.244636, 5.289235, 5.330095, 5.364451, 5.390327, 5.406764, 
    5.413841, 5.412899, 5.408258, 5.395083, 5.37753, 5.357601, 5.33689, 
    5.31798, 5.300873, 5.28678, 5.275898, 5.269395, 5.267859, 5.271605, 
    5.28021, 5.293866, 5.31147, 5.332596, 5.354544, 5.375515, 5.393538, 
    5.406585, 5.412741, 5.410409, 5.398545, 5.376884, 5.346107, 5.307889, 
    5.264752, 5.219728, 5.175877, 5.135812, 5.10137, 5.073483, 5.052285, 
    5.037354,
  // momentumY(9,2, 0-49)
    5.026684, 5.039216, 5.057403, 5.082047, 5.113499, 5.151348, 5.194202, 
    5.239692, 5.284729, 5.326012, 5.360569, 5.386237, 5.401902, 5.407519, 
    5.403984, 5.393466, 5.38223, 5.362339, 5.339471, 5.315671, 5.292365, 
    5.272373, 5.254879, 5.240854, 5.229998, 5.223449, 5.221773, 5.225418, 
    5.234077, 5.248452, 5.26766, 5.291913, 5.318253, 5.345037, 5.370354, 
    5.392126, 5.40825, 5.416761, 5.416035, 5.405025, 5.383495, 5.35221, 
    5.312987, 5.268557, 5.222194, 5.177207, 5.136419, 5.101797, 5.074339, 
    5.054193,
  // momentumY(9,3, 0-49)
    5.037796, 5.054545, 5.077931, 5.108358, 5.145469, 5.18788, 5.233158, 
    5.278073, 5.319133, 5.353187, 5.377922, 5.392138, 5.395739, 5.389587, 
    5.375238, 5.355539, 5.338708, 5.313167, 5.286374, 5.260293, 5.236083, 
    5.216662, 5.200305, 5.187636, 5.177845, 5.171894, 5.170265, 5.173514, 
    5.181518, 5.195473, 5.21482, 5.240509, 5.269487, 5.300368, 5.331426, 
    5.360679, 5.385998, 5.405237, 5.416381, 5.417744, 5.408212, 5.3875, 
    5.356378, 5.316756, 5.271558, 5.224334, 5.17869, 5.137706, 5.103526, 
    5.07722,
  // momentumY(9,4, 0-49)
    5.052035, 5.073641, 5.102532, 5.138441, 5.180034, 5.224841, 5.269492, 
    5.310276, 5.3438, 5.367561, 5.380238, 5.381697, 5.372798, 5.355103, 
    5.330607, 5.30267, 5.281563, 5.251438, 5.221951, 5.194925, 5.171211, 
    5.153751, 5.139843, 5.129701, 5.121983, 5.117336, 5.116074, 5.11881, 
    5.125641, 5.138234, 5.156425, 5.182015, 5.211965, 5.245227, 5.280334, 
    5.31548, 5.34862, 5.37757, 5.400111, 5.414134, 5.417838, 5.409997, 
    5.390258, 5.359409, 5.319504, 5.273733, 5.225988, 5.18022, 5.139762, 
    5.106874,
  // momentumY(9,5, 0-49)
    5.06927, 5.096024, 5.130133, 5.170412, 5.21444, 5.258764, 5.299453, 
    5.332823, 5.356091, 5.367723, 5.367478, 5.356185, 5.335419, 5.307194, 
    5.273708, 5.238726, 5.214715, 5.180921, 5.149723, 5.122785, 5.100636, 
    5.086227, 5.075836, 5.069233, 5.064543, 5.061961, 5.061525, 5.063834, 
    5.069201, 5.079716, 5.095667, 5.119814, 5.149218, 5.18323, 5.220694, 
    5.260019, 5.299302, 5.336403, 5.369049, 5.394906, 5.411742, 5.417627, 
    5.411244, 5.392218, 5.361438, 5.321201, 5.275047, 5.227249, 5.182064, 
    5.142961,
  // momentumY(9,6, 0-49)
    5.088974, 5.120697, 5.159075, 5.201886, 5.245714, 5.28647, 5.320168, 
    5.343662, 5.355105, 5.354039, 5.341181, 5.318075, 5.28674, 5.249392, 
    5.208251, 5.167442, 5.141766, 5.105011, 5.072841, 5.046739, 5.026933, 
    5.016384, 5.01034, 5.008129, 5.007359, 5.007643, 5.008629, 5.010802, 
    5.014644, 5.022597, 5.035425, 5.056958, 5.084433, 5.117664, 5.155847, 
    5.197634, 5.241279, 5.284737, 5.325753, 5.361929, 5.390816, 5.410064, 
    5.417652, 5.412226, 5.393486, 5.362525, 5.321963, 5.275724, 5.22841, 
    5.184418,
  // momentumY(9,7, 0-49)
    5.110209, 5.146196, 5.187303, 5.230341, 5.2712, 5.305634, 5.330105, 
    5.342353, 5.341588, 5.328314, 5.30397, 5.270539, 5.230231, 5.185272, 
    5.137776, 5.092242, 5.065883, 5.026673, 4.994061, 4.969322, 4.952398, 
    4.94629, 4.94522, 4.948102, 4.952066, 4.956038, 4.959166, 4.961686, 
    4.96418, 4.969313, 4.978322, 4.996211, 5.020468, 5.051454, 5.088767, 
    5.131334, 5.177573, 5.225541, 5.273042, 5.317697, 5.356995, 5.388387, 
    5.409444, 5.418111, 5.413079, 5.394205, 5.362855, 5.321998, 5.275874, 
    5.22923,
  // momentumY(9,8, 0-49)
    5.131696, 5.170769, 5.212703, 5.253581, 5.289032, 5.315145, 5.329186, 
    5.329929, 5.317555, 5.293313, 5.25909, 5.217057, 5.16942, 5.118283, 
    5.06558, 5.016235, 4.989789, 4.94848, 4.915803, 4.892795, 4.879127, 
    4.877858, 4.882214, 4.890742, 4.900167, 4.908644, 4.914731, 4.918277, 
    4.919837, 4.922133, 4.926813, 4.940151, 4.959956, 4.987245, 5.022112, 
    5.063804, 5.110915, 5.161597, 5.213713, 5.264927, 5.312754, 5.354599, 
    5.387856, 5.410053, 5.419156, 5.413955, 5.394502, 5.362439, 5.321009, 
    5.274606,
  // momentumY(9,9, 0-49)
    5.152001, 5.192673, 5.233472, 5.270114, 5.29842, 5.315174, 5.318628, 
    5.308538, 5.285864, 5.252336, 5.21005, 5.161165, 5.107756, 5.051719, 
    4.994766, 4.942291, 4.915819, 4.872682, 4.84023, 4.81922, 4.809059, 
    4.812881, 4.822952, 4.837524, 4.85301, 4.866771, 4.876707, 4.882144, 
    4.883457, 4.883184, 4.883249, 4.891264, 4.905428, 4.927546, 4.95835, 
    4.997493, 5.043778, 5.095445, 5.150386, 5.2063, 5.260748, 5.311169, 
    5.354927, 5.389367, 5.412012, 5.420855, 5.414785, 5.39402, 5.360405, 
    5.317352,
  // momentumY(9,10, 0-49)
    5.169785, 5.210491, 5.248452, 5.279398, 5.299693, 5.307023, 5.300615, 
    5.281043, 5.249805, 5.208882, 5.160379, 5.106323, 5.048559, 4.988734, 
    4.928304, 4.873112, 4.845929, 4.801261, 4.769295, 4.750492, 4.743991, 
    4.753007, 4.768904, 4.789725, 4.811697, 4.831421, 4.846126, 4.854508, 
    4.856575, 4.854371, 4.849869, 4.852006, 4.859412, 4.874855, 4.899894, 
    4.934735, 4.978467, 5.029416, 5.085478, 5.144336, 5.203576, 5.260691, 
    5.313084, 5.358071, 5.392953, 5.41521, 5.422825, 5.414724, 5.391241, 
    5.354405,
  // momentumY(9,11, 0-49)
    5.184051, 5.223395, 5.257313, 5.281863, 5.294163, 5.292828, 5.27793, 
    5.25065, 5.212797, 5.166412, 5.113485, 5.055821, 4.994998, 4.932372, 
    4.869107, 4.811265, 4.781673, 4.735917, 4.704734, 4.688303, 4.685516, 
    4.699636, 4.72124, 4.748251, 4.776879, 4.803067, 4.823434, 4.835981, 
    4.840165, 4.837159, 4.828632, 4.824708, 4.824437, 4.831717, 4.849192, 
    4.877854, 4.917208, 4.965708, 5.021219, 5.081358, 5.143673, 5.205681, 
    5.264839, 5.318503, 5.363908, 5.398248, 5.41888, 5.423704, 5.411665, 
    5.383304,
  // momentumY(9,12, 0-49)
    5.194335, 5.231282, 5.260574, 5.278791, 5.28386, 5.275225, 5.253618, 
    5.220604, 5.178126, 5.128154, 5.072487, 5.012671, 4.949991, 4.885493, 
    4.82, 4.759103, 4.724104, 4.677974, 4.647959, 4.634027, 4.634865, 
    4.653734, 4.680614, 4.713413, 4.74852, 4.781399, 4.808202, 4.826231, 
    4.834251, 4.832163, 4.82086, 4.811296, 4.802845, 4.800652, 4.808741, 
    4.829211, 4.862217, 4.906439, 4.959705, 5.019504, 5.083271, 5.148478, 
    5.212607, 5.273064, 5.327098, 5.371778, 5.404087, 5.421196, 5.420952, 
    5.402519,
  // momentumY(9,13, 0-49)
    5.20077, 5.234771, 5.259482, 5.27208, 5.271227, 5.25703, 5.230669, 
    5.19392, 5.148717, 5.09689, 5.04002, 4.97939, 4.916002, 4.850582, 
    4.783556, 4.718486, 4.673654, 4.628222, 4.599886, 4.588519, 4.592689, 
    4.615596, 4.646937, 4.684716, 4.725712, 4.765153, 4.798926, 4.823727, 
    4.837541, 4.838665, 4.826695, 4.812769, 4.796377, 4.783873, 4.780921, 
    4.791139, 4.815689, 4.853671, 4.902922, 4.960753, 5.024401, 5.091208, 
    5.158616, 5.22405, 5.284799, 5.337901, 5.380161, 5.408309, 5.419418, 
    5.411558,
  // momentumY(9,14, 0-49)
    5.204044, 5.235059, 5.255784, 5.26395, 5.258807, 5.240928, 5.211757, 
    5.173126, 5.126891, 5.074712, 5.01796, 4.9577, 4.894693, 4.829371, 
    4.761736, 4.690343, 4.630024, 4.586733, 4.560706, 4.551862, 4.558817, 
    4.584635, 4.619225, 4.660789, 4.706684, 4.75217, 4.793106, 4.82573, 
    4.84728, 4.85427, 4.84457, 4.828547, 4.805531, 4.782758, 4.767636, 
    4.765727, 4.779678, 4.809348, 4.852722, 4.90692, 4.968901, 5.035783, 
    5.104878, 5.173582, 5.2392, 5.2988, 5.349137, 5.386735, 5.408215, 5.410872,
  // momentumY(9,15, 0-49)
    5.205245, 5.233704, 5.251448, 5.256646, 5.248955, 5.229216, 5.198977, 
    5.160035, 5.114126, 5.062756, 5.007135, 4.948183, 4.886503, 4.822322, 
    4.75529, 4.674098, 4.592133, 4.552732, 4.529696, 4.523179, 4.532108, 
    4.559325, 4.595654, 4.639558, 4.689092, 4.739789, 4.787691, 4.828758, 
    4.859601, 4.875039, 4.871017, 4.856003, 4.828897, 4.797172, 4.769747, 
    4.754407, 4.755836, 4.775146, 4.810735, 4.859603, 4.918382, 4.983872, 
    5.053164, 5.123552, 5.192328, 5.2566, 5.31316, 5.358506, 5.389058, 5.40165,
  // momentumY(9,16, 0-49)
    5.205641, 5.232349, 5.248367, 5.25215, 5.243571, 5.223566, 5.193663, 
    5.155571, 5.1109, 5.061044, 5.007129, 4.950017, 4.890282, 4.828084, 
    4.762897, 4.667199, 4.558082, 4.524595, 4.505179, 4.500589, 4.510473, 
    4.537367, 4.573853, 4.618652, 4.670533, 4.725457, 4.779788, 4.82938, 
    4.870381, 4.896234, 4.90115, 4.890569, 4.862889, 4.82492, 4.786451, 
    4.75743, 4.745025, 4.7522, 4.7782, 4.820086, 4.874176, 4.936878, 
    5.004986, 5.075613, 5.145999, 5.21328, 5.274343, 5.325768, 5.363969, 
    5.385563,
  // momentumY(9,17, 0-49)
    5.206429, 5.23244, 5.24809, 5.25195, 5.243927, 5.22491, 5.196322, 
    5.159752, 5.116711, 5.068528, 5.016322, 4.960996, 4.903182, 4.84309, 
    4.780164, 4.665139, 4.525096, 4.499957, 4.484663, 4.481379, 4.491128, 
    4.516054, 4.551351, 4.595904, 4.649085, 4.707342, 4.767391, 4.825082, 
    4.876275, 4.913509, 4.929801, 4.926649, 4.902213, 4.861757, 4.814963, 
    4.77341, 4.746902, 4.740796, 4.755741, 4.789182, 4.837222, 4.895868, 
    4.96155, 5.03114, 5.101774, 5.170614, 5.234653, 5.290627, 5.335063, 
    5.36453,
  // momentumY(9,18, 0-49)
    5.208497, 5.234978, 5.251599, 5.256881, 5.250602, 5.233477, 5.206757, 
    5.171896, 5.13033, 5.083377, 5.032204, 4.977786, 4.920807, 4.861402, 
    4.798707, 4.662005, 4.489505, 4.475817, 4.465091, 4.462282, 4.47091, 
    4.492671, 4.525987, 4.569733, 4.623669, 4.684685, 4.74978, 4.814837, 
    4.875535, 4.924022, 4.952873, 4.959058, 4.941103, 4.902152, 4.850769, 
    4.799243, 4.759669, 4.740109, 4.743153, 4.767068, 4.80796, 4.861491, 
    4.9237, 4.991181, 5.060933, 5.130117, 5.195842, 5.255026, 5.304377, 
    5.340523,
  // momentumY(9,19, 0-49)
    5.212205, 5.240322, 5.25919, 5.267125, 5.263608, 5.249043, 5.224416, 
    5.191014, 5.150217, 5.103388, 5.051769, 4.996344, 4.937584, 4.874966, 
    4.806328, 4.651233, 4.447761, 4.448816, 4.443101, 4.439723, 4.446472, 
    4.464695, 4.496089, 4.539269, 4.594101, 4.657805, 4.727543, 4.799196, 
    4.868299, 4.927033, 4.968306, 4.984324, 4.974784, 4.940611, 4.888542, 
    4.830527, 4.780185, 4.748146, 4.739299, 4.753189, 4.786242, 4.833904, 
    4.891861, 4.956418, 5.024415, 5.092998, 5.159379, 5.220663, 5.273758, 
    5.315415,
  // momentumY(9,20, 0-49)
    5.212728, 5.239095, 5.257136, 5.265122, 5.262591, 5.250175, 5.229265, 
    5.201706, 5.169541, 5.134852, 5.099675, 5.065902, 5.035129, 5.008301, 
    4.984965, 0, 4.281867, 4.296238, 4.319592, 4.349007, 4.384036, 4.42006, 
    4.463272, 4.513869, 4.573604, 4.641306, 4.715052, 4.791258, 4.865699, 
    4.931174, 4.981727, 5.005177, 5.003088, 4.974547, 4.924257, 4.862964, 
    4.804741, 4.762134, 4.742292, 4.746347, 4.771365, 4.812787, 4.866036, 
    4.927151, 4.99281, 5.06013, 5.12641, 5.188928, 5.244792, 5.290888,
  // momentumY(9,21, 0-49)
    5.21802, 5.246518, 5.267158, 5.277958, 5.278198, 5.26831, 5.249588, 
    5.223853, 5.193182, 5.159711, 5.125531, 5.092601, 5.062645, 5.036921, 
    5.015751, 0, 4.280171, 4.286097, 4.301404, 4.32449, 4.355588, 4.38597, 
    4.42638, 4.475754, 4.535542, 4.604822, 4.681754, 4.762756, 4.84341, 
    4.91684, 4.978211, 5.011083, 5.019394, 5.000573, 4.957034, 4.897546, 
    4.835649, 4.785192, 4.75563, 4.750137, 4.766894, 4.801638, 4.849658, 
    4.906757, 4.969437, 5.034751, 5.100053, 5.162745, 5.22009, 5.269087,
  // momentumY(9,22, 0-49)
    5.22302, 5.253256, 5.275841, 5.288589, 5.290601, 5.282212, 5.264708, 
    5.239964, 5.210128, 5.177406, 5.143931, 5.111705, 5.082527, 5.057864, 
    5.038573, 0, 4.278119, 4.278525, 4.288034, 4.306596, 4.335303, 4.361061, 
    4.399333, 4.447818, 4.507654, 4.578084, 4.657235, 4.741405, 4.825919, 
    4.904216, 4.972783, 5.011243, 5.026633, 5.015471, 4.978484, 4.922526, 
    4.859972, 4.804983, 4.768548, 4.755605, 4.765541, 4.794574, 4.838022, 
    4.891535, 4.95148, 5.014856, 5.079045, 5.141546, 5.199745, 5.250741,
  // momentumY(9,23, 0-49)
    5.226744, 5.258028, 5.281734, 5.295559, 5.298512, 5.290893, 5.27401, 
    5.249787, 5.220436, 5.188205, 5.155255, 5.1236, 5.095076, 5.07127, 
    5.053352, 0, 4.279414, 4.276551, 4.281965, 4.297147, 4.32407, 4.345681, 
    4.381749, 4.428933, 4.488155, 4.558842, 4.639098, 4.725091, 4.811872, 
    4.893102, 4.966422, 5.00808, 5.028121, 5.022609, 4.991148, 4.939076, 
    4.877542, 4.820482, 4.779746, 4.76159, 4.766459, 4.791107, 4.830965, 
    4.881619, 4.93934, 5.001071, 5.064211, 5.126318, 5.184858, 5.237008,
  // momentumY(9,24, 0-49)
    5.228496, 5.259939, 5.283836, 5.297881, 5.301076, 5.293717, 5.277114, 
    5.253204, 5.224204, 5.192366, 5.159845, 5.128648, 5.100616, 5.077384, 
    5.060251, 0, 4.283651, 4.279233, 4.282315, 4.295458, 4.321284, 4.339952, 
    4.374256, 4.42016, 4.47849, 4.548845, 4.629343, 4.716074, 4.803885, 
    4.886553, 4.962506, 5.005624, 5.028133, 5.025902, 4.997901, 4.948527, 
    4.888073, 4.830173, 4.787071, 4.765799, 4.767502, 4.789327, 4.826833, 
    4.875592, 4.931826, 4.992456, 5.054884, 5.116711, 5.175456, 5.228333,
  // momentumY(9,25, 0-49)
    5.22796, 5.258594, 5.281716, 5.295139, 5.297939, 5.290426, 5.27388, 
    5.250185, 5.221498, 5.190021, 5.157872, 5.127028, 5.099308, 5.07633, 
    5.059365, 0, 4.289196, 4.284725, 4.287505, 4.300285, 4.325872, 4.343461, 
    4.376945, 4.422066, 4.479642, 4.549365, 4.629392, 4.715792, 4.803343, 
    4.885863, 4.962089, 5.004999, 5.027723, 5.026116, 4.998996, 4.950472, 
    4.89053, 4.832613, 4.789001, 4.766916, 4.767715, 4.788686, 4.825451, 
    4.87359, 4.929327, 4.989579, 5.051758, 5.113479, 5.17228, 5.22539,
  // momentumY(9,26, 0-49)
    5.225247, 5.254143, 5.275551, 5.287515, 5.289261, 5.281141, 5.26438, 
    5.240758, 5.21231, 5.18114, 5.149289, 5.11869, 5.091106, 5.068068, 
    5.050664, 0, 4.295433, 4.292458, 4.29705, 4.311205, 4.33739, 4.355901, 
    4.389616, 4.434559, 4.491645, 4.560555, 4.639478, 4.724538, 4.810594, 
    4.891437, 4.965577, 5.006762, 5.027511, 5.023829, 4.99484, 4.945057, 
    4.88476, 4.827417, 4.78503, 4.764428, 4.766649, 4.788824, 4.826549, 
    4.875436, 4.931742, 4.99241, 5.054859, 5.116698, 5.175449, 5.22833,
  // momentumY(9,27, 0-49)
    5.220861, 5.247246, 5.266091, 5.275759, 5.275703, 5.266364, 5.248924, 
    5.225036, 5.196589, 5.16555, 5.133861, 5.103376, 5.075775, 5.052415, 
    5.034029, 0, 4.302463, 4.302832, 4.311277, 4.328385, 4.355904, 4.377017, 
    4.411754, 4.456905, 4.513578, 4.58136, 4.658477, 4.741166, 4.824496, 
    4.902151, 4.97192, 5.009845, 5.026492, 5.018219, 4.984942, 4.932204, 
    4.871093, 4.815196, 4.775881, 4.759018, 4.764867, 4.790172, 4.830435, 
    4.881328, 4.939181, 5.000987, 5.064165, 5.126294, 5.184847, 5.237001,
  // momentumY(9,28, 0-49)
    5.215629, 5.238973, 5.254549, 5.261092, 5.258357, 5.246945, 5.228058, 
    5.203263, 5.174317, 5.143045, 5.111273, 5.080747, 5.053013, 5.029168, 
    5.009374, 0, 4.311146, 4.317119, 4.331298, 4.35264, 4.382026, 4.406691, 
    4.442622, 4.4878, 4.543655, 4.609676, 4.684156, 4.763472, 4.842965, 
    4.916097, 4.979532, 5.0127, 5.023324, 5.008373, 4.969041, 4.912435, 
    4.850762, 4.797608, 4.763256, 4.75213, 4.763408, 4.793327, 4.837316, 
    4.891145, 4.951268, 5.014741, 5.078983, 5.141513, 5.199726, 5.250731,
  // momentumY(9,29, 0-49)
    5.210575, 5.230656, 5.242446, 5.245065, 5.238635, 5.224026, 5.202578, 
    5.175876, 5.145615, 5.11352, 5.081297, 5.050559, 5.022669, 4.99836, 
    4.977002, 0, 4.32097, 4.335202, 4.357126, 4.384002, 4.415863, 4.444396, 
    4.481161, 4.525657, 4.579839, 4.643129, 4.713893, 4.78861, 4.862862, 
    4.929764, 4.984661, 5.011045, 5.013606, 4.990396, 4.944409, 4.88464, 
    4.824273, 4.776336, 4.749413, 4.746114, 4.764445, 4.80021, 4.84885, 
    4.906308, 4.96919, 5.034617, 5.099981, 5.162707, 5.22007, 5.269075,
  // momentumY(9,30, 0-49)
    5.211185, 5.232265, 5.243868, 5.245254, 5.236584, 5.218601, 5.192334, 
    5.158899, 5.119413, 5.074954, 5.0265, 4.974833, 4.92029, 4.862335, 
    4.799018, 4.650102, 4.46623, 4.474145, 4.474097, 4.474111, 4.482029, 
    4.496277, 4.523712, 4.562758, 4.613616, 4.67399, 4.741224, 4.811243, 
    4.879523, 4.938704, 4.982891, 5.000132, 4.992626, 4.960247, 4.908324, 
    4.847715, 4.791922, 4.752495, 4.735684, 4.742134, 4.768816, 4.811302, 
    4.865192, 4.926679, 4.992549, 5.059987, 5.126332, 5.188886, 5.244769, 
    5.290876,
  // momentumY(9,31, 0-49)
    5.20908, 5.227884, 5.236427, 5.234247, 5.221874, 5.200438, 5.171289, 
    5.135762, 5.095062, 5.050255, 5.002267, 4.951888, 4.899677, 4.845722, 
    4.789222, 4.658228, 4.501397, 4.496706, 4.493328, 4.495354, 4.506206, 
    4.525119, 4.554814, 4.594297, 4.643971, 4.701432, 4.764091, 4.828028, 
    4.888942, 4.939219, 4.972041, 4.980291, 4.964257, 4.925714, 4.87197, 
    4.814879, 4.767239, 4.738547, 4.732779, 4.749048, 4.783735, 4.832435, 
    4.89102, 4.955945, 5.024151, 5.092851, 5.159298, 5.220619, 5.273735, 
    5.315403,
  // momentumY(9,32, 0-49)
    5.209422, 5.227388, 5.234317, 5.229859, 5.214752, 5.190379, 5.15834, 
    5.120173, 5.077215, 5.030576, 4.981167, 4.929723, 4.876769, 4.822464, 
    4.766259, 4.657221, 4.530038, 4.515179, 4.508562, 4.511379, 4.524328, 
    4.547682, 4.579953, 4.620469, 4.669526, 4.724418, 4.782448, 4.839732, 
    4.892161, 4.932154, 4.95264, 4.951416, 4.927637, 4.885253, 4.833202, 
    4.783412, 4.747004, 4.730926, 4.736993, 4.76317, 4.805598, 4.860101, 
    4.922898, 4.990724, 5.060675, 5.129973, 5.195764, 5.254982, 5.304353, 
    5.340511,
  // momentumY(9,33, 0-49)
    5.211784, 5.230331, 5.23714, 5.231805, 5.215128, 5.188638, 5.154125, 
    5.113319, 5.067709, 5.018507, 4.966658, 4.912882, 4.857656, 4.801088, 
    4.742635, 4.653386, 4.555256, 4.532505, 4.522496, 4.524918, 4.538918, 
    4.565711, 4.600144, 4.641606, 4.68998, 4.742125, 4.795075, 4.84495, 
    4.887879, 4.916761, 4.925084, 4.915268, 4.8861, 4.843475, 4.797151, 
    4.758084, 4.735029, 4.73236, 4.75014, 4.785647, 4.835072, 4.894595, 
    4.960809, 5.030715, 5.101532, 5.170478, 5.234578, 5.290584, 5.33504, 
    5.364517,
  // momentumY(9,34, 0-49)
    5.215219, 5.235668, 5.243885, 5.23924, 5.222435, 5.195026, 5.158927, 
    5.11603, 5.067999, 5.016191, 4.961662, 4.905194, 4.847309, 4.788183, 
    4.727444, 4.6529, 4.580625, 4.55162, 4.538008, 4.538926, 4.552721, 
    4.581357, 4.616908, 4.658594, 4.70565, 4.754443, 4.80167, 4.843497, 
    4.87642, 4.894343, 4.89206, 4.875939, 4.844918, 4.806159, 4.769204, 
    4.743195, 4.734305, 4.744707, 4.773262, 4.816971, 4.872271, 4.935742, 
    5.004318, 5.075227, 5.145776, 5.213154, 5.274272, 5.325727, 5.363947, 
    5.38555,
  // momentumY(9,35, 0-49)
    5.218414, 5.241881, 5.252987, 5.250708, 5.235466, 5.208694, 5.172336, 
    5.12841, 5.078754, 5.02491, 4.968103, 4.90927, 4.849085, 4.787934, 
    4.725807, 4.660797, 4.609091, 4.575197, 4.557967, 4.556472, 4.56875, 
    4.597325, 4.632507, 4.673204, 4.717884, 4.762468, 4.803359, 4.83689, 
    4.860095, 4.868361, 4.85827, 4.839107, 4.810142, 4.778883, 4.753745, 
    4.741656, 4.746446, 4.768659, 4.806472, 4.856906, 4.916722, 4.98287, 
    5.052571, 5.123204, 5.192127, 5.256485, 5.313095, 5.358469, 5.389037, 
    5.401639,
  // momentumY(9,36, 0-49)
    5.219895, 5.247176, 5.262488, 5.264244, 5.252396, 5.228087, 5.193159, 
    5.149686, 5.099665, 5.044836, 4.98664, 4.926233, 4.864524, 4.80219, 
    4.739642, 4.680242, 4.642906, 4.605454, 4.584847, 4.580313, 4.589905, 
    4.616549, 4.649711, 4.687962, 4.729007, 4.768494, 4.802673, 4.828212, 
    4.842849, 4.843726, 4.829322, 4.810611, 4.787079, 4.765726, 4.753314, 
    4.754615, 4.771617, 4.803811, 4.849074, 4.904593, 4.967452, 5.034897, 
    5.104344, 5.173264, 5.239013, 5.29869, 5.349073, 5.3867, 5.408195, 
    5.410862,
  // momentumY(9,37, 0-49)
    5.218255, 5.249717, 5.27024, 5.277552, 5.270936, 5.25105, 5.219474, 
    5.178236, 5.129437, 5.075015, 5.016646, 4.955743, 4.893483, 4.830852, 
    4.76865, 4.712382, 4.683611, 4.643882, 4.620321, 4.612436, 4.618487, 
    4.641649, 4.671282, 4.705679, 4.741915, 4.775605, 4.803057, 4.82145, 
    4.829312, 4.825551, 4.810279, 4.794975, 4.779095, 4.768571, 4.768416, 
    4.7816, 4.808813, 4.848932, 4.899767, 4.958707, 5.023099, 5.090394, 
    5.158112, 5.223743, 5.284613, 5.33779, 5.380095, 5.408271, 5.419396, 
    5.411546,
  // momentumY(9,38, 0-49)
    5.212383, 5.247881, 5.274166, 5.288225, 5.288517, 5.274992, 5.248788, 
    5.21174, 5.165967, 5.113562, 5.056436, 4.996264, 4.934503, 4.87243, 
    4.811168, 4.756728, 4.73197, 4.691082, 4.665075, 4.653807, 4.65584, 
    4.674464, 4.699435, 4.72888, 4.759443, 4.786973, 4.808064, 4.820529, 
    4.823663, 4.81791, 4.804527, 4.794577, 4.787253, 4.787226, 4.797941, 
    4.821002, 4.856258, 4.902263, 4.956853, 5.017594, 5.082009, 5.147655, 
    5.212077, 5.272727, 5.326886, 5.371646, 5.404006, 5.421148, 5.420925, 
    5.402503,
  // momentumY(9,39, 0-49)
    5.20167, 5.240501, 5.272511, 5.294001, 5.302503, 5.297089, 5.278226, 
    5.247378, 5.20655, 5.157911, 5.103568, 5.045445, 4.985273, 4.924599, 
    4.864816, 4.811718, 4.787943, 4.746778, 4.718848, 4.70439, 4.702281, 
    4.715828, 4.73548, 4.759322, 4.783782, 4.805178, 4.82057, 4.828451, 
    4.828772, 4.823126, 4.813404, 4.809672, 4.810735, 4.820044, 4.839785, 
    4.870599, 4.911798, 4.96177, 5.018401, 5.079369, 5.142285, 5.204723, 
    5.264188, 5.318067, 5.363621, 5.398062, 5.418763, 5.423631, 5.411623, 
    5.383276,
  // momentumY(9,40, 0-49)
    5.186132, 5.22708, 5.264103, 5.293013, 5.310456, 5.314495, 5.304725, 
    5.282016, 5.248078, 5.205032, 5.155106, 5.100437, 5.043005, 4.984615, 
    4.926899, 4.87519, 4.850765, 4.809989, 4.780656, 4.763356, 4.757268, 
    4.765635, 4.779768, 4.797813, 4.816178, 4.8318, 4.84232, 4.846885, 
    4.845916, 4.841768, 4.836526, 4.838995, 4.847562, 4.864634, 4.891436, 
    4.927948, 4.973135, 5.025293, 5.082327, 5.141959, 5.201804, 5.259393, 
    5.312152, 5.357416, 5.392503, 5.414909, 5.422629, 5.414599, 5.391162, 
    5.354355,
  // momentumY(9,41, 0-49)
    5.166451, 5.207902, 5.248558, 5.28407, 5.310394, 5.324593, 5.325236, 
    5.312375, 5.287194, 5.251593, 5.207793, 5.158082, 5.10465, 5.049539, 
    4.994611, 4.944724, 4.91911, 4.879265, 4.849064, 4.829385, 4.819679, 
    4.823095, 4.831874, 4.844314, 4.856938, 4.867391, 4.873917, 4.876226, 
    4.875024, 4.873092, 4.872416, 4.880478, 4.895287, 4.918398, 4.950332, 
    4.990605, 5.037953, 5.090587, 5.146398, 5.203084, 5.258206, 5.309211, 
    5.353455, 5.388292, 5.41125, 5.42033, 5.414435, 5.393792, 5.360259, 
    5.317256,
  // momentumY(9,42, 0-49)
    5.143857, 5.184021, 5.226386, 5.266863, 5.301079, 5.325276, 5.336976, 
    5.335222, 5.320437, 5.294066, 5.258155, 5.215016, 5.166993, 5.116336, 
    5.06512, 5.017797, 4.99126, 4.952888, 4.922406, 4.90091, 4.888094, 
    4.887012, 4.890862, 4.898168, 4.905657, 4.911681, 4.915056, 4.915931, 
    4.915131, 4.915613, 4.919096, 4.931798, 4.951411, 4.978819, 5.014019, 
    5.056201, 5.103926, 5.155319, 5.208214, 5.260242, 5.308877, 5.35149, 
    5.38544, 5.408236, 5.417833, 5.413025, 5.393868, 5.362019, 5.320735, 
    5.274421,
  // momentumY(9,43, 0-49)
    5.119925, 5.157089, 5.198948, 5.24208, 5.282256, 5.315266, 5.337736, 
    5.347641, 5.344442, 5.32887, 5.302574, 5.267717, 5.226689, 5.18188, 
    5.135561, 5.09184, 5.065246, 5.028996, 4.998917, 4.976262, 4.960958, 
    4.95599, 4.955519, 4.958347, 4.961455, 4.963848, 4.964833, 4.96487, 
    4.964771, 4.967505, 4.974444, 4.990649, 5.013561, 5.043531, 5.080167, 
    5.122412, 5.168684, 5.217022, 5.265179, 5.3107, 5.350989, 5.383418, 
    5.405475, 5.415052, 5.410805, 5.392574, 5.361722, 5.321233, 5.275365, 
    5.228883,
  // momentumY(9,44, 0-49)
    5.096272, 5.129057, 5.168241, 5.211352, 5.254784, 5.29438, 5.326228, 
    5.34737, 5.35621, 5.352563, 5.337418, 5.312571, 5.280278, 5.24296, 
    5.203005, 5.164229, 5.138921, 5.105624, 5.076772, 5.053725, 5.036647, 
    5.028522, 5.024458, 5.023581, 5.023133, 5.022689, 5.021945, 5.021548, 
    5.022201, 5.026792, 5.036315, 5.054803, 5.079486, 5.110286, 5.146511, 
    5.186906, 5.22978, 5.273088, 5.314514, 5.351556, 5.381634, 5.402251, 
    5.411257, 5.407187, 5.389662, 5.359727, 5.319985, 5.274365, 5.22749, 
    5.183779,
  // momentumY(9,45, 0-49)
    5.074281, 5.101814, 5.136524, 5.17699, 5.220571, 5.263685, 5.302406, 
    5.333194, 5.353523, 5.36219, 5.359307, 5.346044, 5.324288, 5.296298, 
    5.264447, 5.232249, 5.209951, 5.180675, 5.154027, 5.131465, 5.113417, 
    5.102954, 5.096113, 5.092372, 5.089212, 5.08668, 5.084756, 5.084169, 
    5.085434, 5.091334, 5.102482, 5.122004, 5.14693, 5.17682, 5.210737, 
    5.247275, 5.284656, 5.320791, 5.353364, 5.379928, 5.39808, 5.405691, 
    5.401236, 5.384155, 5.355194, 5.316544, 5.271692, 5.224903, 5.180446, 
    5.141823,
  // momentumY(9,46, 0-49)
    5.0549, 5.07686, 5.105901, 5.141548, 5.18226, 5.22542, 5.26764, 5.305339, 
    5.335418, 5.355771, 5.36553, 5.365007, 5.355437, 5.338662, 5.316822, 
    5.293051, 5.275785, 5.251806, 5.228491, 5.207395, 5.189259, 5.177374, 
    5.168643, 5.162926, 5.157879, 5.153938, 5.151259, 5.150574, 5.152169, 
    5.158724, 5.17048, 5.189789, 5.213448, 5.240694, 5.270373, 5.30097, 
    5.330666, 5.357411, 5.379015, 5.393284, 5.398237, 5.392398, 5.375129, 
    5.346938, 5.309633, 5.26622, 5.22047, 5.176284, 5.136996, 5.104896,
  // momentumY(9,47, 0-49)
    5.038558, 5.055104, 5.07795, 5.107332, 5.142719, 5.182619, 5.224613, 
    5.265657, 5.302625, 5.332863, 5.354623, 5.367231, 5.371015, 5.367095, 
    5.3571, 5.343633, 5.333583, 5.316318, 5.297566, 5.279008, 5.261748, 
    5.249465, 5.23981, 5.233042, 5.226902, 5.222136, 5.219, 5.218166, 
    5.219665, 5.226124, 5.237422, 5.255292, 5.276211, 5.299119, 5.322676, 
    5.345291, 5.365184, 5.380476, 5.389296, 5.389965, 5.381234, 5.362558, 
    5.334355, 5.298147, 5.256485, 5.212605, 5.169889, 5.131297, 5.098928, 
    5.073874,
  // momentumY(9,48, 0-49)
    5.025191, 5.036808, 5.053524, 5.076003, 5.104483, 5.138533, 5.17689, 
    5.217495, 5.257764, 5.295023, 5.326963, 5.351994, 5.369394, 5.379289, 
    5.382505, 5.380936, 5.380241, 5.371087, 5.358146, 5.343263, 5.327931, 
    5.316406, 5.306894, 5.300048, 5.293569, 5.288468, 5.285032, 5.28385, 
    5.284679, 5.29018, 5.29989, 5.31511, 5.331882, 5.348882, 5.364614, 
    5.377472, 5.385822, 5.388123, 5.38307, 5.369785, 5.348024, 5.318344, 
    5.282197, 5.241826, 5.199984, 5.1595, 5.122818, 5.091662, 5.06691, 
    5.048687,
  // momentumY(9,49, 0-49)
    5.012385, 5.018913, 5.028864, 5.043107, 5.062448, 5.087427, 5.118075, 
    5.153737, 5.193004, 5.233839, 5.273879, 5.31083, 5.342823, 5.368688, 
    5.388059, 5.402215, 5.418763, 5.421006, 5.415788, 5.405649, 5.392869, 
    5.385442, 5.379874, 5.377387, 5.372908, 5.368307, 5.363704, 5.359727, 
    5.355256, 5.355647, 5.359989, 5.371101, 5.38187, 5.390671, 5.395897, 
    5.396035, 5.389802, 5.3763, 5.355184, 5.326793, 5.292233, 5.253324, 
    5.212403, 5.171985, 5.134371, 5.101318, 5.073847, 5.052252, 5.036246, 
    5.025198,
  // momentumY(10,0, 0-49)
    5.063582, 5.085031, 5.112928, 5.146696, 5.184947, 5.225497, 5.265574, 
    5.302221, 5.332746, 5.355133, 5.368267, 5.371976, 5.366912, 5.354355, 
    5.335983, 5.3139, 5.291661, 5.267425, 5.244224, 5.223267, 5.205225, 
    5.190944, 5.179907, 5.172104, 5.167113, 5.164995, 5.165788, 5.169702, 
    5.176876, 5.187829, 5.202584, 5.221438, 5.243492, 5.268015, 5.293913, 
    5.31977, 5.34392, 5.364543, 5.379786, 5.387915, 5.38752, 5.377726, 
    5.358419, 5.3304, 5.295416, 5.256012, 5.215207, 5.176044, 5.141145, 
    5.112394,
  // momentumY(10,1, 0-49)
    5.079928, 5.105417, 5.137311, 5.174423, 5.214681, 5.255301, 5.293159, 
    5.325284, 5.349298, 5.363727, 5.368092, 5.362825, 5.349079, 5.32849, 
    5.302971, 5.274961, 5.249591, 5.22163, 5.19565, 5.1729, 5.153946, 
    5.139993, 5.129792, 5.123188, 5.119247, 5.117973, 5.119292, 5.123413, 
    5.130458, 5.141384, 5.156361, 5.176321, 5.200119, 5.227235, 5.256737, 
    5.287312, 5.31734, 5.344975, 5.368256, 5.385231, 5.394138, 5.393606, 
    5.382902, 5.362143, 5.332445, 5.295923, 5.255486, 5.214435, 5.175961, 
    5.142664,
  // momentumY(10,2, 0-49)
    5.100276, 5.12977, 5.1649, 5.203756, 5.243615, 5.281312, 5.313743, 
    5.338332, 5.35337, 5.358143, 5.352868, 5.338513, 5.316582, 5.288897, 
    5.257421, 5.224789, 5.197577, 5.167107, 5.139554, 5.116156, 5.097363, 
    5.084681, 5.076171, 5.071518, 5.069331, 5.069472, 5.071693, 5.076145, 
    5.082903, 5.093283, 5.107612, 5.127469, 5.151559, 5.179631, 5.210985, 
    5.244498, 5.27869, 5.311812, 5.34193, 5.367047, 5.385226, 5.394764, 
    5.394402, 5.383549, 5.362504, 5.332596, 5.296147, 5.256245, 5.216292, 
    5.179459,
  // momentumY(10,3, 0-49)
    5.123564, 5.156494, 5.193518, 5.232036, 5.268888, 5.30088, 5.325299, 
    5.340286, 5.344973, 5.33944, 5.324524, 5.3016, 5.27236, 5.238668, 
    5.202416, 5.166353, 5.138496, 5.1065, 5.078358, 5.055256, 5.03751, 
    5.026891, 5.020802, 5.018765, 5.018983, 5.021102, 5.024645, 5.029631, 
    5.036055, 5.045497, 5.058444, 5.077137, 5.100204, 5.127726, 5.159303, 
    5.194069, 5.230758, 5.267785, 5.303344, 5.335496, 5.362273, 5.381793, 
    5.39242, 5.392964, 5.382909, 5.362636, 5.33356, 5.298093, 5.259374, 
    5.220767,
  // momentumY(10,4, 0-49)
    5.148277, 5.183551, 5.220681, 5.256588, 5.288019, 5.312116, 5.326862, 
    5.331258, 5.325281, 5.309696, 5.285806, 5.25523, 5.219736, 5.181118, 
    5.141133, 5.102629, 5.075132, 5.042326, 5.01433, 4.99224, 4.976225, 
    4.968293, 4.965206, 4.966337, 4.969534, 4.974173, 4.979482, 4.985287, 
    4.991461, 4.999736, 5.010735, 5.027388, 5.048301, 5.073945, 5.104287, 
    5.138782, 5.176426, 5.215847, 5.255407, 5.293285, 5.327562, 5.356293, 
    5.377622, 5.389924, 5.392003, 5.383332, 5.364291, 5.336296, 5.301751, 
    5.263733,
  // momentumY(10,5, 0-49)
    5.17261, 5.208737, 5.244016, 5.275208, 5.299335, 5.314187, 5.318586, 
    5.31239, 5.29629, 5.271561, 5.239791, 5.202709, 5.162052, 5.119503, 
    5.076645, 5.036462, 5.010109, 4.97695, 4.949606, 4.929027, 4.91522, 
    4.910427, 4.91076, 4.915475, 4.92213, 4.929779, 4.937321, 4.944317, 
    4.950469, 4.957533, 4.96622, 4.980175, 4.998003, 5.020619, 5.048433, 
    5.081285, 5.118479, 5.158883, 5.201038, 5.243255, 5.283694, 5.320426, 
    5.351492, 5.375001, 5.389269, 5.393025, 5.385661, 5.367476, 5.339813, 
    5.305001,
  // momentumY(10,6, 0-49)
    5.194726, 5.230039, 5.261647, 5.286497, 5.302191, 5.307335, 5.301603, 
    5.285583, 5.260492, 5.227921, 5.189589, 5.147222, 5.102467, 5.056863, 
    5.011828, 4.97053, 4.945855, 4.912601, 4.886216, 4.867458, 4.85615, 
    4.854763, 4.858765, 4.867326, 4.877797, 4.888885, 4.899129, 4.907778, 
    4.914294, 4.920318, 4.926564, 4.9374, 4.951415, 4.97002, 4.994144, 
    5.024087, 5.059518, 5.099563, 5.142944, 5.188095, 5.233257, 5.276544, 
    5.315973, 5.349518, 5.375189, 5.391176, 5.396054, 5.389062, 5.370367, 
    5.341236,
  // momentumY(10,7, 0-49)
    5.213053, 5.245964, 5.27248, 5.290026, 5.296961, 5.292734, 5.27777, 
    5.253204, 5.220595, 5.181672, 5.138168, 5.091727, 5.04387, 4.995987, 
    4.949328, 4.907313, 4.88458, 4.851351, 4.826089, 4.809305, 4.800615, 
    4.802724, 4.810457, 4.822952, 4.837451, 4.852314, 4.865723, 4.876563, 
    4.88401, 4.889411, 4.893355, 4.900923, 4.910622, 4.924387, 4.94375, 
    4.969565, 5.001939, 5.040301, 5.083554, 5.130239, 5.178657, 5.226962, 
    5.27318, 5.315236, 5.350972, 5.378225, 5.394969, 5.399563, 5.391072, 
    5.369621,
  // momentumY(10,8, 0-49)
    5.226548, 5.255755, 5.276319, 5.286304, 5.284873, 5.272231, 5.249386, 
    5.217844, 5.179329, 5.135591, 5.088283, 5.038926, 4.98889, 4.939411, 
    4.891582, 4.849094, 4.828224, 4.795094, 4.771032, 4.756248, 4.750131, 
    4.755633, 4.766952, 4.783258, 4.801815, 4.820665, 4.837659, 4.851306, 
    4.860435, 4.865911, 4.868018, 4.872491, 4.877636, 4.885912, 4.899523, 
    4.919997, 4.947987, 4.983297, 5.02504, 5.071846, 5.122056, 5.173835, 
    5.225216, 5.274106, 5.318265, 5.355324, 5.38286, 5.39859, 5.40069, 
    5.388237,
  // momentumY(10,9, 0-49)
    5.234836, 5.259479, 5.273821, 5.276622, 5.26777, 5.248077, 5.218955, 
    5.182111, 5.139313, 5.09224, 5.042422, 4.991228, 4.93987, 4.889423, 
    4.840813, 4.797938, 4.778379, 4.745469, 4.722646, 4.709779, 4.706027, 
    4.714598, 4.729111, 4.748862, 4.77128, 4.794157, 4.815078, 4.832183, 
    4.843925, 4.850475, 4.851599, 4.853556, 4.854271, 4.856665, 4.863659, 
    4.877585, 4.899804, 4.930608, 4.969382, 5.014863, 5.0654, 5.119133, 
    5.17407, 5.228092, 5.27892, 5.324071, 5.360898, 5.386709, 5.399065, 
    5.396215,
  // momentumY(10,10, 0-49)
    5.238247, 5.257951, 5.266341, 5.262815, 5.247848, 5.222678, 5.188955, 
    5.148462, 5.102916, 5.053882, 5.002743, 4.950707, 4.898828, 4.848012, 
    4.798991, 4.755602, 4.736162, 4.703743, 4.682203, 4.671069, 4.66929, 
    4.68035, 4.697388, 4.71993, 4.745744, 4.772466, 4.797513, 4.818703, 
    4.834116, 4.843032, 4.844454, 4.844961, 4.841871, 4.838394, 4.838163, 
    4.844429, 4.859446, 4.88419, 4.918439, 4.961081, 5.01046, 5.064648, 
    5.121579, 5.17908, 5.234825, 5.286284, 5.330706, 5.365195, 5.38696, 
    5.393692,
  // momentumY(10,11, 0-49)
    5.237722, 5.252574, 5.255694, 5.247005, 5.227397, 5.198365, 5.161659, 
    5.119038, 5.072123, 5.022343, 4.970935, 4.918961, 4.86732, 4.81674, 
    4.767717, 4.723385, 4.702055, 4.670654, 4.650481, 4.64079, 4.640394, 
    4.653071, 4.671667, 4.696053, 4.724506, 4.754633, 4.783804, 4.809594, 
    4.829752, 4.842523, 4.845928, 4.846569, 4.840914, 4.832191, 4.824595, 
    4.822354, 4.828823, 4.845907, 4.873978, 4.912177, 4.958867, 5.012014, 
    5.069425, 5.128822, 5.187816, 5.243847, 5.294146, 5.335773, 5.365799, 
    5.381611,
  // momentumY(10,12, 0-49)
    5.234626, 5.245103, 5.243909, 5.231354, 5.20858, 5.177192, 5.138937, 
    5.095491, 5.048359, 4.998839, 4.948044, 4.896914, 4.84622, 4.796515, 
    4.748018, 4.701878, 4.675796, 4.646248, 4.627597, 4.618956, 4.619151, 
    4.632289, 4.651206, 4.676237, 4.706321, 4.739155, 4.772195, 4.802876, 
    4.828703, 4.846828, 4.854155, 4.856939, 4.85062, 4.838054, 4.82369, 
    4.812641, 4.809513, 4.817426, 4.837632, 4.869717, 4.912129, 4.962729, 
    5.019142, 5.078934, 5.139617, 5.198605, 5.253157, 5.300396, 5.33741, 
    5.361478,
  // momentumY(10,13, 0-49)
    5.230535, 5.237388, 5.232965, 5.21782, 5.193212, 5.160748, 5.122097, 
    5.078829, 5.032333, 4.983805, 4.934273, 4.884608, 4.835494, 4.787343, 
    4.740097, 4.690714, 4.656355, 4.629813, 4.612917, 4.604844, 4.60468, 
    4.616896, 4.634736, 4.65907, 4.689609, 4.724247, 4.760649, 4.796208, 
    4.828288, 4.853024, 4.866192, 4.873289, 4.868722, 4.854521, 4.834921, 
    4.81561, 4.802438, 4.8, 4.810771, 4.835072, 4.871596, 4.918133, 4.972108, 
    5.030878, 5.091822, 5.152305, 5.209641, 5.261067, 5.303789, 5.335109,
  // momentumY(10,14, 0-49)
    5.22699, 5.231134, 5.224566, 5.207964, 5.182598, 5.150006, 5.111754, 
    5.069297, 5.023933, 4.976803, 4.928903, 4.881094, 4.834053, 4.788131, 
    4.743088, 4.688396, 4.642111, 4.619964, 4.605116, 4.597078, 4.595531, 
    4.605345, 4.620689, 4.643006, 4.672795, 4.708239, 4.747289, 4.787376, 
    4.82584, 4.857959, 4.878545, 4.891905, 4.89165, 4.878604, 4.856218, 
    4.830238, 4.807499, 4.794166, 4.79429, 4.80929, 4.838372, 4.879369, 
    4.929523, 4.985952, 5.04586, 5.106551, 5.16538, 5.219721, 5.266939, 
    5.304432,
  // momentumY(10,15, 0-49)
    5.225293, 5.227697, 5.219958, 5.202792, 5.177416, 5.145269, 5.107808, 
    5.066401, 5.02229, 4.976607, 4.930377, 4.88452, 4.839792, 4.79663, 
    4.75483, 4.69235, 4.631154, 4.614925, 4.602443, 4.593904, 4.58998, 
    4.595966, 4.607544, 4.62669, 4.65465, 4.689934, 4.730808, 4.7748, 
    4.819294, 4.85896, 4.887938, 4.908922, 4.915213, 4.906217, 4.884106, 
    4.854033, 4.823288, 4.799448, 4.788349, 4.792909, 4.813193, 4.847295, 
    4.892347, 4.94524, 5.002972, 5.062758, 5.12198, 5.17813, 5.228736, 
    5.271329,
  // momentumY(10,16, 0-49)
    5.226336, 5.227925, 5.219817, 5.202703, 5.177724, 5.146221, 5.109568, 
    5.06908, 5.025991, 4.981462, 4.936589, 4.892404, 4.84983, 4.809532, 
    4.771629, 4.699264, 4.621652, 4.61295, 4.603134, 4.593575, 4.586397, 
    4.587306, 4.594104, 4.609207, 4.634496, 4.668808, 4.710706, 4.757823, 
    4.807619, 4.854417, 4.892068, 4.921228, 4.935552, 4.933044, 4.914313, 
    4.883314, 4.847099, 4.81419, 4.792173, 4.785765, 4.796284, 4.822381, 
    4.861237, 4.909564, 4.964163, 5.022121, 5.08082, 5.137845, 5.190862, 
    5.237532,
  // momentumY(10,17, 0-49)
    5.230514, 5.23212, 5.224253, 5.207549, 5.183083, 5.152126, 5.116007, 
    5.076031, 5.033445, 4.989463, 4.945265, 4.902009, 4.860803, 4.822589, 
    4.787977, 4.705591, 4.612271, 4.612747, 4.605839, 4.594719, 4.583512, 
    4.578328, 4.579618, 4.590136, 4.612224, 4.645008, 4.687278, 4.736743, 
    4.790919, 4.844021, 4.890014, 4.927098, 4.949994, 4.955523, 4.94271, 
    4.913936, 4.875333, 4.835699, 4.804019, 4.7869, 4.787251, 4.804621, 
    4.836472, 4.879438, 4.930146, 4.985555, 5.04301, 5.100143, 5.154733, 
    5.204546,
  // momentumY(10,18, 0-49)
    5.237718, 5.240082, 5.232924, 5.216834, 5.19283, 5.162156, 5.126127, 
    5.086053, 5.043212, 4.998859, 4.954231, 4.910549, 4.86899, 4.830619, 
    4.796376, 4.707914, 4.602833, 4.613844, 4.60993, 4.59652, 4.580455, 
    4.568354, 4.563672, 4.569397, 4.588124, 4.619167, 4.66143, 4.712628, 
    4.770273, 4.82866, 4.882247, 4.92637, 4.957467, 4.971514, 4.966166, 
    4.942143, 4.904187, 4.860658, 4.821369, 4.794617, 4.785073, 4.793501, 
    4.817908, 4.85501, 4.901318, 4.953671, 5.009349, 5.066003, 5.121474, 
    5.173612,
  // momentumY(10,19, 0-49)
    5.247415, 5.251267, 5.245289, 5.230013, 5.20642, 5.175728, 5.139245, 
    5.098292, 5.054173, 5.008155, 4.961453, 4.915181, 4.870294, 4.827582, 
    4.788054, 4.702839, 4.595904, 4.617163, 4.615731, 4.598713, 4.576507, 
    4.556717, 4.545831, 4.546948, 4.562612, 4.592149, 4.634409, 4.687026, 
    4.747424, 4.810097, 4.870316, 4.920206, 4.958426, 4.980475, 4.982996, 
    4.965231, 4.930353, 4.885727, 4.841322, 4.806689, 4.788195, 4.788025, 
    4.80498, 4.836047, 4.87772, 4.926739, 4.980312, 5.036072, 5.091892, 
    5.14567,
  // momentumY(10,20, 0-49)
    5.253863, 5.255918, 5.248505, 5.232355, 5.208736, 5.179231, 5.145556, 
    5.109469, 5.072702, 5.036943, 5.003791, 4.974656, 4.950539, 4.931577, 
    4.916345, 0, 4.529047, 4.533604, 4.533447, 4.529254, 4.524078, 4.517531, 
    4.516744, 4.524277, 4.543463, 4.574782, 4.617994, 4.671397, 4.732827, 
    4.797443, 4.86176, 4.91475, 4.957507, 4.985386, 4.994432, 4.982762, 
    4.952068, 4.908407, 4.861261, 4.820816, 4.794822, 4.786893, 4.796811, 
    4.82201, 4.859082, 4.904712, 4.956047, 5.010677, 5.066474, 5.121367,
  // momentumY(10,21, 0-49)
    5.263675, 5.267076, 5.260616, 5.245088, 5.221847, 5.192562, 5.159019, 
    5.122997, 5.086214, 5.050299, 5.016766, 4.986938, 4.961788, 4.941614, 
    4.925509, 0, 4.57267, 4.567389, 4.555607, 4.539651, 4.524162, 4.505689, 
    4.496675, 4.498558, 4.514233, 4.543977, 4.587254, 4.642064, 4.705884, 
    4.773979, 4.843802, 4.901035, 4.949372, 4.984136, 5.000959, 4.997036, 
    4.972662, 4.932421, 4.884916, 4.840544, 4.808241, 4.793121, 4.796153, 
    4.815408, 4.847692, 4.889668, 4.938398, 4.991401, 5.046501, 5.101614,
  // momentumY(10,22, 0-49)
    5.271476, 5.27575, 5.269802, 5.254496, 5.231293, 5.201962, 5.168361, 
    5.132299, 5.095483, 5.059496, 5.025783, 4.995612, 4.969961, 4.949296, 
    4.933185, 0, 4.606127, 4.593786, 4.574115, 4.550414, 4.528358, 4.500781, 
    4.48548, 4.482813, 4.495416, 4.523509, 4.566337, 4.621633, 4.686522, 
    4.756358, 4.829571, 4.888551, 4.939791, 4.978797, 5.001094, 5.003343, 
    4.984809, 4.94875, 4.902673, 4.85667, 4.820312, 4.799883, 4.797452, 
    4.8118, 4.840026, 4.878856, 4.925291, 4.976785, 5.031116, 5.086174,
  // momentumY(10,23, 0-49)
    5.276399, 5.281113, 5.275375, 5.260115, 5.236866, 5.207469, 5.173829, 
    5.13778, 5.101011, 5.065071, 5.031356, 5.001098, 4.975291, 4.954518, 
    4.93868, 0, 4.630615, 4.613832, 4.58922, 4.560673, 4.534565, 4.500163, 
    4.480029, 4.473634, 4.483511, 4.509951, 4.552076, 4.607405, 4.672744, 
    4.743471, 4.818842, 4.878325, 4.930957, 4.972464, 4.998406, 5.005173, 
    4.991349, 4.959182, 4.915194, 4.868976, 4.830346, 4.80637, 4.800004, 
    4.810667, 4.83577, 4.87212, 4.916699, 4.966904, 5.020463, 5.075243,
  // momentumY(10,24, 0-49)
    5.277895, 5.282643, 5.276915, 5.261662, 5.238444, 5.20912, 5.175599, 
    5.139707, 5.103124, 5.067368, 5.033813, 5.003671, 4.977938, 4.957258, 
    4.941692, 0, 4.644578, 4.625749, 4.598795, 4.567974, 4.540061, 4.501756, 
    4.478832, 4.470163, 4.478271, 4.503554, 4.545105, 4.600323, 4.665806, 
    4.736924, 4.813501, 4.87292, 4.926011, 4.96866, 4.996484, 5.005741, 
    4.994654, 4.964887, 4.922336, 4.876217, 4.836404, 4.810391, 4.801668, 
    4.810068, 4.83323, 4.868037, 4.911464, 4.96088, 5.013984, 5.068623,
  // momentumY(10,25, 0-49)
    5.275751, 5.280137, 5.274252, 5.259029, 5.235986, 5.20693, 5.173734, 
    5.138188, 5.10195, 5.066529, 5.033287, 5.003433, 4.977952, 4.957484, 
    4.942075, 0, 4.646362, 4.627713, 4.600918, 4.57033, 4.542782, 4.504051, 
    4.480865, 4.47187, 4.479598, 4.504527, 4.545787, 4.600784, 4.666057, 
    4.736995, 4.813643, 4.872583, 4.925354, 4.967914, 4.995914, 5.005612, 
    4.995152, 4.966033, 4.923948, 4.877962, 4.837917, 4.81139, 4.802017, 
    4.809758, 4.832334, 4.866657, 4.909718, 4.958877, 5.011829, 5.066416,
  // momentumY(10,26, 0-49)
    5.270087, 5.273705, 5.267471, 5.252261, 5.229498, 5.200881, 5.168194, 
    5.133167, 5.097431, 5.062489, 5.029718, 5.00033, 4.975293, 4.955161, 
    4.939804, 0, 4.636261, 4.619933, 4.595723, 4.567776, 4.542617, 4.506954, 
    4.486037, 4.478699, 4.487489, 4.512912, 4.554196, 4.60886, 4.67358, 
    4.743774, 4.819333, 4.877504, 4.92928, 4.970582, 4.997083, 5.005145, 
    4.993102, 4.962729, 4.919972, 4.874004, 4.834575, 4.809024, 4.800726, 
    4.809459, 4.832855, 4.867812, 4.911335, 4.960805, 5.013942, 5.0686,
  // momentumY(10,27, 0-49)
    5.261351, 5.26376, 5.256897, 5.241565, 5.219057, 5.190928, 5.158837, 
    5.124437, 5.089321, 5.054998, 5.022872, 4.994169, 4.969829, 4.950259, 
    4.934984, 0, 4.616155, 4.604306, 4.585077, 4.56209, 4.541208, 4.511642, 
    4.495096, 4.490992, 4.501941, 4.528447, 4.569895, 4.624023, 4.687788, 
    4.756649, 4.829976, 4.887001, 4.937045, 4.975907, 4.999275, 5.003732, 
    4.988097, 4.954829, 4.910524, 4.864675, 4.826832, 4.803771, 4.798227, 
    4.809523, 4.835066, 4.871701, 4.916456, 4.966763, 5.020384, 5.0752,
  // momentumY(10,28, 0-49)
    5.250287, 5.251001, 5.243098, 5.227319, 5.204828, 5.177031, 5.145455, 
    5.111665, 5.077218, 5.043633, 5.012346, 4.984618, 4.961354, 4.942771, 
    4.927911, 0, 4.589266, 4.58401, 4.572131, 4.556344, 4.541521, 4.520256, 
    4.509414, 4.509357, 4.5229, 4.55061, 4.592104, 4.645408, 4.707838, 
    4.774844, 4.844988, 4.900376, 4.947849, 4.983022, 5.001625, 5.000618, 
    4.979618, 4.942165, 4.895842, 4.850533, 4.815399, 4.796301, 4.795027, 
    4.81025, 4.839077, 4.87829, 4.924963, 4.976596, 5.031007, 5.086114,
  // momentumY(10,29, 0-49)
    5.237892, 5.236384, 5.226872, 5.210082, 5.187092, 5.159198, 5.127821, 
    5.094449, 5.060609, 5.027836, 4.997607, 4.971239, 4.949625, 4.9328, 
    4.919292, 0, 4.557674, 4.560971, 4.558987, 4.552932, 4.546215, 4.534846, 
    4.530406, 4.534475, 4.550333, 4.578779, 4.61976, 4.671615, 4.73202, 
    4.796323, 4.862085, 4.914719, 4.958258, 4.988181, 5.000409, 4.992544, 
    4.965331, 4.923674, 4.876193, 4.832937, 4.80229, 4.788859, 4.793301, 
    4.813599, 4.846585, 4.889009, 4.938014, 4.991178, 5.046374, 5.101542,
  // momentumY(10,30, 0-49)
    5.229731, 5.229138, 5.220243, 5.203627, 5.180113, 5.150661, 5.116294, 
    5.078084, 5.037141, 4.994608, 4.951617, 4.909244, 4.868432, 4.829989, 
    4.794954, 4.714292, 4.616234, 4.637926, 4.637839, 4.622587, 4.602194, 
    4.580849, 4.568728, 4.568097, 4.581463, 4.608438, 4.648096, 4.698241, 
    4.756376, 4.817419, 4.877771, 4.926244, 4.964109, 4.986963, 4.99125, 
    4.975613, 4.942276, 4.897612, 4.851018, 4.812195, 4.788252, 4.782269, 
    4.793753, 4.820078, 4.857902, 4.904008, 4.955632, 5.010437, 5.066337, 
    5.121289,
  // momentumY(10,31, 0-49)
    5.219232, 5.216277, 5.205369, 5.187213, 5.162733, 5.132943, 5.098883, 
    5.061612, 5.022202, 4.98176, 4.94143, 4.902367, 4.865702, 4.832438, 
    4.803414, 4.719196, 4.623185, 4.63613, 4.634095, 4.622359, 4.607735, 
    4.594142, 4.588014, 4.591664, 4.607731, 4.635858, 4.675278, 4.723969, 
    4.779628, 4.836938, 4.891286, 4.934981, 4.966794, 4.982536, 4.979336, 
    4.957036, 4.91935, 4.873874, 4.830328, 4.797622, 4.781393, 4.783288, 
    4.801867, 4.834084, 4.87652, 4.926019, 4.979887, 5.035825, 5.091748, 
    5.145588,
  // momentumY(10,32, 0-49)
    5.212204, 5.207666, 5.195166, 5.175536, 5.149817, 5.119109, 5.084501, 
    5.047058, 5.007833, 4.967883, 4.928288, 4.890134, 4.854459, 4.822115, 
    4.793561, 4.715725, 4.631017, 4.635134, 4.631091, 4.622012, 4.61214, 
    4.605616, 4.605232, 4.613331, 4.632458, 4.662114, 4.70151, 4.748676, 
    4.801376, 4.854101, 4.901446, 4.939006, 4.963384, 4.970959, 4.959958, 
    4.931739, 4.891537, 4.847791, 4.809901, 4.785426, 4.77831, 4.788849, 
    4.814866, 4.853093, 4.900144, 4.952962, 5.008929, 5.065755, 5.121329, 
    5.173527,
  // momentumY(10,33, 0-49)
    5.20914, 5.203825, 5.190194, 5.169207, 5.142048, 5.109946, 5.074082, 
    5.035568, 4.995455, 4.954757, 4.914469, 4.875549, 4.838848, 4.804925, 
    4.77372, 4.706617, 4.637273, 4.633828, 4.628059, 4.621222, 4.615577, 
    4.615524, 4.620589, 4.633079, 4.655277, 4.686444, 4.725629, 4.770813, 
    4.819751, 4.866857, 4.906264, 4.936515, 4.952563, 4.951732, 4.933675, 
    4.901386, 4.861358, 4.822259, 4.792506, 4.777924, 4.780762, 4.800201, 
    4.83359, 4.877619, 4.929025, 4.984875, 5.042601, 5.0999, 5.154591, 
    5.204463,
  // momentumY(10,34, 0-49)
    5.210141, 5.204962, 5.190825, 5.168797, 5.140215, 5.106468, 5.068875, 
    5.028635, 4.986836, 4.944474, 4.902484, 4.861712, 4.82285, 4.786231, 
    4.751455, 4.695054, 4.642087, 4.632432, 4.625143, 4.620174, 4.618269, 
    4.623944, 4.634017, 4.650625, 4.67562, 4.707963, 4.746448, 4.788954, 
    4.833173, 4.873645, 4.904438, 4.926645, 4.934232, 4.925783, 4.902545, 
    4.868981, 4.83229, 4.800661, 4.780991, 4.77725, 4.790213, 4.818267, 
    4.858552, 4.907861, 4.963102, 5.021472, 5.080428, 5.137609, 5.190722, 
    5.237449,
  // momentumY(10,35, 0-49)
    5.214813, 5.2108, 5.196992, 5.174516, 5.144845, 5.109542, 5.070085, 
    5.0278, 4.983854, 4.939272, 4.894969, 4.851746, 4.810218, 4.770653, 
    4.732632, 4.684653, 4.646751, 4.632051, 4.62333, 4.619743, 4.620919, 
    4.631336, 4.64574, 4.665937, 4.693183, 4.726111, 4.763205, 4.802227, 
    4.84081, 4.873873, 4.895854, 4.909962, 4.909899, 4.895682, 4.870054, 
    4.838493, 4.808202, 4.78625, 4.777755, 4.784982, 4.807583, 4.843489, 
    4.889846, 4.943633, 5.00196, 5.062129, 5.121593, 5.177893, 5.228593, 
    5.271242,
  // momentumY(10,36, 0-49)
    5.222264, 5.220515, 5.208066, 5.186024, 5.155957, 5.119577, 5.078528, 
    5.03429, 4.988141, 4.941181, 4.894366, 4.848512, 4.804265, 4.76197, 
    4.721433, 4.679046, 4.653185, 4.63448, 4.62433, 4.621491, 4.624862, 
    4.638769, 4.656545, 4.67952, 4.708213, 4.740936, 4.775853, 4.810642, 
    4.842913, 4.868268, 4.881892, 4.888682, 4.882713, 4.865387, 4.840581, 
    4.814148, 4.792623, 4.781571, 4.784374, 4.801928, 4.833148, 4.875787, 
    4.927128, 4.984381, 5.044846, 5.105902, 5.164972, 5.219464, 5.266778, 
    5.30433,
  // momentumY(10,37, 0-49)
    5.231169, 5.232775, 5.222847, 5.202373, 5.172933, 5.13634, 5.094387, 
    5.048704, 5.000711, 4.951622, 4.902481, 4.854186, 4.807487, 4.762895, 
    4.720541, 4.681284, 4.663596, 4.641848, 4.63024, 4.627433, 4.631958, 
    4.647927, 4.667863, 4.692542, 4.721674, 4.753293, 4.785275, 4.815282, 
    4.840997, 4.858955, 4.865395, 4.866431, 4.85696, 4.839487, 4.818485, 
    4.799541, 4.78807, 4.788061, 4.801427, 4.82809, 4.86656, 4.914594, 
    4.969669, 5.029223, 5.090712, 5.15157, 5.209159, 5.260755, 5.303586, 
    5.334973,
  // momentumY(10,38, 0-49)
    5.239892, 5.24584, 5.239644, 5.222045, 5.194521, 5.158906, 5.117092, 
    5.070849, 5.021742, 4.971128, 4.920183, 4.869933, 4.821266, 4.774899, 
    4.73128, 4.693408, 4.680095, 4.656179, 4.643091, 4.639637, 4.644267, 
    4.660845, 4.6816, 4.706756, 4.735232, 4.764845, 4.793278, 4.818267, 
    4.837685, 4.849177, 4.850168, 4.847516, 4.837119, 4.822165, 4.80716, 
    4.796963, 4.795705, 4.805967, 4.828554, 4.862772, 4.906951, 4.958941, 
    5.016412, 5.076992, 5.138256, 5.197663, 5.252513, 5.29996, 5.337116, 
    5.361272,
  // momentumY(10,39, 0-49)
    5.246655, 5.257724, 5.256416, 5.243073, 5.218928, 5.18572, 5.145367, 
    5.099737, 5.050538, 4.999286, 4.947315, 4.895807, 4.845814, 4.798248, 
    4.753822, 4.71631, 4.704317, 4.678978, 4.664438, 4.659803, 4.663629, 
    4.679513, 4.699796, 4.724214, 4.750978, 4.777809, 4.802306, 4.822383, 
    4.83622, 4.842612, 4.840141, 4.835948, 4.826879, 4.816355, 4.808491, 
    4.8072, 4.815392, 4.83454, 4.864683, 4.904767, 4.953069, 5.007549, 
    5.066037, 5.126289, 5.185953, 5.242501, 5.293189, 5.335102, 5.365329, 
    5.381271,
  // momentumY(10,40, 0-49)
    5.249744, 5.266394, 5.270947, 5.263197, 5.243958, 5.214726, 5.177338, 
    5.133704, 5.085651, 5.034855, 4.982824, 4.930913, 4.880349, 4.832219, 
    4.787439, 4.749863, 4.737173, 4.711016, 4.69513, 4.68898, 4.691325, 
    4.705497, 4.724216, 4.746839, 4.771021, 4.794501, 4.81493, 4.830498, 
    4.839759, 4.842586, 4.838536, 4.834641, 4.828501, 4.823401, 4.822832, 
    4.829747, 4.846045, 4.872379, 4.908298, 4.952549, 5.003408, 5.058919, 
    5.117007, 5.175501, 5.232083, 5.284229, 5.329195, 5.364105, 5.386174, 
    5.393111,
  // momentumY(10,41, 0-49)
    5.247719, 5.269979, 5.281053, 5.280043, 5.267168, 5.243511, 5.210688, 
    5.170568, 5.125053, 5.075967, 5.024994, 4.973671, 4.923398, 4.875422, 
    4.830817, 4.79321, 4.778804, 4.752316, 4.735268, 4.727466, 4.727908, 
    4.739669, 4.756018, 4.776052, 4.797035, 4.816849, 4.833313, 4.844961, 
    4.85074, 4.851439, 4.847338, 4.845059, 4.842711, 4.843216, 4.849365, 
    4.863264, 4.886032, 4.917758, 4.95768, 5.004436, 5.056305, 5.111372, 
    5.167601, 5.222831, 5.274746, 5.320846, 5.358463, 5.384906, 5.397736, 
    5.395216,
  // momentumY(10,42, 0-49)
    5.239619, 5.267014, 5.284798, 5.291317, 5.286037, 5.269451, 5.242799, 
    5.207787, 5.166325, 5.120343, 5.071693, 5.02209, 4.973096, 4.926105, 
    4.88232, 4.845045, 4.828703, 4.802299, 4.784326, 4.774885, 4.773208, 
    4.78215, 4.795608, 4.812541, 4.829976, 4.846041, 4.858818, 4.867209, 
    4.870528, 4.870278, 4.867199, 4.867313, 4.869003, 4.87472, 4.886584, 
    4.906005, 4.933528, 4.968866, 5.01106, 5.058681, 5.109999, 5.1631, 
    5.215928, 5.266298, 5.311891, 5.350265, 5.378949, 5.395628, 5.398466, 
    5.386536,
  // momentumY(10,43, 0-49)
    5.225125, 5.256631, 5.280723, 5.295022, 5.298166, 5.289894, 5.270908, 
    5.242608, 5.206801, 5.165462, 5.120562, 5.073971, 5.027399, 4.982369, 
    4.940185, 4.903838, 4.885886, 4.85994, 4.841307, 4.830328, 4.826455, 
    4.832383, 4.842665, 4.856229, 4.869998, 4.882415, 4.891881, 4.897665, 
    4.899386, 4.899063, 4.897659, 4.900507, 4.90607, 4.916288, 4.932685, 
    4.956121, 4.986723, 5.023946, 5.066707, 5.113532, 5.16267, 5.212178, 
    5.259955, 5.303786, 5.34137, 5.370416, 5.388793, 5.394788, 5.38742, 
    5.366787,
  // momentumY(10,44, 0-49)
    5.204635, 5.238729, 5.268057, 5.289697, 5.30149, 5.302343, 5.292276, 
    5.272214, 5.243718, 5.20869, 5.169145, 5.127045, 5.08421, 5.042264, 
    5.0026, 4.967926, 4.949046, 4.92391, 4.904885, 4.892501, 4.88643, 
    4.88929, 4.896282, 4.906398, 4.916552, 4.925547, 4.932125, 4.93589, 
    4.936687, 4.936886, 4.937493, 4.94312, 4.952159, 4.966044, 4.985777, 
    5.011779, 5.043863, 5.081303, 5.122929, 5.167236, 5.212452, 5.256604, 
    5.297564, 5.333117, 5.361072, 5.379413, 5.386541, 5.381553, 5.364513, 
    5.336632,
  // momentumY(10,45, 0-49)
    5.179212, 5.214012, 5.246877, 5.274645, 5.294554, 5.304733, 5.304421, 
    5.293918, 5.274354, 5.247395, 5.214958, 5.179004, 5.14139, 5.103791, 
    5.067675, 5.035524, 5.016601, 4.992625, 4.973468, 4.959824, 4.951601, 
    4.951439, 4.955157, 4.961893, 4.9686, 4.974474, 4.978585, 4.980832, 
    4.981196, 4.982283, 4.985005, 4.993274, 5.005284, 5.021986, 5.043922, 
    5.071142, 5.103206, 5.139245, 5.178025, 5.218019, 5.257449, 5.294353, 
    5.326642, 5.352213, 5.369123, 5.375821, 5.371424, 5.355994, 5.330694, 
    5.29772,
  // momentumY(10,46, 0-49)
    5.15041, 5.183906, 5.218145, 5.250115, 5.276795, 5.295731, 5.305416, 
    5.305406, 5.296213, 5.27905, 5.255547, 5.227502, 5.196701, 5.164815, 
    5.133346, 5.104626, 5.08668, 5.064239, 5.04522, 5.03049, 5.020214, 
    5.017181, 5.017759, 5.021304, 5.024827, 5.027922, 5.029962, 5.031085, 
    5.031336, 5.033477, 5.038228, 5.048871, 5.063292, 5.081979, 5.10506, 
    5.132253, 5.162891, 5.19597, 5.230196, 5.264036, 5.295753, 5.323472, 
    5.345274, 5.359347, 5.364205, 5.358969, 5.343636, 5.319263, 5.287948, 
    5.25254,
  // momentumY(10,47, 0-49)
    5.119985, 5.150326, 5.183611, 5.217366, 5.248749, 5.275069, 5.294239, 
    5.305062, 5.307268, 5.30139, 5.288529, 5.270121, 5.247734, 5.222944, 
    5.197252, 5.1729, 5.157071, 5.136595, 5.11804, 5.102479, 5.090351, 
    5.084734, 5.082446, 5.08311, 5.083791, 5.084471, 5.08479, 5.085076, 
    5.085362, 5.088531, 5.095047, 5.107666, 5.123862, 5.143695, 5.166904, 
    5.192897, 5.220782, 5.249414, 5.27744, 5.303342, 5.32549, 5.342224, 
    5.351979, 5.353467, 5.345912, 5.329299, 5.304561, 5.273603, 5.239101, 
    5.204047,
  // momentumY(10,48, 0-49)
    5.089595, 5.115337, 5.145545, 5.178566, 5.212147, 5.243782, 5.271115, 
    5.29231, 5.306252, 5.312603, 5.311698, 5.304386, 5.291848, 5.275453, 
    5.25664, 5.23762, 5.225192, 5.207209, 5.189566, 5.173572, 5.159956, 
    5.152224, 5.147508, 5.145734, 5.143994, 5.142636, 5.141529, 5.141139, 
    5.141435, 5.145405, 5.153227, 5.167259, 5.184483, 5.204558, 5.226863, 
    5.250508, 5.274375, 5.297177, 5.317502, 5.333895, 5.344922, 5.349295, 
    5.346019, 5.33458, 5.315123, 5.288604, 5.256801, 5.222151, 5.187412, 
    5.155191,
  // momentumY(10,49, 0-49)
    5.053679, 5.072524, 5.096591, 5.125384, 5.157755, 5.191944, 5.225796, 
    5.257071, 5.283777, 5.304451, 5.318295, 5.325191, 5.325613, 5.320494, 
    5.311103, 5.300251, 5.299141, 5.285053, 5.268355, 5.251288, 5.235315, 
    5.227765, 5.223431, 5.222784, 5.22031, 5.217353, 5.213843, 5.210539, 
    5.206765, 5.208167, 5.214479, 5.229855, 5.247833, 5.267559, 5.287977, 
    5.307836, 5.32576, 5.340317, 5.350102, 5.353841, 5.350516, 5.339516, 
    5.320797, 5.295008, 5.263525, 5.228363, 5.191968, 5.156848, 5.125219, 
    5.098701,
  // momentumY(11,0, 0-49)
    5.173462, 5.206308, 5.240257, 5.272574, 5.300474, 5.321579, 5.334246, 
    5.337715, 5.33208, 5.318138, 5.297173, 5.270765, 5.240604, 5.208375, 
    5.175654, 5.144077, 5.116427, 5.090436, 5.068562, 5.051296, 5.038685, 
    5.030923, 5.027062, 5.026567, 5.028524, 5.032345, 5.037494, 5.043713, 
    5.050945, 5.059712, 5.070448, 5.084126, 5.100892, 5.121141, 5.144976, 
    5.172139, 5.202004, 5.233603, 5.265666, 5.296687, 5.325003, 5.348888, 
    5.366683, 5.376942, 5.378628, 5.371307, 5.355311, 5.331816, 5.302765, 
    5.270608,
  // momentumY(11,1, 0-49)
    5.194742, 5.228152, 5.26071, 5.289646, 5.312393, 5.32699, 5.332311, 
    5.328114, 5.314935, 5.29389, 5.266475, 5.234376, 5.199319, 5.162972, 
    5.126867, 5.092795, 5.064954, 5.037652, 5.015035, 4.997619, 4.985379, 
    4.97889, 4.976613, 4.977965, 4.981647, 4.987005, 4.993341, 5.000309, 
    5.007703, 5.0163, 5.026547, 5.039942, 5.056371, 5.076459, 5.100532, 
    5.128533, 5.160006, 5.194112, 5.229676, 5.265248, 5.299183, 5.329723, 
    5.355093, 5.373639, 5.383974, 5.385177, 5.376961, 5.359829, 5.335091, 
    5.304753,
  // momentumY(11,2, 0-49)
    5.215133, 5.247335, 5.276393, 5.299809, 5.315543, 5.322279, 5.319528, 
    5.307566, 5.287278, 5.259983, 5.227242, 5.190721, 5.152076, 5.112883, 
    5.074576, 5.039062, 5.011899, 4.983998, 4.961249, 4.944171, 4.93268, 
    4.927715, 4.927212, 4.93057, 4.936181, 4.943317, 4.951117, 4.959096, 
    4.966879, 4.975387, 4.985026, 4.997762, 5.013227, 5.032263, 5.055445, 
    5.082962, 5.114574, 5.149624, 5.187086, 5.225627, 5.263697, 5.299596, 
    5.33156, 5.357855, 5.376884, 5.387331, 5.388323, 5.37959, 5.3616, 5.335593,
  // momentumY(11,3, 0-49)
    5.23278, 5.262092, 5.285949, 5.302372, 5.310034, 5.308362, 5.297498, 
    5.278173, 5.251532, 5.218977, 5.182038, 5.142278, 5.101216, 5.060287, 
    5.020789, 4.984736, 4.959036, 4.931108, 4.908727, 4.892389, 4.881948, 
    4.878703, 4.880101, 4.885571, 4.893275, 4.902404, 4.911927, 4.921201, 
    4.929637, 4.9382, 4.947193, 4.959, 4.972971, 4.990158, 5.011407, 
    5.037199, 5.067567, 5.102092, 5.139944, 5.17996, 5.220726, 5.260663, 
    5.298082, 5.331253, 5.358465, 5.378115, 5.388823, 5.389595, 5.380008, 
    5.360395,
  // momentumY(11,4, 0-49)
    5.246124, 5.271151, 5.28868, 5.297393, 5.296728, 5.286824, 5.26838, 
    5.242476, 5.21042, 5.173625, 5.133534, 5.091561, 5.049062, 5.007304, 
    4.967432, 4.931567, 4.908005, 4.880484, 4.858866, 4.843581, 4.83441, 
    4.833011, 4.836378, 4.843999, 4.853899, 4.86519, 4.876671, 4.887522, 
    4.896918, 4.905757, 4.914163, 4.924904, 4.936983, 4.951648, 4.970031, 
    4.992957, 5.020799, 5.053441, 5.090303, 5.130426, 5.172563, 5.215267, 
    5.256948, 5.295912, 5.330392, 5.358579, 5.378705, 5.389174, 5.388783, 
    5.376987,
  // momentumY(11,5, 0-49)
    5.254175, 5.273928, 5.284616, 5.285609, 5.277045, 5.259663, 5.234583, 
    5.203132, 5.1667, 5.126667, 5.08436, 5.041042, 4.997897, 4.956021, 
    4.916396, 4.881262, 4.860361, 4.83355, 4.812981, 4.798963, 4.791189, 
    4.79168, 4.796989, 4.80671, 4.818825, 4.832373, 4.846004, 4.858711, 
    4.86942, 4.878846, 4.88686, 4.896566, 4.906542, 4.918179, 4.932914, 
    4.951959, 4.976102, 5.005606, 5.040208, 5.079185, 5.121468, 5.165733, 
    5.210474, 5.254028, 5.294588, 5.330204, 5.358836, 5.378459, 5.387281, 
    5.384035,
  // momentumY(11,6, 0-49)
    5.256631, 5.270588, 5.274484, 5.268309, 5.25277, 5.229043, 5.198534, 
    5.162709, 5.122982, 5.080671, 5.036992, 4.993062, 4.949906, 4.90846, 
    4.869534, 4.835497, 4.817565, 4.791654, 4.772311, 4.759662, 4.753291, 
    4.755591, 4.762683, 4.77432, 4.788547, 4.804348, 4.820257, 4.835084, 
    4.847507, 4.857955, 4.865939, 4.874877, 4.882786, 4.891138, 4.901649, 
    4.915957, 4.935346, 4.960551, 4.991693, 5.028335, 5.069591, 5.114242, 
    5.160832, 5.2077, 5.252995, 5.294673, 5.33052, 5.358258, 5.375719, 
    5.381134,
  // momentumY(11,7, 0-49)
    5.253899, 5.261981, 5.259573, 5.247164, 5.225865, 5.197128, 5.162515, 
    5.123538, 5.081592, 5.037923, 4.993641, 4.949739, 4.907105, 4.866518, 
    4.828615, 4.795863, 4.780922, 4.756021, 4.737971, 4.726662, 4.721548, 
    4.72541, 4.733949, 4.747142, 4.763211, 4.781125, 4.799346, 4.816528, 
    4.831117, 4.843144, 4.851673, 4.860385, 4.866592, 4.871735, 4.877743, 
    4.88669, 4.900416, 4.920234, 4.94675, 4.979874, 5.018923, 5.062773, 
    5.109976, 5.158839, 5.207454, 5.253706, 5.295303, 5.329849, 5.355006, 
    5.36871,
  // momentumY(11,8, 0-49)
    5.246972, 5.249469, 5.241543, 5.224041, 5.198316, 5.165953, 5.128552, 
    5.087615, 5.044479, 5.000314, 4.956141, 4.912849, 4.871207, 4.831842, 
    4.795206, 4.763745, 4.751428, 4.727627, 4.710842, 4.700696, 4.696517, 
    4.701485, 4.710924, 4.725105, 4.742551, 4.762268, 4.782706, 4.802408, 
    4.81963, 4.83391, 4.843769, 4.853097, 4.858361, 4.860801, 4.86244, 
    4.865728, 4.873104, 4.886553, 4.907292, 4.935679, 4.971288, 5.01309, 
    5.059626, 5.109141, 5.159651, 5.208991, 5.254846, 5.29482, 5.326542, 
    5.347835,
  // momentumY(11,9, 0-49)
    5.237248, 5.234728, 5.222235, 5.200835, 5.17199, 5.1373, 5.09833, 
    5.056515, 5.013119, 4.96924, 4.925823, 4.883679, 4.843467, 4.805668, 
    4.770514, 4.740153, 4.729591, 4.707032, 4.691422, 4.682123, 4.678374, 
    4.683771, 4.693341, 4.707723, 4.725875, 4.746894, 4.769297, 4.791569, 
    4.811847, 4.829095, 4.841227, 4.852277, 4.857747, 4.858494, 4.856425, 
    4.854231, 4.854913, 4.861206, 4.875076, 4.897473, 4.92833, 4.966763, 
    5.011302, 5.060114, 5.111127, 5.162135, 5.210836, 5.254894, 5.292007, 
    5.319999,
  // momentumY(11,10, 0-49)
    5.226325, 5.219534, 5.203464, 5.179299, 5.148501, 5.112608, 5.073096, 
    5.031306, 4.988426, 4.94549, 4.903389, 4.862872, 4.824508, 4.788627, 
    4.755206, 4.725522, 4.715262, 4.694233, 4.679683, 4.670805, 4.666822, 
    4.671776, 4.680524, 4.694141, 4.712152, 4.733792, 4.757727, 4.782455, 
    4.806074, 4.826941, 4.84233, 4.856339, 4.863483, 4.86403, 4.859515, 
    4.852623, 4.846785, 4.845483, 4.851567, 4.866756, 4.891508, 4.925184, 
    4.966353, 5.013109, 5.063296, 5.114656, 5.164914, 5.211822, 5.253187, 
    5.286903,
  // momentumY(11,11, 0-49)
    5.215777, 5.205538, 5.186835, 5.160881, 5.129076, 5.092853, 5.05357, 
    5.01247, 4.970669, 4.929159, 4.888799, 4.850304, 4.814176, 4.780593, 
    4.749253, 4.719546, 4.70758, 4.688578, 4.67502, 4.666077, 4.661113, 
    4.664628, 4.671499, 4.683293, 4.700191, 4.72163, 4.746493, 4.773363, 
    4.800385, 4.825321, 4.844834, 4.86298, 4.873383, 4.875564, 4.870417, 
    4.860304, 4.848796, 4.840018, 4.837758, 4.844696, 4.862033, 4.889554, 
    4.925972, 4.969349, 5.01745, 5.067966, 5.118637, 5.167293, 5.211854, 
    5.250307,
  // momentumY(11,12, 0-49)
    5.206971, 5.194101, 5.173579, 5.146593, 5.114454, 5.078471, 5.039887, 
    4.99986, 4.959449, 4.919629, 4.88126, 4.845059, 4.811492, 4.78062, 
    4.751868, 4.72114, 4.705098, 4.688858, 4.676319, 4.666856, 4.660173, 
    4.661228, 4.665177, 4.674097, 4.688881, 4.709216, 4.734272, 4.762765, 
    4.792983, 4.822137, 4.846368, 4.869545, 4.884646, 4.890373, 4.886761, 
    4.875495, 4.859918, 4.844513, 4.833935, 4.83196, 4.84078, 4.860842, 
    4.891177, 4.929914, 4.974764, 5.023362, 5.073436, 5.12287, 5.169671, 
    5.211904,
  // momentumY(11,13, 0-49)
    5.200899, 5.186135, 5.164429, 5.136922, 5.104827, 5.069341, 5.031617, 
    4.992749, 4.953773, 4.915673, 4.879345, 4.845548, 4.814764, 4.787011, 
    4.761545, 4.728561, 4.7061, 4.693552, 4.682205, 4.671872, 4.662838, 
    4.660499, 4.66059, 4.665687, 4.677411, 4.695735, 4.72017, 4.749611, 
    4.782543, 4.815727, 4.844905, 4.873561, 4.8944, 4.905334, 4.90543, 
    4.895422, 4.878002, 4.857599, 4.839486, 4.828537, 4.828136, 4.839681, 
    4.862757, 4.895705, 4.936254, 4.981984, 5.030586, 5.079952, 5.128131, 
    5.173246,
  // momentumY(11,14, 0-49)
    5.198095, 5.182048, 5.159592, 5.13182, 5.099866, 5.064854, 5.027873, 
    4.989992, 4.952253, 4.915678, 4.881233, 4.849756, 4.82182, 4.797526, 
    4.776157, 4.739671, 4.70902, 4.701211, 4.69137, 4.679989, 4.668147, 
    4.661624, 4.657088, 4.65757, 4.665394, 4.680862, 4.703853, 4.733477, 
    4.768441, 4.805169, 4.839162, 4.873245, 4.9003, 4.917571, 4.923186, 
    4.916782, 4.900061, 4.876922, 4.852844, 4.83361, 4.823883, 4.826264, 
    4.841175, 4.867381, 4.902731, 4.944778, 4.991159, 5.039723, 5.088521, 
    5.135692,
  // momentumY(11,15, 0-49)
    5.198611, 5.181742, 5.158781, 5.130789, 5.098861, 5.064082, 5.027527, 
    4.990268, 4.953382, 4.917949, 4.885024, 4.855564, 4.83031, 4.809587, 
    4.793001, 4.752295, 4.712822, 4.710817, 4.702914, 4.690477, 4.67556, 
    4.664219, 4.654443, 4.649671, 4.652883, 4.664748, 4.685534, 4.714571, 
    4.750784, 4.790377, 4.82878, 4.867803, 4.900972, 4.92504, 4.93734, 
    4.936428, 4.922827, 4.899501, 4.871641, 4.845568, 4.827119, 4.820251, 
    4.826494, 4.845283, 4.874737, 4.912448, 4.955987, 5.003134, 5.051886, 
    5.100367,
  // momentumY(11,16, 0-49)
    5.202085, 5.184723, 5.161361, 5.133057, 5.10091, 5.066013, 5.029459, 
    4.99235, 4.955808, 4.920977, 4.889006, 4.860992, 4.837896, 4.820388, 
    4.808672, 4.76449, 4.717262, 4.722044, 4.716553, 4.703173, 4.685042, 
    4.668344, 4.652804, 4.642239, 4.640246, 4.647893, 4.665833, 4.693597, 
    4.730288, 4.771996, 4.814262, 4.857442, 4.896148, 4.926826, 4.946223, 
    4.951967, 4.943392, 4.922285, 4.893093, 4.862197, 4.836313, 4.820743, 
    4.818316, 4.829373, 4.852494, 4.885402, 4.925627, 4.970856, 5.019004, 
    5.068143,
  // momentumY(11,17, 0-49)
    5.207882, 5.190274, 5.166554, 5.137811, 5.105181, 5.069798, 5.032796, 
    4.995312, 4.95851, 4.923584, 4.891758, 4.864257, 4.842258, 4.826826, 
    4.818871, 4.77463, 4.723094, 4.735348, 4.732672, 4.718445, 4.696949, 
    4.674356, 4.652512, 4.635655, 4.627968, 4.630945, 4.645575, 4.671546, 
    4.708066, 4.751193, 4.796754, 4.843171, 4.886521, 4.923114, 4.949328, 
    4.962093, 4.959697, 4.942693, 4.914481, 4.881027, 4.849508, 4.826371, 
    4.815795, 4.819218, 4.835872, 4.863728, 4.900331, 4.943276, 4.990375, 
    5.039623,
  // momentumY(11,18, 0-49)
    5.215275, 5.197681, 5.173691, 5.144443, 5.111129, 5.074939, 5.037043, 
    4.998607, 4.960812, 4.924872, 4.892043, 4.863613, 4.840909, 4.825321, 
    4.818491, 4.781203, 4.73237, 4.751977, 4.752251, 4.737044, 4.711777, 
    4.682581, 4.653769, 4.630121, 4.616386, 4.614459, 4.625572, 4.649482, 
    4.685395, 4.729392, 4.777759, 4.826488, 4.873441, 4.914927, 4.947153, 
    4.966595, 4.970727, 4.958978, 4.933579, 4.899727, 4.8646, 4.835458, 
    4.817726, 4.814026, 4.824396, 4.847192, 4.880045, 4.920485, 4.966215, 
    5.015142,
  // momentumY(11,19, 0-49)
    5.223647, 5.206471, 5.182448, 5.152765, 5.118663, 5.081373, 5.042089, 
    5.001988, 4.962242, 4.924037, 4.888577, 4.857102, 4.830956, 4.811839, 
    4.802468, 4.782428, 4.748799, 4.774101, 4.776849, 4.759989, 4.72988, 
    4.692934, 4.656215, 4.62528, 4.605374, 4.598666, 4.606437, 4.628368, 
    4.663541, 4.708077, 4.758886, 4.809097, 4.858589, 4.903782, 4.940869, 
    4.966106, 4.976411, 4.9703, 4.948884, 4.916395, 4.87963, 4.846251, 
    4.822695, 4.812732, 4.817303, 4.835267, 4.864427, 4.902291, 4.94647, 
    4.994776,
  // momentumY(11,20, 0-49)
    5.228605, 5.209377, 5.183713, 5.153066, 5.118945, 5.08285, 5.046243, 
    5.010551, 4.977164, 4.947405, 4.922451, 4.903156, 4.889757, 4.881487, 
    4.876232, 0, 4.74619, 4.746288, 4.737542, 4.720608, 4.697607, 4.668127, 
    4.638677, 4.612827, 4.595506, 4.58938, 4.596458, 4.617135, 4.651025, 
    4.694868, 4.746641, 4.79661, 4.846766, 4.893705, 4.933717, 4.963015, 
    4.978206, 4.977147, 4.959987, 4.929938, 4.893122, 4.857208, 4.829299, 
    4.814166, 4.813659, 4.827224, 4.852918, 4.888282, 4.930861, 4.978384,
  // momentumY(11,21, 0-49)
    5.2353, 5.216488, 5.190962, 5.160259, 5.125952, 5.089577, 5.052596, 
    5.016393, 4.982272, 4.951435, 4.92492, 4.903454, 4.887238, 4.875626, 
    4.866798, 0, 4.797721, 4.792305, 4.77688, 4.75208, 4.720561, 4.678942, 
    4.639472, 4.605354, 4.581752, 4.571404, 4.576097, 4.595869, 4.629888, 
    4.674782, 4.72919, 4.780305, 4.832267, 4.881819, 4.925358, 4.959108, 
    4.979494, 4.983882, 4.97161, 4.944922, 4.909168, 4.871809, 4.840419, 
    4.820678, 4.815356, 4.824558, 4.846657, 4.879263, 4.919861, 4.966089,
  // momentumY(11,22, 0-49)
    5.239971, 5.221348, 5.19583, 5.165015, 5.130526, 5.093925, 5.056665, 
    5.020096, 4.985459, 4.95387, 4.926275, 4.903344, 4.885296, 4.871654, 
    4.860947, 0, 4.835303, 4.825794, 4.806291, 4.777096, 4.740961, 4.690882, 
    4.644479, 4.604306, 4.575753, 4.561767, 4.564087, 4.582548, 4.615982, 
    4.660958, 4.716836, 4.767711, 4.819979, 4.870557, 4.915993, 4.952604, 
    4.976768, 4.985557, 4.977713, 4.954643, 4.920895, 4.883494, 4.850173, 
    4.82724, 4.818252, 4.823944, 4.84304, 4.873272, 4.912107, 4.957114,
  // momentumY(11,23, 0-49)
    5.242476, 5.223934, 5.198411, 5.167542, 5.132972, 5.096276, 5.058898, 
    5.022161, 4.987256, 4.95525, 4.927035, 4.903254, 4.884159, 4.869406, 
    4.857812, 0, 4.860757, 4.848539, 4.826694, 4.795172, 4.756673, 4.700799, 
    4.649669, 4.605175, 4.572934, 4.556139, 4.556563, 4.573909, 4.606749, 
    4.651597, 4.708432, 4.75862, 4.810601, 4.861441, 4.90783, 4.9462, 
    4.97295, 4.984998, 4.980686, 4.960799, 4.929197, 4.892447, 4.858245, 
    4.833289, 4.82172, 4.824795, 4.841565, 4.869889, 4.907241, 4.951149,
  // momentumY(11,24, 0-49)
    5.242755, 5.224256, 5.198783, 5.167976, 5.133484, 5.096869, 5.059566, 
    5.022881, 4.987978, 4.955898, 4.927505, 4.903431, 4.883943, 4.868771, 
    4.856884, 0, 4.873823, 4.860311, 4.837456, 4.80504, 4.765738, 4.706779, 
    4.653216, 4.606438, 4.572193, 4.55386, 4.553253, 4.570012, 4.602548, 
    4.647337, 4.704798, 4.75439, 4.805976, 4.856723, 4.903411, 4.942552, 
    4.970578, 4.984347, 4.981996, 4.963964, 4.933707, 4.897477, 4.862895, 
    4.836847, 4.823806, 4.825346, 4.840734, 4.867923, 4.904401, 4.947665,
  // momentumY(11,25, 0-49)
    5.240794, 5.22232, 5.196975, 5.166369, 5.132127, 5.095788, 5.058773, 
    5.022375, 4.987755, 4.955944, 4.927806, 4.903964, 4.884675, 4.869664, 
    4.8579, 0, 4.873703, 4.860322, 4.837665, 4.805562, 4.766716, 4.707583, 
    4.654046, 4.607269, 4.572984, 4.554605, 4.553962, 4.570693, 4.603181, 
    4.647916, 4.705504, 4.754699, 4.80592, 4.856369, 4.902862, 4.941946, 
    4.970081, 4.984127, 4.982181, 4.964595, 4.934705, 4.898656, 4.864019, 
    4.837709, 4.824278, 4.825392, 4.84038, 4.86723, 4.903439, 4.946502,
  // momentumY(11,26, 0-49)
    5.236609, 5.218122, 5.192966, 5.162689, 5.128861, 5.092988, 5.056469, 
    5.020595, 4.98654, 4.955349, 4.927902, 4.904818, 4.886321, 4.872047, 
    4.860817, 0, 4.860604, 4.848742, 4.827468, 4.796851, 4.759639, 4.703284, 
    4.652233, 4.607754, 4.575406, 4.558476, 4.558778, 4.576014, 4.608685, 
    4.653347, 4.710508, 4.75958, 4.810529, 4.860532, 4.90638, 4.944607, 
    4.971689, 4.984544, 4.981393, 4.962756, 4.932151, 4.895843, 4.8614, 
    4.835618, 4.82288, 4.824695, 4.8403, 4.867644, 4.904226, 4.947563,
  // momentumY(11,27, 0-49)
    5.230247, 5.211652, 5.186687, 5.156816, 5.12353, 5.088286, 5.052456, 
    5.017334, 4.984122, 4.953905, 4.927598, 4.90583, 4.888774, 4.875917, 
    4.8658, 0, 4.835612, 4.826562, 4.807929, 4.780112, 4.745865, 4.695104, 
    4.648843, 4.608716, 4.580005, 4.565769, 4.567803, 4.585944, 4.618935, 
    4.663445, 4.719617, 4.768734, 4.819421, 4.868762, 4.913473, 4.950031, 
    4.97492, 4.985185, 4.979329, 4.958301, 4.926076, 4.889226, 4.855335, 
    4.83092, 4.819949, 4.823555, 4.84074, 4.869361, 4.906916, 4.950954,
  // momentumY(11,28, 0-49)
    5.221816, 5.202913, 5.178044, 5.148566, 5.115879, 5.081367, 5.046379, 
    5.012208, 4.980105, 4.951216, 4.926524, 4.906692, 4.891847, 4.881296, 
    4.873246, 0, 4.800921, 4.795757, 4.781104, 4.757642, 4.728002, 4.685359, 
    4.64586, 4.611671, 4.58779, 4.577054, 4.5813, 4.600579, 4.633968, 
    4.678254, 4.733004, 4.782204, 4.832494, 4.880813, 4.923745, 4.957682, 
    4.979128, 4.985353, 4.975339, 4.950729, 4.91621, 4.878789, 4.846007, 
    4.823902, 4.815784, 4.822229, 4.841906, 4.872549, 4.91166, 4.956846,
  // momentumY(11,29, 0-49)
    5.211528, 5.191969, 5.166947, 5.13771, 5.105555, 5.071788, 5.037718, 
    5.004653, 4.97389, 4.946674, 4.924098, 4.906909, 4.895241, 4.888247, 
    4.883862, 0, 4.758096, 4.757624, 4.74851, 4.73148, 4.7087, 4.676564, 
    4.645609, 4.618504, 4.600053, 4.593021, 4.59944, 4.61967, 4.653188, 
    4.696864, 4.749561, 4.798358, 4.847646, 4.894192, 4.934445, 4.964732, 
    4.981649, 4.982831, 4.967932, 4.939481, 4.902971, 4.865784, 4.835213, 
    4.816581, 4.812366, 4.8225, 4.845302, 4.8784, 4.919327, 4.965767,
  // momentumY(11,30, 0-49)
    5.203184, 5.185256, 5.161644, 5.13331, 5.101258, 5.066503, 5.030076, 
    4.993026, 4.956442, 4.921446, 4.889181, 4.860801, 4.837526, 4.82086, 
    4.81322, 4.793564, 4.759291, 4.783369, 4.786592, 4.771524, 4.744068, 
    4.707412, 4.671654, 4.641252, 4.621176, 4.613644, 4.620066, 4.640306, 
    4.673593, 4.716428, 4.766704, 4.814546, 4.862028, 4.905797, 4.942236, 
    4.967708, 4.97907, 4.974526, 4.954614, 4.922864, 4.885518, 4.850087, 
    4.823308, 4.809544, 4.810329, 4.82495, 4.851427, 4.887334, 4.930273, 
    4.978027,
  // momentumY(11,31, 0-49)
    5.191897, 5.173043, 5.149139, 5.121112, 5.08991, 5.056485, 5.021814, 
    4.986914, 4.952852, 4.920757, 4.891789, 4.867128, 4.847923, 4.835331, 
    4.830701, 4.793941, 4.74672, 4.765321, 4.765812, 4.751783, 4.728415, 
    4.699248, 4.671027, 4.647578, 4.633379, 4.630328, 4.639804, 4.661777, 
    4.695667, 4.737928, 4.785717, 4.832349, 4.877781, 4.918511, 4.950845, 
    4.971227, 4.976875, 4.966708, 4.942261, 4.908067, 4.87096, 4.838338, 
    4.81617, 4.807773, 4.813767, 4.832868, 4.862859, 4.901292, 4.945847, 
    4.994394,
  // momentumY(11,32, 0-49)
    5.182117, 5.162619, 5.138494, 5.110645, 5.079966, 5.047355, 5.013735, 
    4.980078, 4.947419, 4.916849, 4.889486, 4.866421, 4.848642, 4.836962, 
    4.832007, 4.788759, 4.739945, 4.751895, 4.749567, 4.736239, 4.716129, 
    4.69341, 4.671788, 4.654728, 4.646223, 4.647764, 4.660519, 4.684406, 
    4.718903, 4.760376, 4.805366, 4.850052, 4.892422, 4.928905, 4.955868, 
    4.970041, 4.969263, 4.95342, 4.925176, 4.889977, 4.854934, 4.826926, 
    4.810857, 4.808888, 4.820767, 4.844739, 4.87844, 4.919459, 4.965571, 
    5.014742,
  // momentumY(11,33, 0-49)
    5.174572, 5.154589, 5.13018, 5.102248, 5.071674, 5.039321, 5.00607, 
    4.972849, 4.940649, 4.910503, 4.883449, 4.860447, 4.842265, 4.829318, 
    4.82152, 4.779136, 4.735283, 4.740807, 4.736142, 4.723701, 4.706699, 
    4.689884, 4.674292, 4.663169, 4.660039, 4.665985, 4.681876, 4.707491, 
    4.742249, 4.782453, 4.824167, 4.866026, 4.904251, 4.935326, 4.955851, 
    4.96308, 4.955732, 4.934846, 4.90422, 4.869962, 4.83904, 4.817427, 
    4.808751, 4.814018, 4.832221, 4.861261, 4.898711, 4.942233, 4.989711, 
    5.039204,
  // momentumY(11,34, 0-49)
    5.170084, 5.149796, 5.125022, 5.096713, 5.065773, 5.033074, 4.999493, 
    4.965929, 4.933328, 4.902668, 4.874899, 4.850855, 4.831088, 4.815667, 
    4.803902, 4.766072, 4.730641, 4.730635, 4.724333, 4.713195, 4.699438, 
    4.68818, 4.678235, 4.672667, 4.674529, 4.684519, 4.703167, 4.730061, 
    4.764484, 4.802741, 4.840598, 4.878656, 4.91169, 4.936383, 4.949773, 
    4.949892, 4.936552, 4.912015, 4.881037, 4.849986, 4.825233, 4.811538, 
    4.81119, 4.824152, 4.848831, 4.882911, 4.923972, 4.969772, 5.0183, 
    5.067683,
  // momentumY(11,35, 0-49)
    5.16936, 5.149054, 5.123928, 5.095007, 5.063273, 5.029659, 4.99507, 
    4.960418, 4.926631, 4.894642, 4.865333, 4.839435, 4.817364, 4.798974, 
    4.783234, 4.750862, 4.725138, 4.7207, 4.713482, 4.704073, 4.693744, 
    4.687737, 4.683125, 4.682759, 4.689171, 4.702719, 4.723572, 4.751113, 
    4.784435, 4.819942, 4.853301, 4.886603, 4.913572, 4.931258, 4.937376, 
    4.930943, 4.912982, 4.886868, 4.857957, 4.832395, 4.815557, 4.810833, 
    4.819266, 4.839981, 4.870982, 4.909855, 4.954227, 5.001952, 5.051094, 
    5.099827,
  // momentumY(11,36, 0-49)
    5.172808, 5.152929, 5.127627, 5.098027, 5.065219, 5.030244, 4.994094, 
    4.95773, 4.922098, 4.888113, 4.856624, 4.828312, 4.803537, 4.782102, 
    4.762949, 4.735329, 4.718907, 4.711125, 4.703607, 4.696209, 4.689353, 
    4.688214, 4.688584, 4.693012, 4.703455, 4.719961, 4.742342, 4.769779, 
    4.801148, 4.833087, 4.861357, 4.889116, 4.909484, 4.920085, 4.919499, 
    4.907862, 4.887349, 4.862151, 4.837749, 4.819602, 4.811847, 4.816537, 
    4.833683, 4.861814, 4.898704, 4.941922, 4.989157, 5.038332, 5.08755, 
    5.134997,
  // momentumY(11,37, 0-49)
    5.180398, 5.161556, 5.136457, 5.106329, 5.072402, 5.035862, 4.997823, 
    4.959341, 4.921418, 4.884993, 4.850913, 4.819863, 4.792229, 4.767898, 
    4.746009, 4.72179, 4.713002, 4.702868, 4.695462, 4.6901, 4.686528, 
    4.689706, 4.694558, 4.703251, 4.717091, 4.735848, 4.758998, 4.785535, 
    4.814129, 4.841794, 4.864573, 4.886342, 4.900098, 4.904203, 4.898227, 
    4.883398, 4.862806, 4.841026, 4.823173, 4.813704, 4.815465, 4.829372, 
    4.854675, 4.889541, 4.931647, 4.978592, 5.028115, 5.07816, 5.126826, 
    5.172269,
  // momentumY(11,38, 0-49)
    5.191592, 5.174534, 5.150224, 5.119972, 5.085162, 5.047144, 5.007191, 
    4.966487, 4.926123, 4.887098, 4.850299, 4.816452, 4.786022, 4.759057, 
    4.735008, 4.712789, 4.70924, 4.697576, 4.690451, 4.686867, 4.686113, 
    4.692836, 4.701461, 4.713706, 4.730173, 4.750387, 4.773516, 4.798402, 
    4.82355, 4.846487, 4.86371, 4.879532, 4.88728, 4.886151, 4.876693, 
    4.861042, 4.842818, 4.826513, 4.816519, 4.816159, 4.827136, 4.849496, 
    4.882006, 4.922656, 4.969118, 5.019029, 5.070147, 5.120387, 5.167787, 
    5.210437,
  // momentumY(11,39, 0-49)
    5.205347, 5.190912, 5.168145, 5.138416, 5.103247, 5.064161, 5.022605, 
    4.979915, 4.937297, 4.895839, 4.856494, 4.820059, 4.787104, 4.757856, 
    4.732081, 4.710703, 4.709868, 4.697269, 4.690359, 4.688056, 4.689408, 
    4.698699, 4.710176, 4.72507, 4.743271, 4.764093, 4.786444, 4.809061, 
    4.830353, 4.848471, 4.860497, 4.870972, 4.873897, 4.869296, 4.858545, 
    4.844366, 4.830497, 4.82097, 4.819266, 4.827655, 4.846931, 4.876558, 
    4.915043, 4.960332, 5.010135, 5.06212, 5.114024, 5.163682, 5.209023, 
    5.248034,
  // momentumY(11,40, 0-49)
    5.220186, 5.209238, 5.188896, 5.160541, 5.125803, 5.086365, 5.043848, 
    4.999744, 4.955394, 4.911988, 4.870568, 4.832009, 4.796983, 4.765884, 
    4.73874, 4.717393, 4.717087, 4.703911, 4.69698, 4.695314, 4.697904, 
    4.708665, 4.721914, 4.738419, 4.75739, 4.777978, 4.798889, 4.81882, 
    4.836173, 4.849782, 4.857394, 4.863602, 4.863284, 4.857172, 4.847208, 
    4.836345, 4.828079, 4.825771, 4.831997, 4.848148, 4.874382, 4.90982, 
    4.95287, 5.001508, 5.053501, 5.106535, 5.158285, 5.206468, 5.248866, 
    5.283354,
  // momentumY(11,41, 0-49)
    5.23431, 5.227661, 5.210699, 5.184736, 5.151451, 5.112651, 5.070111, 
    5.025473, 4.980214, 4.935633, 4.892861, 4.852852, 4.816367, 4.783926, 
    4.755749, 4.733974, 4.732622, 4.719017, 4.711739, 4.710033, 4.712957, 
    4.724083, 4.737983, 4.755019, 4.773808, 4.793388, 4.812348, 4.829412, 
    4.84305, 4.852812, 4.85709, 4.860407, 4.858553, 4.852761, 4.845245, 
    4.838876, 4.836684, 4.841298, 4.854504, 4.87704, 4.908657, 4.948308, 
    4.994401, 5.044983, 5.097881, 5.150779, 5.201279, 5.246957, 5.285442, 
    5.314502,
  // momentumY(11,42, 0-49)
    5.245757, 5.244094, 5.231469, 5.209024, 5.178406, 5.141475, 5.100114, 
    5.056091, 5.011003, 4.966255, 4.923054, 4.882427, 4.845201, 4.811985, 
    4.783129, 4.76075, 4.75743, 4.7434, 4.735441, 4.733069, 4.735492, 
    4.745985, 4.759491, 4.776057, 4.793811, 4.811748, 4.828418, 4.84264, 
    4.853035, 4.859815, 4.861965, 4.863824, 4.861996, 4.857988, 4.854019, 
    4.852657, 4.856369, 4.867102, 4.886012, 4.913383, 4.948726, 4.99094, 
    5.038484, 5.089493, 5.141856, 5.193256, 5.241224, 5.283213, 5.316723, 
    5.33947,
  // momentumY(11,43, 0-49)
    5.252583, 5.256382, 5.248981, 5.231237, 5.20464, 5.171007, 5.132254, 
    5.090226, 5.046606, 5.002879, 4.96032, 4.92001, 4.882821, 4.849424, 
    4.820261, 4.797302, 4.791629, 4.777101, 4.768164, 4.764614, 4.765842, 
    4.774894, 4.787142, 4.802403, 4.818435, 4.834261, 4.848473, 4.860041, 
    4.867776, 4.872492, 4.873652, 4.875337, 4.87478, 4.873552, 4.873688, 
    4.877326, 4.886364, 4.902164, 4.925396, 4.95604, 4.993475, 5.036603, 
    5.083958, 5.133768, 5.18399, 5.232327, 5.276277, 5.313229, 5.340635, 
    5.356261,
  // momentumY(11,44, 0-49)
    5.253074, 5.262515, 5.261069, 5.249179, 5.228035, 5.199276, 5.164745, 
    5.12628, 5.085594, 5.044218, 5.003467, 4.964456, 4.928098, 4.895112, 
    4.866016, 4.842618, 4.834599, 4.819472, 4.809327, 4.804217, 4.803734, 
    4.810767, 4.821117, 4.834463, 4.848287, 4.861711, 4.873432, 4.882618, 
    4.888287, 4.891765, 4.892875, 4.89539, 4.896967, 4.89908, 4.90345, 
    4.911751, 4.925344, 4.945101, 4.971322, 5.003768, 5.041742, 5.084168, 
    5.129661, 5.176544, 5.222858, 5.266371, 5.304625, 5.335056, 5.355216, 
    5.363077,
  // momentumY(11,45, 0-49)
    5.245976, 5.260865, 5.26584, 5.260825, 5.246549, 5.224311, 5.19573, 
    5.162527, 5.126361, 5.08875, 5.05102, 5.014307, 4.97956, 4.947553, 
    4.918889, 4.895254, 4.885153, 4.869344, 4.85784, 4.850928, 4.848397, 
    4.853063, 4.861111, 4.872155, 4.883486, 4.894375, 4.903677, 4.910774, 
    4.914892, 4.917789, 4.919525, 4.923557, 4.927764, 4.933413, 4.941857, 
    4.954303, 4.971632, 4.994293, 5.02229, 5.055206, 5.092278, 5.13245, 
    5.174401, 5.216556, 5.257073, 5.293852, 5.324604, 5.34698, 5.358833, 
    5.358551,
  // momentumY(11,46, 0-49)
    5.230698, 5.250425, 5.261923, 5.264531, 5.258378, 5.244246, 5.223355, 
    5.197155, 5.167138, 5.134735, 5.101245, 5.067813, 5.035434, 5.004955, 
    4.977088, 4.953472, 4.941727, 4.925207, 4.912287, 4.903466, 4.898721, 
    4.900876, 4.90643, 4.914997, 4.923724, 4.932077, 4.939089, 4.944373, 
    4.94734, 4.950113, 4.952881, 4.958815, 4.965834, 4.974938, 4.987098, 
    5.003079, 5.023328, 5.047932, 5.076622, 5.108816, 5.143669, 5.180115, 
    5.216885, 5.252507, 5.285301, 5.313405, 5.334856, 5.347742, 5.35046, 
    5.342037,
  // momentumY(11,47, 0-49)
    5.207477, 5.23103, 5.248695, 5.259253, 5.262141, 5.257459, 5.24584, 
    5.228285, 5.205985, 5.18019, 5.152124, 5.122934, 5.093671, 5.065282, 
    5.03861, 5.015327, 5.00253, 4.985361, 4.971079, 4.96038, 4.953408, 
    4.953086, 4.956131, 4.962209, 4.968366, 4.974279, 4.979176, 4.982888, 
    4.984988, 4.987902, 4.991867, 4.999817, 5.009564, 5.021826, 5.037194, 
    5.056029, 5.07839, 5.104032, 5.132427, 5.162814, 5.194239, 5.225595, 
    5.255641, 5.283024, 5.306286, 5.323929, 5.334507, 5.336784, 5.329955, 
    5.313877,
  // momentumY(11,48, 0-49)
    5.177426, 5.203481, 5.226476, 5.244749, 5.257052, 5.262691, 5.261548, 
    5.253999, 5.240782, 5.222868, 5.201346, 5.177341, 5.151967, 5.126286, 
    5.101289, 5.078762, 5.06565, 5.04801, 5.03255, 5.020142, 5.011084, 
    5.008462, 5.009127, 5.012832, 5.016562, 5.020209, 5.023188, 5.025537, 
    5.026949, 5.030105, 5.035226, 5.045074, 5.057245, 5.072175, 5.090107, 
    5.111032, 5.134658, 5.16043, 5.187572, 5.215123, 5.242, 5.267024, 
    5.288981, 5.30666, 5.318905, 5.324718, 5.323361, 5.314494, 5.298303, 
    5.275572,
  // momentumY(11,49, 0-49)
    5.130487, 5.157133, 5.184359, 5.21029, 5.233043, 5.250996, 5.26301, 
    5.268517, 5.267499, 5.260395, 5.247995, 5.231311, 5.211483, 5.189702, 
    5.167173, 5.146682, 5.140685, 5.122538, 5.104847, 5.089356, 5.0769, 
    5.074059, 5.074942, 5.079597, 5.082418, 5.084044, 5.083921, 5.082497, 
    5.079126, 5.079224, 5.082874, 5.095003, 5.110043, 5.128022, 5.148745, 
    5.171737, 5.196276, 5.221437, 5.24613, 5.269165, 5.289305, 5.305318, 
    5.316079, 5.32065, 5.318389, 5.309089, 5.293078, 5.271255, 5.245065, 
    5.216325,
  // momentumY(12,0, 0-49)
    5.283156, 5.303393, 5.315825, 5.319623, 5.31465, 5.301387, 5.280786, 
    5.254111, 5.222781, 5.188264, 5.151982, 5.115261, 5.079288, 5.045088, 
    5.013504, 4.985375, 4.962522, 4.942296, 4.926528, 4.915215, 4.908121, 
    4.905272, 4.90585, 4.909438, 4.915286, 4.922814, 4.93137, 4.940413, 
    4.949502, 4.958674, 4.967987, 4.978175, 4.989471, 5.002637, 5.018452, 
    5.037585, 5.060488, 5.087313, 5.117883, 5.15169, 5.18792, 5.225489, 
    5.263074, 5.299156, 5.332043, 5.359944, 5.381062, 5.393738, 5.396669, 
    5.389134,
  // momentumY(12,1, 0-49)
    5.289672, 5.306209, 5.313846, 5.31217, 5.301459, 5.28255, 5.256652, 
    5.225194, 5.189679, 5.15159, 5.112332, 5.073187, 5.035285, 4.999592, 
    4.966884, 4.938138, 4.916506, 4.896032, 4.880301, 4.86932, 4.862805, 
    4.861174, 4.863127, 4.868292, 4.875661, 4.884639, 4.894459, 4.904496, 
    4.91414, 4.923573, 4.932739, 4.942745, 4.953437, 4.965678, 4.980408, 
    4.998491, 5.020582, 5.047031, 5.077825, 5.112586, 5.150586, 5.19079, 
    5.231888, 5.272332, 5.310356, 5.344034, 5.371366, 5.390417, 5.399523, 
    5.397548,
  // momentumY(12,2, 0-49)
    5.289351, 5.301156, 5.303457, 5.296273, 5.280246, 5.256473, 5.226311, 
    5.191248, 5.152781, 5.112347, 5.071281, 5.030792, 4.991937, 4.955608, 
    4.922512, 4.893762, 4.873818, 4.853418, 4.837952, 4.827422, 4.821506, 
    4.821013, 4.824201, 4.830774, 4.839534, 4.849892, 4.860994, 4.872135, 
    4.882534, 4.892459, 4.901697, 4.911676, 4.921791, 4.932947, 4.946202, 
    4.962606, 4.983036, 5.008065, 5.037891, 5.072294, 5.110664, 5.152039, 
    5.195147, 5.238437, 5.280128, 5.318251, 5.350725, 5.375486, 5.390674, 
    5.394858,
  // momentumY(12,3, 0-49)
    5.282612, 5.289087, 5.285932, 5.273549, 5.252862, 5.225129, 5.191766, 
    5.154241, 5.113979, 5.072326, 5.030522, 4.989674, 4.950751, 4.914566, 
    4.881744, 4.85353, 4.835714, 4.815639, 4.800602, 4.790585, 4.785224, 
    4.785729, 4.789946, 4.797691, 4.807655, 4.819279, 4.831649, 4.843991, 
    4.855368, 4.866057, 4.875648, 4.885847, 4.895519, 4.905539, 4.917031, 
    4.931207, 4.949178, 4.971781, 4.999463, 5.032219, 5.069589, 5.110712, 
    5.154368, 5.199042, 5.24297, 5.2842, 5.320669, 5.350304, 5.37118, 5.381702,
  // momentumY(12,4, 0-49)
    5.270433, 5.271401, 5.263016, 5.245987, 5.221428, 5.190666, 5.15511, 
    5.116154, 5.07512, 5.033241, 4.991632, 4.951296, 4.9131, 4.877757, 
    4.845793, 4.818586, 4.803279, 4.783717, 4.769216, 4.759707, 4.754789, 
    4.756079, 4.761035, 4.769634, 4.780541, 4.793252, 4.806829, 4.820447, 
    4.833023, 4.844786, 4.855074, 4.865842, 4.87534, 4.884321, 4.893908, 
    4.905432, 4.92024, 4.93947, 4.963875, 4.993721, 5.02876, 5.068261, 
    5.111091, 5.155785, 5.200624, 5.243716, 5.283067, 5.316677, 5.342657, 
    5.359342,
  // momentumY(12,5, 0-49)
    5.254186, 5.249829, 5.236703, 5.215734, 5.188132, 5.155237, 5.118395, 
    5.078903, 5.037965, 4.996687, 4.956069, 4.916993, 4.880211, 4.84632, 
    4.815726, 4.789899, 4.777379, 4.758461, 4.744543, 4.735467, 4.730793, 
    4.732566, 4.737878, 4.74691, 4.758401, 4.771935, 4.786589, 4.801508, 
    4.815494, 4.828657, 4.840042, 4.851838, 4.861586, 4.869823, 4.877574, 
    4.886226, 4.897335, 4.912361, 4.932431, 4.958163, 4.989584, 5.026161, 
    5.066878, 5.110339, 5.154894, 5.19872, 5.239929, 5.276628, 5.30701, 
    5.329417,
  // momentumY(12,6, 0-49)
    5.235466, 5.226234, 5.209022, 5.184886, 5.155065, 5.120851, 5.083508, 
    5.044224, 5.004089, 4.964089, 4.925107, 4.88791, 4.853123, 4.821205, 
    4.792401, 4.768209, 4.758565, 4.740386, 4.727033, 4.718237, 4.713521, 
    4.715374, 4.720548, 4.729478, 4.741088, 4.755076, 4.770578, 4.786751, 
    4.802309, 4.817187, 4.830103, 4.84348, 4.854072, 4.862099, 4.868368, 
    4.874223, 4.881364, 4.891574, 4.906406, 4.926915, 4.953505, 4.985915, 
    5.023302, 5.064378, 5.107562, 5.151116, 5.193247, 5.232182, 5.266211, 
    5.293715,
  // momentumY(12,7, 0-49)
    5.215919, 5.202434, 5.181869, 5.155337, 5.124051, 5.089231, 5.052039, 
    5.013558, 4.974773, 4.936571, 4.899731, 4.864904, 4.832586, 4.803066, 
    4.776391, 4.753929, 4.746964, 4.729606, 4.716753, 4.708011, 4.702882, 
    4.704314, 4.708754, 4.716944, 4.728096, 4.742053, 4.758061, 4.775326, 
    4.792534, 4.809388, 4.824256, 4.839813, 4.851985, 4.860579, 4.86606, 
    4.869582, 4.872879, 4.878002, 4.88695, 4.901301, 4.921952, 4.949025, 
    4.981931, 5.019534, 5.060344, 5.102702, 5.144898, 5.185256, 5.222154, 
    5.254018,
  // momentumY(12,8, 0-49)
    5.197084, 5.180053, 5.15687, 5.128651, 5.096552, 5.0617, 5.02516, 
    4.987918, 4.950877, 4.914841, 4.880503, 4.848413, 4.818925, 4.792144, 
    4.76786, 4.747036, 4.742175, 4.725766, 4.713326, 4.70436, 4.698389, 
    4.698829, 4.701871, 4.708604, 4.71863, 4.731961, 4.748012, 4.766073, 
    4.784878, 4.803852, 4.82102, 4.839316, 4.853869, 4.863999, 4.869711, 
    4.871802, 4.871869, 4.872107, 4.874922, 4.882471, 4.896258, 4.916928, 
    4.944264, 4.977354, 5.014838, 5.055129, 5.096582, 5.137584, 5.17657, 
    5.212003,
  // momentumY(12,9, 0-49)
    5.180264, 5.160401, 5.13527, 5.105958, 5.07355, 5.03908, 5.003524, 
    4.967793, 4.932725, 4.899067, 4.86745, 4.838332, 4.811933, 4.788154, 
    4.766489, 4.747004, 4.743248, 4.728023, 4.715933, 4.706465, 4.699218, 
    4.698076, 4.699035, 4.70357, 4.711748, 4.723778, 4.739289, 4.757714, 
    4.777895, 4.798965, 4.818629, 4.840088, 4.857762, 4.870472, 4.877666, 
    4.879622, 4.877593, 4.873718, 4.870685, 4.871213, 4.877508, 4.890886, 
    4.911653, 4.939244, 4.972483, 5.00987, 5.049802, 5.090693, 5.131, 5.169196,
  // momentumY(12,10, 0-49)
    5.166411, 5.144372, 5.117849, 5.087887, 5.0555, 5.021643, 4.987225, 
    4.9531, 4.920068, 4.888845, 4.86002, 4.833982, 4.810833, 4.790262, 
    4.771456, 4.752806, 4.748785, 4.735146, 4.723433, 4.713244, 4.704352, 
    4.701074, 4.699321, 4.700947, 4.706553, 4.716559, 4.730864, 4.749084, 
    4.770245, 4.79319, 4.815342, 4.840149, 4.861498, 4.877731, 4.887707, 
    4.891069, 4.888515, 4.881875, 4.873897, 4.867746, 4.866354, 4.871841, 
    4.885215, 4.906405, 4.934523, 4.968196, 5.005853, 5.045899, 5.086775, 
    5.126939,
  // momentumY(12,11, 0-49)
    5.156057, 5.132392, 5.104886, 5.074547, 5.042329, 5.009131, 4.975822, 
    4.943227, 4.912133, 4.883249, 4.85715, 4.83418, 4.814344, 4.797164, 
    4.781535, 4.763055, 4.757185, 4.745727, 4.734569, 4.723561, 4.712773, 
    4.706907, 4.701915, 4.700012, 4.70236, 4.709619, 4.721997, 4.739341, 
    4.760933, 4.785336, 4.809756, 4.837816, 4.863089, 4.883525, 4.89742, 
    4.90373, 4.902445, 4.894832, 4.883407, 4.871558, 4.862848, 4.860272, 
    4.865705, 4.879758, 4.901966, 4.931159, 4.965813, 5.004309, 5.045033, 
    5.086396,
  // momentumY(12,12, 0-49)
    5.149285, 5.12441, 5.096178, 5.065566, 5.033495, 5.000843, 4.968459, 
    4.937173, 4.907782, 4.881011, 4.857444, 4.837414, 4.820879, 4.807252, 
    4.795251, 4.776213, 4.766981, 4.758471, 4.748212, 4.73646, 4.723689, 
    4.714914, 4.706287, 4.700346, 4.698822, 4.702633, 4.712355, 4.728104, 
    4.74946, 4.774756, 4.801041, 4.831972, 4.861088, 4.886032, 4.904624, 
    4.915174, 4.916892, 4.910286, 4.897347, 4.881368, 4.866335, 4.856068, 
    4.853416, 4.859857, 4.875521, 4.899554, 4.930533, 4.966812, 5.006703, 
    5.048541,
  // momentumY(12,13, 0-49)
    5.145769, 5.119963, 5.09112, 5.060205, 5.028135, 4.995795, 4.964047, 
    4.933748, 4.905724, 4.880737, 4.859405, 4.842088, 4.828754, 4.818828, 
    4.811018, 4.790828, 4.777141, 4.772433, 4.763588, 4.751352, 4.736684, 
    4.724803, 4.712266, 4.701881, 4.695943, 4.695662, 4.70202, 4.715442, 
    4.735847, 4.761384, 4.789021, 4.822229, 4.854795, 4.884152, 4.90777, 
    4.923401, 4.929517, 4.925776, 4.913407, 4.895278, 4.875484, 4.858485, 
    4.848105, 4.846823, 4.855548, 4.87389, 4.900612, 4.934071, 4.9725, 5.01414,
  // momentumY(12,14, 0-49)
    5.144871, 5.118295, 5.088853, 5.057521, 5.02524, 4.992924, 4.961475, 
    4.931789, 4.904742, 4.881144, 4.861664, 4.846729, 4.836396, 4.830227, 
    4.827164, 4.805708, 4.787249, 4.787188, 4.780379, 4.768078, 4.751752, 
    4.736667, 4.720029, 4.704872, 4.694035, 4.689069, 4.691406, 4.701812, 
    4.720558, 4.745669, 4.774117, 4.808887, 4.844282, 4.877623, 4.906136, 
    4.927167, 4.938556, 4.939137, 4.929252, 4.911079, 4.888462, 4.866208, 
    4.848984, 4.840306, 4.842016, 4.854346, 4.876366, 4.906497, 4.942909, 
    4.983748,
  // momentumY(12,15, 0-49)
    5.145796, 5.118527, 5.088447, 5.056561, 5.023852, 4.991281, 4.959796, 
    4.930346, 4.903856, 4.881192, 4.863095, 4.850088, 4.842387, 4.839818, 
    4.841783, 4.819959, 4.797536, 4.802824, 4.798692, 4.786848, 4.769209, 
    4.750873, 4.72998, 4.709755, 4.693579, 4.683396, 4.681126, 4.687901, 
    4.70434, 4.728413, 4.75718, 4.792764, 4.83025, 4.866904, 4.899821, 
    4.926082, 4.943048, 4.948842, 4.942933, 4.92663, 4.903234, 4.877543, 
    4.854808, 4.839509, 4.834488, 4.840753, 4.857808, 4.884229, 4.918171, 
    4.957691,
  // momentumY(12,16, 0-49)
    5.14775, 5.119838, 5.089086, 5.056542, 5.023234, 4.99017, 4.958349, 
    4.928762, 4.902383, 4.88013, 4.862822, 4.851107, 4.845402, 4.84588, 
    4.852536, 4.832886, 4.808788, 4.819836, 4.818934, 4.808081, 4.789505, 
    4.767872, 4.742556, 4.716972, 4.695046, 4.67918, 4.671813, 4.674458, 
    4.688052, 4.710579, 4.739286, 4.774993, 4.813807, 4.852983, 4.889573, 
    4.920512, 4.942851, 4.954165, 4.953143, 4.940207, 4.917892, 4.890668, 
    4.864047, 4.843275, 4.83217, 4.832603, 4.844646, 4.867138, 4.898277, 
    4.936063,
  // momentumY(12,17, 0-49)
    5.150093, 5.121617, 5.090219, 5.056981, 5.022968, 4.989228, 4.956792, 
    4.926682, 4.899899, 4.877413, 4.860113, 4.84878, 4.844049, 4.846456, 
    4.856596, 4.843801, 4.822259, 4.838977, 4.841652, 4.832212, 4.813004, 
    4.787975, 4.758004, 4.726743, 4.698685, 4.676764, 4.663949, 4.662121, 
    4.672501, 4.693131, 4.72155, 4.756793, 4.796225, 4.837117, 4.876529, 
    4.911358, 4.938486, 4.955118, 4.959318, 4.950685, 4.930918, 4.903908, 
    4.875101, 4.850234, 4.833983, 4.829096, 4.836311, 4.854834, 4.882985, 
    4.918743,
  // momentumY(12,18, 0-49)
    5.152446, 5.123583, 5.091654, 5.057766, 5.023003, 4.988423, 4.955067, 
    4.923962, 4.896122, 4.872548, 4.854192, 4.841951, 4.836679, 4.839291, 
    4.851016, 4.851833, 4.839601, 4.861182, 4.867465, 4.859635, 4.839867, 
    4.81117, 4.776155, 4.738822, 4.704293, 4.676091, 4.657684, 4.651282, 
    4.65831, 4.676892, 4.704975, 4.739322, 4.778765, 4.820615, 4.861983, 
    4.8998, 4.930897, 4.952261, 4.961515, 4.957573, 4.941316, 4.915917, 
    4.886491, 4.85898, 4.838706, 4.829237, 4.832021, 4.846715, 4.871841, 
    4.905409,
  // momentumY(12,19, 0-49)
    5.154763, 5.125841, 5.093623, 5.059199, 5.023643, 4.987998, 4.95329, 
    4.920535, 4.890742, 4.864912, 4.844035, 4.829114, 4.82127, 4.821993, 
    4.833523, 4.855882, 4.862566, 4.887558, 4.897141, 4.890828, 4.870145, 
    4.837114, 4.796288, 4.752288, 4.710979, 4.67649, 4.652683, 4.64197, 
    4.645842, 4.66249, 4.690382, 4.723572, 4.762553, 4.804698, 4.847201, 
    4.887078, 4.921197, 4.946469, 4.960234, 4.960886, 4.948586, 4.925761, 
    4.897009, 4.868209, 4.845094, 4.831927, 4.83085, 4.842024, 4.864239, 
    4.895589,
  // momentumY(12,20, 0-49)
    5.154693, 5.1242, 5.09093, 5.056166, 5.021146, 4.987069, 4.955105, 
    4.926386, 4.901967, 4.88274, 4.869288, 4.861674, 4.859224, 4.860402, 
    4.862944, 0, 4.887241, 4.889175, 4.884861, 4.87331, 4.854144, 4.824542, 
    4.78899, 4.749675, 4.711314, 4.677715, 4.653001, 4.640221, 4.641569, 
    4.655976, 4.682993, 4.71405, 4.751464, 4.792706, 4.835068, 4.875674, 
    4.911485, 4.939419, 4.956679, 4.961297, 4.952844, 4.933036, 4.905849, 
    4.876883, 4.852042, 4.836103, 4.831837, 4.839926, 4.859478, 4.888717,
  // momentumY(12,21, 0-49)
    5.155864, 5.125593, 5.092457, 5.057732, 5.02263, 4.988307, 4.955864, 
    4.926349, 4.90071, 4.879722, 4.863865, 4.853156, 4.846985, 4.843976, 
    4.841977, 0, 4.928431, 4.928067, 4.921334, 4.906662, 4.883474, 4.84574, 
    4.802858, 4.756638, 4.712227, 4.67375, 4.64543, 4.630235, 4.630127, 
    4.64397, 4.671875, 4.702372, 4.7396, 4.78107, 4.82414, 4.866025, 
    4.903787, 4.934397, 4.954999, 4.963388, 4.958678, 4.941965, 4.916625, 
    4.887901, 4.861739, 4.843331, 4.83602, 4.841007, 4.857741, 4.884601,
  // momentumY(12,22, 0-49)
    5.156168, 5.126009, 5.092949, 5.05825, 5.023098, 4.988604, 4.955816, 
    4.925714, 4.899168, 4.876884, 4.859283, 4.846379, 4.837635, 4.831826, 
    4.826962, 0, 4.95737, 4.955109, 4.947015, 4.931, 4.906226, 4.863213, 
    4.81588, 4.765259, 4.716686, 4.674536, 4.643195, 4.62569, 4.623909, 
    4.63674, 4.664946, 4.694184, 4.7305, 4.771442, 4.814431, 4.856776, 
    4.895633, 4.928053, 4.951179, 4.962662, 4.96128, 4.947614, 4.924472, 
    4.896675, 4.870069, 4.850082, 4.840516, 4.843034, 4.857418, 4.882221,
  // momentumY(12,23, 0-49)
    5.155862, 5.125789, 5.092804, 5.058161, 5.023019, 4.988459, 4.955489, 
    4.925042, 4.897942, 4.874845, 4.856148, 4.84187, 4.831531, 4.824033, 
    4.817537, 0, 4.976377, 4.972693, 4.963794, 4.947212, 4.921901, 4.875348, 
    4.825215, 4.771749, 4.720391, 4.675718, 4.642266, 4.623123, 4.620123, 
    4.632184, 4.660638, 4.688662, 4.724012, 4.764284, 4.806946, 4.849384, 
    4.888843, 4.92245, 4.947373, 4.961187, 4.962439, 4.951327, 4.930201, 
    4.903494, 4.876895, 4.855958, 4.8448, 4.845447, 4.857971, 4.881085,
  // momentumY(12,24, 0-49)
    5.155117, 5.125144, 5.092268, 5.057733, 5.022682, 4.988179, 4.955212, 
    4.924688, 4.897405, 4.873996, 4.85484, 4.839958, 4.828905, 4.820646, 
    4.81344, 0, 4.985891, 4.981441, 4.972165, 4.95543, 4.930089, 4.881607, 
    4.830071, 4.775189, 4.722447, 4.676545, 4.642097, 4.622215, 4.618693, 
    4.630451, 4.65923, 4.686486, 4.721179, 4.760937, 4.803261, 4.84558, 
    4.885197, 4.919293, 4.945075, 4.960088, 4.962771, 4.953119, 4.93321, 
    4.907235, 4.880754, 4.85936, 4.84734, 4.846935, 4.858387, 4.880515,
  // momentumY(12,25, 0-49)
    5.154003, 5.124162, 5.091442, 5.057076, 5.022206, 4.987893, 4.955125, 
    4.924804, 4.897723, 4.874507, 4.855525, 4.840787, 4.829843, 4.821658, 
    4.814504, 0, 4.985445, 4.981015, 4.971813, 4.955236, 4.930161, 4.881445, 
    4.829905, 4.775073, 4.722418, 4.676649, 4.642362, 4.622644, 4.61925, 
    4.63111, 4.66012, 4.687131, 4.721565, 4.761066, 4.803155, 4.84528, 
    4.884767, 4.918823, 4.94467, 4.959867, 4.962834, 4.953512, 4.933909, 
    4.908139, 4.88171, 4.860214, 4.847972, 4.847279, 4.858426, 4.880264,
  // momentumY(12,26, 0-49)
    5.152479, 5.122794, 5.090271, 5.056139, 5.021544, 4.98756, 4.955191, 
    4.925356, 4.898864, 4.876347, 4.858164, 4.84431, 4.834285, 4.826993, 
    4.820641, 0, 4.975043, 4.971416, 4.962752, 4.946657, 4.92212, 4.874942, 
    4.824836, 4.771557, 4.72049, 4.676219, 4.64323, 4.624537, 4.621883, 
    4.634203, 4.663285, 4.690606, 4.725205, 4.764738, 4.80672, 4.848597, 
    4.887678, 4.921165, 4.946287, 4.960632, 4.962692, 4.952519, 4.932245, 
    4.906088, 4.879598, 4.858325, 4.846496, 4.846295, 4.857932, 4.880213,
  // momentumY(12,27, 0-49)
    5.150397, 5.120863, 5.088561, 5.054716, 5.020484, 4.986965, 4.955193, 
    4.926123, 4.900596, 4.879271, 4.862515, 4.85029, 4.842027, 4.836516, 
    4.831839, 0, 4.955084, 4.952917, 4.945256, 4.930057, 4.906505, 4.862667, 
    4.815493, 4.76527, 4.717227, 4.67572, 4.645051, 4.628139, 4.626747, 
    4.639816, 4.668792, 4.696878, 4.731983, 4.77176, 4.813708, 4.855239, 
    4.893616, 4.925999, 4.949613, 4.96211, 4.962144, 4.950032, 4.928223, 
    4.901196, 4.874612, 4.853933, 4.843158, 4.844211, 4.857095, 4.880501,
  // momentumY(12,28, 0-49)
    5.147523, 5.118073, 5.085974, 5.052443, 5.018648, 4.985715, 4.954721, 
    4.926675, 4.902474, 4.882824, 4.868122, 4.858309, 4.85273, 4.850033, 
    4.848179, 0, 4.926608, 4.926298, 4.920071, 4.906347, 4.884541, 4.845834, 
    4.803155, 4.757463, 4.713751, 4.676086, 4.648576, 4.634062, 4.63437, 
    4.648452, 4.677229, 4.706404, 4.742229, 4.782332, 4.82418, 4.865112, 
    4.902321, 4.932904, 4.95409, 4.963649, 4.960521, 4.945456, 4.921401, 
    4.893226, 4.866715, 4.847156, 4.838172, 4.84128, 4.85618, 4.881395,
  // momentumY(12,29, 0-49)
    5.143562, 5.11403, 5.082041, 5.048799, 5.015478, 4.983227, 4.953168, 
    4.926374, 4.903827, 4.886317, 4.874309, 4.867758, 4.86593, 4.867328, 
    4.869853, 0, 4.889934, 4.891613, 4.88732, 4.875996, 4.857266, 4.825638, 
    4.789297, 4.749714, 4.711526, 4.678509, 4.654641, 4.642774, 4.644877, 
    4.659924, 4.688231, 4.718379, 4.754757, 4.794957, 4.836395, 4.876332, 
    4.911868, 4.940042, 4.958111, 4.964036, 4.957141, 4.938742, 4.912372, 
    4.883308, 4.857393, 4.839608, 4.833077, 4.838827, 4.856208, 4.883573,
  // momentumY(12,30, 0-49)
    5.140514, 5.112536, 5.081708, 5.049011, 5.015432, 4.981946, 4.949521, 
    4.919111, 4.891653, 4.868042, 4.849143, 4.835805, 4.82899, 4.830027, 
    4.841019, 4.861464, 4.864655, 4.888956, 4.899061, 4.894265, 4.875897, 
    4.843383, 4.804152, 4.761779, 4.721758, 4.68805, 4.664435, 4.653369, 
    4.656442, 4.672151, 4.699848, 4.730855, 4.767568, 4.807538, 4.848127, 
    4.886528, 4.91977, 4.944874, 4.959198, 4.960996, 4.950107, 4.928501, 
    4.900321, 4.871173, 4.846792, 4.831698, 4.828403, 4.837403, 4.857709, 
    4.887527,
  // momentumY(12,31, 0-49)
    5.134956, 5.106979, 5.076535, 5.044599, 5.012144, 4.980138, 4.949538, 
    4.921287, 4.896299, 4.875444, 4.859525, 4.84926, 4.845331, 4.848502, 
    4.859925, 4.859009, 4.845135, 4.865917, 4.872577, 4.866015, 4.848228, 
    4.820029, 4.786397, 4.750472, 4.717049, 4.68944, 4.671017, 4.664021, 
    4.67, 4.687367, 4.714871, 4.746837, 4.783939, 4.823677, 4.863338, 
    4.900009, 4.93064, 4.952261, 4.962398, 4.959703, 4.944641, 4.919906, 
    4.890231, 4.861438, 4.83902, 4.826921, 4.826994, 4.839206, 4.862264, 
    4.894248,
  // momentumY(12,32, 0-49)
    5.129212, 5.101433, 5.071481, 5.040294, 5.008811, 4.97796, 4.948673, 
    4.921868, 4.898431, 4.87919, 4.864866, 4.856045, 4.853179, 4.856658, 
    4.867016, 4.852871, 4.831022, 4.847097, 4.850173, 4.841893, 4.824452, 
    4.79999, 4.771226, 4.741108, 4.713883, 4.692271, 4.679163, 4.676469, 
    4.685562, 4.704714, 4.732142, 4.764843, 4.801892, 4.840762, 4.878683, 
    4.912685, 4.939712, 4.956912, 4.96214, 4.954616, 4.93555, 4.908378, 
    4.878297, 4.851113, 4.831837, 4.823677, 4.827783, 4.84363, 4.869668, 
    4.90391,
  // momentumY(12,33, 0-49)
    5.12343, 5.095872, 5.066374, 5.035829, 5.005118, 4.975122, 4.946723, 
    4.920801, 4.898202, 4.879708, 4.865957, 4.8574, 4.854257, 4.856545, 
    4.864198, 4.843874, 4.820434, 4.831309, 4.831038, 4.821383, 4.804472, 
    4.783561, 4.75934, 4.73466, 4.713286, 4.697415, 4.689446, 4.690929, 
    4.70299, 4.723768, 4.751048, 4.784074, 4.82048, 4.857722, 4.89301, 
    4.92337, 4.945841, 4.957834, 4.957703, 4.945395, 4.922944, 4.894461, 
    4.865391, 4.841245, 4.82632, 4.822978, 4.831672, 4.851446, 4.880571, 
    4.91704,
  // momentumY(12,34, 0-49)
    5.118104, 5.090694, 5.0615, 5.031375, 5.001149, 4.971647, 4.943697, 
    4.918133, 4.895763, 4.877318, 4.863366, 4.854235, 4.849931, 4.850104, 
    4.854072, 4.83257, 4.811661, 4.817543, 4.81448, 4.804032, 4.788081, 
    4.770701, 4.75087, 4.731368, 4.715502, 4.705021, 4.701844, 4.707161, 
    4.721816, 4.74386, 4.770767, 4.803555, 4.838606, 4.873378, 4.905098, 
    4.930877, 4.947974, 4.954234, 4.948682, 4.932118, 4.907397, 4.87913, 
    4.852721, 4.83309, 4.823634, 4.825835, 4.8395, 4.863335, 4.895511, 
    4.934046,
  // momentumY(12,35, 0-49)
    5.113986, 5.086621, 5.057515, 5.027502, 4.997377, 4.967923, 4.939924, 
    4.914174, 4.891447, 4.872436, 4.85766, 4.847354, 4.841359, 4.839027, 
    4.839162, 4.81933, 4.803371, 4.80494, 4.799863, 4.789345, 4.774886, 
    4.761084, 4.745565, 4.731028, 4.720322, 4.714813, 4.715966, 4.724633, 
    4.74135, 4.764152, 4.790324, 4.822191, 4.855091, 4.886513, 4.913769, 
    4.934159, 4.945316, 4.945704, 4.935174, 4.915422, 4.890007, 4.863766, 
    4.841733, 4.827977, 4.824899, 4.833127, 4.851935, 4.879796, 4.914845, 
    4.955168,
  // momentumY(12,36, 0-49)
    5.111942, 5.084561, 5.055326, 5.025081, 4.994619, 4.964703, 4.936105, 
    4.909595, 4.885931, 4.865786, 4.849653, 4.83772, 4.829732, 4.824864, 
    4.821609, 4.804615, 4.794687, 4.792881, 4.786672, 4.776821, 4.764374, 
    4.754197, 4.742932, 4.733154, 4.727239, 4.726232, 4.731174, 4.742603, 
    4.760743, 4.7837, 4.808667, 4.838854, 4.868789, 4.896034, 4.918074, 
    4.932533, 4.937595, 4.932491, 4.91799, 4.896621, 4.872406, 4.850078, 
    4.833977, 4.827167, 4.831044, 4.845499, 4.8694, 4.901079, 4.938695, 
    4.980416,
  // momentumY(12,37, 0-49)
    5.112801, 5.08544, 5.055923, 5.025138, 4.993912, 4.963036, 4.933292, 
    4.905466, 4.880316, 4.858521, 4.840577, 4.826664, 4.81651, 4.809246, 
    4.803285, 4.789212, 4.785302, 4.781154, 4.774646, 4.766088, 4.756061, 
    4.7495, 4.742392, 4.737138, 4.735608, 4.738574, 4.746701, 4.76024, 
    4.779102, 4.801551, 4.82479, 4.852537, 4.878767, 4.901183, 4.917546, 
    4.92596, 4.9253, 4.915676, 4.898742, 4.877671, 4.856634, 4.839904, 
    4.830922, 4.831695, 4.84272, 4.863298, 4.892019, 4.927155, 4.966915, 
    5.009552,
  // momentumY(12,38, 0-49)
    5.117163, 5.089993, 5.060169, 5.028653, 4.996345, 4.964101, 4.932761, 
    4.903154, 4.876072, 4.852218, 4.83211, 4.815961, 4.803544, 4.794055, 
    4.786015, 4.774364, 4.77559, 4.770068, 4.763923, 4.757067, 4.749672, 
    4.746599, 4.743455, 4.742412, 4.744793, 4.75115, 4.761802, 4.776754, 
    4.795622, 4.81691, 4.837911, 4.862556, 4.884535, 4.90178, 4.912446, 
    4.915242, 4.909836, 4.897208, 4.879747, 4.860974, 4.844863, 4.834976, 
    4.833762, 4.842255, 4.86022, 4.886531, 4.919603, 4.957696, 4.999078, 
    5.042069,
  // momentumY(12,39, 0-49)
    5.125264, 5.098615, 5.068628, 5.036368, 5.002841, 4.969013, 4.935816, 
    4.904154, 4.874874, 4.84872, 4.826249, 4.807725, 4.793006, 4.781432, 
    4.771742, 4.761746, 4.766644, 4.760505, 4.755105, 4.750071, 4.74527, 
    4.745384, 4.745862, 4.74859, 4.754327, 4.763429, 4.775914, 4.791576, 
    4.809772, 4.829317, 4.847673, 4.868758, 4.88626, 4.898421, 4.903902, 
    4.902092, 4.893451, 4.879701, 4.863706, 4.849003, 4.839085, 4.836678, 
    4.843287, 4.859147, 4.883482, 4.914883, 4.951668, 4.992102, 5.034494, 
    5.077206,
  // momentumY(12,40, 0-49)
    5.136877, 5.111238, 5.081432, 5.048639, 5.014005, 4.978633, 4.943581, 
    4.909848, 4.878351, 4.849883, 4.825041, 4.804149, 4.787166, 4.773599, 
    4.76246, 4.753274, 4.760116, 4.753808, 4.749212, 4.745819, 4.743309, 
    4.746111, 4.749687, 4.755607, 4.764044, 4.775191, 4.788807, 4.804513, 
    4.821455, 4.83882, 4.854307, 4.871682, 4.884876, 4.892533, 4.893868, 
    4.888951, 4.878927, 4.866021, 4.853262, 4.843918, 4.840827, 4.845891, 
    4.859829, 4.882285, 4.912125, 4.94777, 4.987484, 5.029533, 5.072239, 
    5.113965,
  // momentumY(12,41, 0-49)
    5.151308, 5.127309, 5.098226, 5.065358, 5.030005, 4.993429, 4.956825, 
    4.921301, 4.887843, 4.857288, 4.830274, 4.807172, 4.78804, 4.772555, 
    4.759991, 4.750806, 4.757907, 4.751545, 4.747518, 4.745323, 4.744565, 
    4.749381, 4.755365, 4.763759, 4.774164, 4.786629, 4.800695, 4.81586, 
    4.83112, 4.846073, 4.858711, 4.872571, 4.882043, 4.886209, 4.884839, 
    4.878588, 4.869079, 4.858769, 4.850559, 4.847245, 4.850982, 4.862956, 
    4.883301, 4.911276, 4.945533, 4.98441, 5.026139, 5.068966, 5.111191, 
    5.151146,
  // momentumY(12,42, 0-49)
    5.167433, 5.145825, 5.118198, 5.085958, 5.05056, 5.013422, 4.975871, 
    4.939118, 4.904213, 4.872023, 4.84321, 4.818187, 4.797098, 4.779766, 
    4.765706, 4.755823, 4.761775, 4.755195, 4.751298, 4.749695, 4.749995, 
    4.756035, 4.763631, 4.773695, 4.7853, 4.798368, 4.81227, 4.826428, 
    4.839757, 4.852291, 4.862344, 4.873213, 4.879873, 4.881848, 4.879389, 
    4.873567, 4.866244, 4.859843, 4.856923, 4.859726, 4.86978, 4.887712, 
    4.91327, 4.945491, 4.982934, 5.023899, 5.066599, 5.109246, 5.150087, 
    5.187401,
  // momentumY(12,43, 0-49)
    5.183809, 5.165433, 5.140165, 5.109489, 5.074985, 5.038198, 5.000572, 
    4.963393, 4.927755, 4.894545, 4.864434, 4.837869, 4.815063, 4.795979, 
    4.780333, 4.769211, 4.773004, 4.765872, 4.76158, 4.759906, 4.760523, 
    4.766987, 4.77537, 4.786294, 4.798351, 4.811367, 4.824594, 4.837421, 
    4.848752, 4.859057, 4.866989, 4.875616, 4.880549, 4.881706, 4.879692, 
    4.875801, 4.871909, 4.870196, 4.872773, 4.881325, 4.896852, 4.919589, 
    4.94904, 4.984147, 5.023449, 5.065253, 5.107759, 5.149135, 5.187568, 
    5.22127,
  // momentumY(12,44, 0-49)
    5.198803, 5.184547, 5.162685, 5.134711, 5.102264, 5.066974, 5.03035, 
    4.993721, 4.9582, 4.924677, 4.893834, 4.866149, 4.841905, 4.821187, 
    4.803893, 4.791168, 4.792223, 4.784158, 4.778965, 4.776611, 4.77686, 
    4.783025, 4.79144, 4.802482, 4.814332, 4.826746, 4.838907, 4.85022, 
    4.859634, 4.868042, 4.874416, 4.881635, 4.88592, 4.887495, 4.887174, 
    4.886299, 4.886583, 4.889843, 4.897708, 4.911355, 4.931366, 4.957692, 
    4.989709, 5.026331, 5.066129, 5.10744, 5.148468, 5.187353, 5.222224, 
    5.251262,
  // momentumY(12,45, 0-49)
    5.210752, 5.201502, 5.184183, 5.160196, 5.131147, 5.098663, 5.064255, 
    5.029252, 4.994759, 4.961669, 4.930681, 4.902313, 4.876929, 4.854733, 
    4.835791, 4.821271, 4.819385, 4.810057, 4.803559, 4.800041, 4.799366, 
    4.804659, 4.81249, 4.82304, 4.834153, 4.845552, 4.856387, 4.866125, 
    4.873801, 4.880695, 4.886077, 4.892675, 4.897229, 4.900172, 4.9024, 
    4.905163, 4.909904, 4.918032, 4.9307, 4.948648, 4.972125, 5.000875, 
    5.034193, 5.071006, 5.109934, 5.149368, 5.187541, 5.222595, 5.252655, 
    5.275915,
  // momentumY(12,46, 0-49)
    5.218122, 5.214686, 5.20306, 5.184418, 5.160201, 5.131918, 5.101005, 
    5.068739, 5.036206, 5.004301, 4.973755, 4.945153, 4.91895, 4.895483, 
    4.874975, 4.858628, 4.853901, 4.843082, 4.835012, 4.830008, 4.828019, 
    4.832044, 4.838839, 4.848449, 4.858446, 4.868553, 4.87793, 4.886125, 
    4.892288, 4.898044, 4.902914, 4.909524, 4.915015, 4.919935, 4.925162, 
    4.93177, 4.940877, 4.953484, 4.970314, 4.991725, 5.017685, 5.047775, 
    5.081226, 5.116975, 5.153697, 5.189855, 5.223742, 5.253561, 5.277506, 
    5.293887,
  // momentumY(12,47, 0-49)
    5.21968, 5.222688, 5.21781, 5.205827, 5.18786, 5.16517, 5.139026, 
    5.110605, 5.080956, 5.050987, 5.021486, 4.993125, 4.966475, 4.942011, 
    4.920112, 4.902047, 4.89479, 4.88238, 4.87262, 4.865965, 4.86244, 
    4.86497, 4.870446, 4.87882, 4.88747, 4.896142, 4.904027, 4.910778, 
    4.91566, 4.9206, 4.925312, 4.932374, 4.939193, 4.946368, 4.954691, 
    4.965012, 4.978126, 4.994638, 5.014892, 5.038917, 5.066428, 5.09685, 
    5.129348, 5.162853, 5.19609, 5.227598, 5.255783, 5.278975, 5.295548, 
    5.304067,
  // momentumY(12,48, 0-49)
    5.214645, 5.224436, 5.227116, 5.222918, 5.212476, 5.196669, 5.176497, 
    5.152991, 5.127141, 5.099882, 5.07207, 5.044486, 5.017835, 4.992734, 
    4.969724, 4.950169, 4.940837, 4.926858, 4.91543, 4.907111, 4.90198, 
    4.902931, 4.906935, 4.913908, 4.921101, 4.9283, 4.934745, 4.940191, 
    4.944019, 4.94839, 4.953168, 4.960919, 4.969209, 4.978634, 4.989865, 
    5.003521, 5.020082, 5.039804, 5.062685, 5.088459, 5.11661, 5.146403, 
    5.176918, 5.207063, 5.235599, 5.261165, 5.28232, 5.297623, 5.305756, 
    5.305692,
  // momentumY(12,49, 0-49)
    5.192284, 5.210041, 5.222421, 5.228807, 5.229014, 5.22324, 5.211989, 
    5.195982, 5.176065, 5.153151, 5.128168, 5.102034, 5.075628, 5.049784, 
    5.025281, 5.004552, 5.000236, 4.983833, 4.969202, 4.957649, 4.949624, 
    4.951151, 4.956371, 4.96534, 4.972784, 4.978915, 4.982822, 4.984548, 
    4.983208, 4.98358, 4.985592, 4.994268, 5.004465, 5.016714, 5.031483, 
    5.049073, 5.069549, 5.092734, 5.118204, 5.145324, 5.173291, 5.201159, 
    5.227886, 5.252362, 5.273417, 5.289875, 5.300619, 5.304664, 5.301308, 
    5.290269,
  // momentumY(13,0, 0-49)
    5.302906, 5.297866, 5.283644, 5.261401, 5.232627, 5.198957, 5.162014, 
    5.123312, 5.084203, 5.045848, 5.009209, 4.975058, 4.943973, 4.916348, 
    4.892391, 4.872317, 4.857236, 4.844203, 4.834624, 4.828238, 4.824745, 
    4.82422, 4.826094, 4.830255, 4.836333, 4.844073, 4.853085, 4.862946, 
    4.873157, 4.88348, 4.893552, 4.903595, 4.913329, 4.923114, 4.933573, 
    4.945522, 4.959881, 4.977537, 4.999209, 5.025342, 5.056015, 5.090916, 
    5.129323, 5.170135, 5.211916, 5.252959, 5.291361, 5.325141, 5.352355, 
    5.371239,
  // momentumY(13,1, 0-49)
    5.28951, 5.280722, 5.263025, 5.237669, 5.206186, 5.170209, 5.131349, 
    5.091095, 5.05077, 5.011506, 4.974237, 4.939699, 4.908432, 4.880779, 
    4.856899, 4.837128, 4.823848, 4.810921, 4.801519, 4.795393, 4.792206, 
    4.792432, 4.795098, 4.800194, 4.807179, 4.81584, 4.825731, 4.836394, 
    4.847203, 4.858047, 4.868423, 4.878859, 4.888578, 4.897897, 4.907441, 
    4.918092, 4.930884, 4.946864, 4.966928, 4.991677, 5.021327, 5.055649, 
    5.093979, 5.135242, 5.178015, 5.220617, 5.26118, 5.297764, 5.328457, 
    5.351484,
  // momentumY(13,2, 0-49)
    5.270072, 5.257787, 5.237234, 5.209664, 5.176543, 5.139416, 5.099804, 
    5.059119, 5.018622, 4.979402, 4.942351, 4.90817, 4.877359, 4.850216, 
    4.826835, 4.807679, 4.796417, 4.78367, 4.774438, 4.768469, 4.765407, 
    4.766132, 4.769279, 4.774964, 4.782534, 4.791835, 4.802403, 4.813765, 
    4.825194, 4.836684, 4.847581, 4.858711, 4.868759, 4.877928, 4.886779, 
    4.896184, 4.907245, 4.921134, 4.938916, 4.961381, 4.988906, 5.021394, 
    5.058273, 5.098534, 5.14082, 5.18352, 5.224868, 5.263035, 5.29622, 
    5.322726,
  // momentumY(13,3, 0-49)
    5.246368, 5.230927, 5.208125, 5.179145, 5.145323, 5.108055, 5.068716, 
    5.028602, 4.988883, 4.950584, 4.914549, 4.881436, 4.851695, 4.825564, 
    4.803069, 4.78479, 4.775711, 4.763161, 4.754032, 4.748058, 4.744871, 
    4.745768, 4.749006, 4.754856, 4.762612, 4.77221, 4.783199, 4.795122, 
    4.807179, 4.819442, 4.831099, 4.843277, 4.85408, 4.863536, 4.872057, 
    4.880424, 4.889727, 4.901223, 4.916138, 4.935462, 4.959786, 4.989203, 
    5.023292, 5.061168, 5.10159, 5.143067, 5.183972, 5.222636, 5.257412, 
    5.286727,
  // momentumY(13,4, 0-49)
    5.220337, 5.202127, 5.177616, 5.147886, 5.114111, 5.077507, 5.039276, 
    5.000571, 4.962453, 4.925858, 4.89157, 4.860184, 4.83209, 4.80745, 
    4.786195, 4.768989, 4.762178, 4.749801, 4.740659, 4.734465, 4.730842, 
    4.731516, 4.734381, 4.73989, 4.747362, 4.756843, 4.767935, 4.780223, 
    4.792881, 4.806018, 4.818665, 4.832267, 4.844315, 4.854602, 4.863307, 
    4.871026, 4.878742, 4.887725, 4.899331, 4.91477, 4.934896, 4.960064, 
    4.990092, 5.024294, 5.061602, 5.100693, 5.140108, 5.178351, 5.21394, 
    5.245433,
  // momentumY(13,5, 0-49)
    5.193888, 5.173308, 5.147536, 5.117548, 5.084359, 5.048999, 5.012493, 
    4.975842, 4.939978, 4.905743, 4.873834, 4.84477, 4.818851, 4.796136, 
    4.776439, 4.760425, 4.755842, 4.743599, 4.734304, 4.72764, 4.723233, 
    4.723243, 4.725216, 4.729818, 4.736472, 4.745353, 4.756155, 4.768545, 
    4.781706, 4.795761, 4.809578, 4.824949, 4.838744, 4.850475, 4.860016, 
    4.867673, 4.874217, 4.880829, 4.88893, 4.899941, 4.915029, 4.9349, 
    4.959711, 4.989072, 5.022166, 5.057874, 5.094924, 5.131988, 5.167728, 
    5.200819,
  // momentumY(13,6, 0-49)
    5.168723, 5.146162, 5.119484, 5.089571, 5.057295, 5.023526, 4.989129, 
    4.954954, 4.92181, 4.890425, 4.861399, 4.835148, 4.811861, 4.791458, 
    4.773588, 4.758794, 4.756223, 4.744107, 4.734529, 4.727149, 4.721606, 
    4.720503, 4.721052, 4.724154, 4.729415, 4.737158, 4.74721, 4.759347, 
    4.772826, 4.78774, 4.802809, 4.820201, 4.836185, 4.849976, 4.861088, 
    4.869447, 4.875493, 4.880192, 4.884932, 4.891296, 4.900784, 4.914537, 
    4.933163, 4.956684, 4.984612, 5.016095, 5.050054, 5.085308, 5.12063, 
    5.154777,
  // momentumY(13,7, 0-49)
    5.146191, 5.122014, 5.094694, 5.065038, 5.033816, 5.001769, 4.969636, 
    4.938137, 4.907962, 4.879731, 4.853929, 4.830854, 4.810551, 4.792776, 
    4.776973, 4.763321, 4.762328, 4.750426, 4.740496, 4.732202, 4.72523, 
    4.722604, 4.721231, 4.72226, 4.725554, 4.73159, 4.740366, 4.751813, 
    4.765307, 4.780891, 4.797148, 4.816651, 4.835127, 4.851506, 4.864916, 
    4.874842, 4.881288, 4.884869, 4.886801, 4.888733, 4.892467, 4.899627, 
    4.911375, 4.928267, 4.950256, 4.976807, 5.007057, 5.039953, 5.074344, 
    5.109021,
  // momentumY(13,8, 0-49)
    5.12719, 5.101721, 5.073936, 5.044599, 5.01441, 4.984032, 4.95411, 
    4.92527, 4.898105, 4.873127, 4.850711, 4.831019, 4.81394, 4.799034, 
    4.785518, 4.77283, 4.772757, 4.761313, 4.751078, 4.74178, 4.733187, 
    4.728723, 4.725017, 4.723469, 4.724253, 4.728013, 4.734952, 4.745189, 
    4.758284, 4.7742, 4.791411, 4.812908, 4.833974, 4.853284, 4.869596, 
    4.881938, 4.889804, 4.893339, 4.893427, 4.891637, 4.889973, 4.890526, 
    4.895082, 4.90484, 4.920309, 4.941354, 4.96736, 4.997399, 5.030363, 
    5.06504,
  // momentumY(13,9, 0-49)
    5.112118, 5.085622, 5.057474, 5.028415, 4.999117, 4.970207, 4.94228, 
    4.915903, 4.891597, 4.869787, 4.850737, 4.834479, 4.820738, 4.808884, 
    4.7979, 4.785911, 4.785915, 4.775369, 4.765037, 4.754792, 4.744537, 
    4.73805, 4.731728, 4.727205, 4.725008, 4.725948, 4.730473, 4.738923, 
    4.7511, 4.766879, 4.784646, 4.8078, 4.831308, 4.853636, 4.873232, 
    4.888683, 4.898961, 4.903659, 4.903191, 4.898856, 4.892699, 4.88718, 
    4.884699, 4.887177, 4.895783, 4.910887, 4.932183, 4.958889, 4.989927, 
    5.024058,
  // momentumY(13,10, 0-49)
    5.100892, 5.073568, 5.045088, 5.016195, 4.987566, 4.959826, 4.933566, 
    4.909325, 4.887583, 4.868696, 4.852839, 4.839923, 4.829534, 4.820874, 
    4.812728, 4.801129, 4.800285, 4.791276, 4.781237, 4.770275, 4.758482, 
    4.749933, 4.740851, 4.733079, 4.727515, 4.725141, 4.726683, 4.732738, 
    4.743409, 4.758473, 4.776271, 4.800553, 4.826117, 4.851284, 4.874251, 
    4.893243, 4.906741, 4.913769, 4.914171, 4.908805, 4.899549, 4.88904, 
    4.880201, 4.875673, 4.877369, 4.886271, 4.902476, 4.925397, 4.954008, 
    4.987036,
  // momentumY(13,11, 0-49)
    5.093023, 5.064999, 5.036164, 5.007285, 4.979065, 4.952162, 4.927186, 
    4.904684, 4.885119, 4.868808, 4.855855, 4.846086, 4.838981, 4.833637, 
    4.828726, 4.817231, 4.814683, 4.807994, 4.798809, 4.787527, 4.774482, 
    4.76396, 4.75211, 4.74093, 4.731703, 4.725581, 4.723604, 4.726661, 
    4.7352, 4.748919, 4.766147, 4.790886, 4.817931, 4.845511, 4.87165, 
    4.894293, 4.911518, 4.921821, 4.924446, 4.919686, 4.909037, 4.895079, 
    4.881061, 4.870255, 4.86534, 4.868004, 4.878853, 4.897589, 4.923282, 
    4.954648,
  // momentumY(13,12, 0-49)
    5.087749, 5.05909, 5.029847, 5.00082, 4.972756, 4.946362, 4.92229, 
    4.901118, 4.883312, 4.869174, 4.858771, 4.851879, 4.847934, 4.846014, 
    4.844818, 4.833281, 4.828422, 4.824882, 4.817225, 4.80616, 4.792282, 
    4.779981, 4.765455, 4.75081, 4.737704, 4.727466, 4.721484, 4.720968, 
    4.72675, 4.738482, 4.754528, 4.778989, 4.806825, 4.836215, 4.865081, 
    4.891179, 4.912287, 4.926467, 4.932404, 4.92977, 4.919513, 4.903913, 
    4.886283, 4.870348, 4.859491, 4.856153, 4.861555, 4.875796, 4.898129, 
    4.927302,
  // momentumY(13,13, 0-49)
    5.084192, 5.054919, 5.025204, 4.995886, 4.967764, 4.941601, 4.918097, 
    4.897873, 4.881418, 4.86904, 4.860798, 4.856464, 4.8555, 4.857069, 
    4.860056, 4.848661, 4.84133, 4.84169, 4.836272, 4.826051, 4.811856, 
    4.798031, 4.780994, 4.762904, 4.745772, 4.731121, 4.720706, 4.716094, 
    4.718533, 4.727675, 4.741975, 4.765423, 4.793318, 4.823824, 4.854806, 
    4.883918, 4.908742, 4.927023, 4.936974, 4.937667, 4.929421, 4.914011, 
    4.894545, 4.874947, 4.859157, 4.850342, 4.850424, 4.860008, 4.878631, 
    4.905142,
  // momentumY(13,14, 0-49)
    5.081517, 5.05163, 5.021392, 4.991681, 4.963344, 4.937195, 4.913986, 
    4.89438, 4.878895, 4.867865, 4.861372, 4.85923, 4.860987, 4.865987, 
    4.87346, 4.863003, 4.853669, 4.858477, 4.855946, 4.847213, 4.833271, 
    4.818205, 4.798866, 4.777408, 4.756172, 4.736881, 4.721683, 4.712525, 
    4.7111, 4.717124, 4.729209, 4.750969, 4.778223, 4.809133, 4.841548, 
    4.873077, 4.901201, 4.923458, 4.937708, 4.942506, 4.937534, 4.923936, 
    4.904391, 4.882751, 4.863289, 4.849806, 4.844934, 4.849881, 4.864576, 
    4.888054,
  // momentumY(13,15, 0-49)
    5.079049, 5.048556, 5.017774, 4.987615, 4.958967, 4.932677, 4.909543, 
    4.890262, 4.875388, 4.865291, 4.8601, 4.859703, 4.863788, 4.871943, 
    4.883821, 4.876032, 4.865983, 4.875477, 4.876322, 4.869667, 4.856545, 
    4.840522, 4.819111, 4.794412, 4.769051, 4.744977, 4.724737, 4.710681, 
    4.704965, 4.707441, 4.716984, 4.73648, 4.762472, 4.793127, 4.826293, 
    4.859575, 4.890423, 4.916268, 4.934734, 4.94397, 4.943079, 4.932546, 
    4.914461, 4.892363, 4.870615, 4.853478, 4.844249, 4.844784, 4.855497, 
    4.875701,
  // momentumY(13,16, 0-49)
    5.076357, 5.04529, 5.013985, 4.983371, 4.954356, 4.927814, 4.90456, 
    4.885322, 4.870687, 4.861065, 4.85665, 4.857431, 4.863256, 4.873969, 
    4.889624, 4.887436, 4.878976, 4.892997, 4.897475, 4.893355, 4.881554, 
    4.864819, 4.841561, 4.813771, 4.784333, 4.755423, 4.729992, 4.710805, 
    4.700493, 4.699131, 4.705956, 4.722753, 4.746984, 4.776818, 4.810111, 
    4.844488, 4.877415, 4.906292, 4.928608, 4.942223, 4.945766, 4.939097, 
    4.923651, 4.902481, 4.879802, 4.860133, 4.84732, 4.843862, 4.850718, 
    4.867552,
  // momentumY(13,17, 0-49)
    5.073276, 5.041718, 5.00995, 4.978906, 4.949494, 4.922585, 4.899002, 
    4.879483, 4.864644, 4.854941, 4.850645, 4.851858, 4.858593, 4.870928, 
    4.889231, 4.896774, 4.893412, 4.911368, 4.919476, 4.918165, 4.908042, 
    4.890761, 4.865815, 4.835064, 4.801618, 4.767901, 4.737255, 4.712861, 
    4.697815, 4.692492, 4.696613, 4.710435, 4.732548, 4.761121, 4.794013, 
    4.828882, 4.86324, 4.894509, 4.920127, 4.937771, 4.94571, 4.943258, 
    4.931211, 4.912036, 4.889621, 4.86853, 4.853006, 4.846128, 4.849413, 
    4.862942,
  // momentumY(13,18, 0-49)
    5.069894, 5.037993, 5.005871, 4.974439, 4.94458, 4.917144, 4.89294, 
    4.872707, 4.857082, 4.846572, 4.841537, 4.842215, 4.848804, 4.861626, 
    4.881323, 4.903514, 4.910012, 4.930978, 4.94249, 4.944072, 4.935783, 
    4.917948, 4.891298, 4.857579, 4.820136, 4.781682, 4.745924, 4.716439, 
    4.696753, 4.687572, 4.689219, 4.699979, 4.719781, 4.746784, 4.778859, 
    4.813701, 4.848888, 4.881894, 4.910168, 4.931293, 4.943286, 4.945026, 
    4.936729, 4.920257, 4.899048, 4.877536, 4.860189, 4.850558, 4.850698, 
    4.861127,
  // momentumY(13,19, 0-49)
    5.066533, 5.034526, 5.002198, 4.970406, 4.939985, 4.911748, 4.886477, 
    4.864903, 4.847689, 4.835394, 4.828495, 4.827422, 4.832679, 4.845, 
    4.865422, 4.907155, 4.92915, 4.952248, 4.966908, 4.971374, 4.964861, 
    4.946195, 4.917465, 4.88041, 4.838736, 4.795547, 4.754904, 4.720706, 
    4.696789, 4.684154, 4.683802, 4.691631, 4.709097, 4.734366, 4.765323, 
    4.799715, 4.83519, 4.869302, 4.899551, 4.923498, 4.939002, 4.944619, 
    4.940077, 4.926665, 4.907319, 4.886206, 4.86786, 4.856178, 4.853689, 
    4.861349,
  // momentumY(13,20, 0-49)
    5.062326, 5.029428, 4.996673, 4.965066, 4.935573, 4.909109, 4.88653, 
    4.868585, 4.85582, 4.848474, 4.846332, 4.848631, 4.854045, 4.860835, 
    4.867209, 0, 4.960554, 4.96489, 4.966611, 4.9642, 4.956264, 4.938369, 
    4.913416, 4.881072, 4.843659, 4.803276, 4.763498, 4.72832, 4.70213, 
    4.68676, 4.684481, 4.689006, 4.70359, 4.72649, 4.755638, 4.788839, 
    4.823808, 4.858182, 4.88953, 4.915427, 4.93366, 4.942553, 4.941444, 
    4.931111, 4.913975, 4.893856, 4.875212, 4.86215, 4.857589, 4.862891,
  // momentumY(13,21, 0-49)
    5.05939, 5.026729, 4.99416, 4.962648, 4.9331, 4.906367, 4.883225, 
    4.864333, 4.850152, 4.840854, 4.836205, 4.83551, 4.837572, 4.840788, 
    4.843318, 0, 4.988412, 4.991874, 4.992982, 4.989769, 4.980573, 4.958037, 
    4.92908, 4.892868, 4.851937, 4.808477, 4.766072, 4.728681, 4.700647, 
    4.683903, 4.681386, 4.684261, 4.697501, 4.719358, 4.747776, 4.780595, 
    4.815596, 4.850495, 4.882943, 4.910565, 4.93112, 4.942796, 4.944633, 
    4.936992, 4.921839, 4.902638, 4.883723, 4.869337, 4.862715, 4.865593,
  // momentumY(13,22, 0-49)
    5.056715, 5.024198, 4.991746, 4.960288, 4.930684, 4.903732, 4.880151, 
    4.860536, 4.845291, 4.834549, 4.828082, 4.825235, 4.824912, 4.825584, 
    4.825378, 0, 5.007531, 5.01016, 5.010991, 5.007695, 4.998391, 4.972798, 
    4.941637, 4.903322, 4.860387, 4.814988, 4.770687, 4.731456, 4.701693, 
    4.683507, 4.680566, 4.681566, 4.693231, 4.713815, 4.741263, 4.773442, 
    4.808179, 4.843255, 4.876388, 4.905256, 4.92762, 4.941576, 4.94595, 
    4.940767, 4.927596, 4.90955, 4.890788, 4.875599, 4.867455, 4.868394,
  // momentumY(13,23, 0-49)
    5.054629, 5.022224, 4.989868, 4.958463, 4.928839, 4.901758, 4.877898, 
    4.857814, 4.841877, 4.830197, 4.822548, 4.818313, 4.816451, 4.815497, 
    4.813565, 0, 5.020011, 5.021922, 5.022535, 5.019291, 5.010156, 4.982364, 
    4.949795, 4.910171, 4.86599, 4.819386, 4.773896, 4.733502, 4.702621, 
    4.683495, 4.680393, 4.679896, 4.690282, 4.709814, 4.73644, 4.768047, 
    4.802501, 4.837631, 4.871211, 4.900962, 4.924655, 4.940331, 4.946666, 
    4.94344, 4.931912, 4.914906, 4.89641, 4.880715, 4.871446, 4.870869,
  // momentumY(13,24, 0-49)
    5.053342, 5.021052, 4.988799, 4.957475, 4.927895, 4.900801, 4.876853, 
    4.856582, 4.840339, 4.828224, 4.820012, 4.8151, 4.812484, 4.810732, 
    4.807968, 0, 5.026357, 5.027834, 5.028316, 5.025136, 5.016194, 4.987086, 
    4.953739, 4.913423, 4.868618, 4.821458, 4.775474, 4.734633, 4.703346, 
    4.683897, 4.680958, 4.67964, 4.689296, 4.708194, 4.734291, 4.765488, 
    4.799673, 4.834713, 4.868412, 4.898533, 4.92286, 4.939422, 4.946823, 
    4.944707, 4.934157, 4.91782, 4.899562, 4.883654, 4.873792, 4.872372,
  // momentumY(13,25, 0-49)
    5.052937, 5.020776, 4.988652, 4.957452, 4.927993, 4.901019, 4.877185, 
    4.857019, 4.840869, 4.828824, 4.820656, 4.815761, 4.813137, 4.811367, 
    4.80859, 0, 5.026131, 5.027595, 5.028104, 5.025001, 5.016189, 4.986772, 
    4.953303, 4.912925, 4.868127, 4.821061, 4.775249, 4.73463, 4.703572, 
    4.684343, 4.681725, 4.680303, 4.68982, 4.708557, 4.734481, 4.76551, 
    4.799545, 4.834464, 4.868091, 4.898201, 4.922594, 4.939297, 4.946908, 
    4.945036, 4.934718, 4.918549, 4.900354, 4.884392, 4.874371, 4.872713,
  // momentumY(13,26, 0-49)
    5.053365, 5.021352, 4.989378, 4.958348, 4.92909, 4.902367, 4.878851, 
    4.859085, 4.843421, 4.831948, 4.824425, 4.82023, 4.81834, 4.817324, 
    4.815344, 0, 5.019228, 5.021117, 5.02184, 5.018843, 5.010098, 4.981457, 
    4.948575, 4.908823, 4.864714, 4.818419, 4.773448, 4.7337, 4.703471, 
    4.684952, 4.682744, 4.681938, 4.691911, 4.710961, 4.737072, 4.768174, 
    4.802174, 4.836944, 4.870301, 4.900016, 4.923895, 4.939982, 4.946925, 
    4.944401, 4.933534, 4.917, 4.89867, 4.8828, 4.873055, 4.871789,
  // momentumY(13,27, 0-49)
    5.054453, 5.022583, 4.990769, 4.959939, 4.930949, 4.904599, 4.881593, 
    4.862506, 4.847711, 4.837303, 4.831028, 4.82823, 4.827834, 4.828379, 
    4.828067, 0, 5.005809, 5.008458, 5.00954, 5.006703, 4.998044, 4.971261, 
    4.939735, 4.901355, 4.858659, 4.813832, 4.770372, 4.732119, 4.703287, 
    4.685929, 4.684206, 4.684655, 4.695604, 4.715379, 4.741986, 4.773363, 
    4.807406, 4.841971, 4.874848, 4.903781, 4.926571, 4.941309, 4.946741, 
    4.942723, 4.93059, 4.913219, 4.894607, 4.879008, 4.86998, 4.869713,
  // momentumY(13,28, 0-49)
    5.055897, 5.024127, 4.992451, 4.961824, 4.933147, 4.907266, 4.884938, 
    4.866787, 4.853227, 4.844376, 4.839968, 4.839299, 4.841219, 4.844214, 
    4.846556, 0, 4.986444, 4.989986, 4.991482, 4.988878, 4.980467, 4.956567, 
    4.927253, 4.891089, 4.850602, 4.80798, 4.766706, 4.730566, 4.703684, 
    4.687934, 4.686851, 4.689076, 4.701419, 4.722225, 4.749526, 4.781257, 
    4.815298, 4.849463, 4.8815, 4.909118, 4.930127, 4.942695, 4.945752, 
    4.939439, 4.925432, 4.906913, 4.88804, 4.873039, 4.865275, 4.866679,
  // momentumY(13,29, 0-49)
    5.057277, 5.025501, 4.993886, 4.963425, 4.935068, 4.909718, 4.888201, 
    4.871215, 4.859243, 4.852449, 4.850572, 4.852848, 4.858019, 4.864477, 
    4.870577, 0, 4.960837, 4.965211, 4.967146, 4.96498, 4.957272, 4.937307, 
    4.911318, 4.878489, 4.841214, 4.801627, 4.763185, 4.72964, 4.705064, 
    4.691149, 4.690714, 4.694875, 4.708726, 4.730634, 4.758652, 4.790708, 
    4.824646, 4.858231, 4.889145, 4.915062, 4.933808, 4.943669, 4.943821, 
    4.934777, 4.918635, 4.898928, 4.87997, 4.865904, 4.859822, 4.863319,
  // momentumY(13,30, 0-49)
    5.059418, 5.028654, 4.997622, 4.96715, 4.938057, 4.911136, 4.887138, 
    4.866747, 4.850553, 4.839038, 4.832601, 4.831628, 4.836618, 4.848354, 
    4.867994, 4.90837, 4.928143, 4.951606, 4.967244, 4.973113, 4.968354, 
    4.949694, 4.92203, 4.886323, 4.846043, 4.804104, 4.764419, 4.730797, 
    4.707057, 4.694342, 4.694369, 4.700532, 4.715995, 4.739077, 4.76782, 
    4.800131, 4.833815, 4.866575, 4.896039, 4.919852, 4.935893, 4.942627, 
    4.93956, 4.927652, 4.909478, 4.888913, 4.870369, 4.857808, 4.853965, 
    4.860042,
  // momentumY(13,31, 0-49)
    5.060282, 5.029759, 4.999126, 4.96925, 4.940992, 4.915175, 4.892564, 
    4.873836, 4.859542, 4.850095, 4.845772, 4.846765, 4.85328, 4.865714, 
    4.884841, 4.905748, 4.911053, 4.932447, 4.945031, 4.948086, 4.941575, 
    4.923994, 4.898461, 4.866093, 4.830063, 4.792876, 4.758057, 4.729052, 
    4.709362, 4.699802, 4.701348, 4.710032, 4.727447, 4.751931, 4.781534, 
    4.814127, 4.847456, 4.879147, 4.906764, 4.927947, 4.940672, 4.94366, 
    4.936833, 4.921684, 4.90129, 4.879853, 4.861801, 4.850834, 4.849262, 
    4.857854,
  // momentumY(13,32, 0-49)
    5.060558, 5.030423, 5.000259, 4.970952, 4.943376, 4.918372, 4.896713, 
    4.879066, 4.865955, 4.857725, 4.854555, 4.856493, 4.863556, 4.875896, 
    4.894008, 4.900531, 4.896977, 4.915523, 4.924882, 4.9252, 4.916963, 
    4.900275, 4.876549, 4.847143, 4.815058, 4.782508, 4.752657, 4.728541, 
    4.713242, 4.707185, 4.710644, 4.721965, 4.741295, 4.766997, 4.797129, 
    4.829546, 4.861939, 4.891879, 4.916902, 4.9347, 4.943443, 4.94221, 
    4.931443, 4.913217, 4.891095, 4.869491, 4.85271, 4.844056, 4.845331, 
    4.856855,
  // momentumY(13,33, 0-49)
    5.059862, 5.03015, 5.000467, 4.971692, 4.944696, 4.920317, 4.899325, 
    4.882373, 4.869952, 4.862354, 4.859664, 4.861796, 4.868586, 4.879933, 
    4.896007, 4.893321, 4.885574, 4.900522, 4.906545, 4.904282, 4.894521, 
    4.878765, 4.856861, 4.8304, 4.802221, 4.774295, 4.749418, 4.730218, 
    4.719326, 4.716811, 4.722351, 4.736221, 4.757266, 4.783872, 4.814105, 
    4.845798, 4.876605, 4.904065, 4.925737, 4.939448, 4.943662, 4.93793, 
    4.923305, 4.902457, 4.879358, 4.858486, 4.843853, 4.838239, 4.842885, 
    4.857669,
  // momentumY(13,34, 0-49)
    5.058055, 5.028715, 4.999457, 4.971143, 4.944623, 4.920722, 4.900189, 
    4.883659, 4.871587, 4.864218, 4.861553, 4.863379, 4.869329, 4.879015, 
    4.892175, 4.88469, 4.876192, 4.887134, 4.889908, 4.885369, 4.874451, 
    4.859777, 4.839851, 4.816452, 4.79222, 4.768898, 4.748909, 4.734482, 
    4.727811, 4.728682, 4.736307, 4.752478, 4.774912, 4.802001, 4.831811, 
    4.862161, 4.890678, 4.914915, 4.93252, 4.941554, 4.94089, 4.930667, 
    4.912594, 4.889904, 4.866834, 4.847734, 4.836153, 4.834247, 4.842685, 
    4.860934,
  // momentumY(13,35, 0-49)
    5.055274, 5.02619, 4.997241, 4.969266, 4.943089, 4.919506, 4.899241, 
    4.882901, 4.870915, 4.863482, 4.860535, 4.861737, 4.866537, 4.874239, 
    4.884109, 4.875016, 4.868087, 4.875023, 4.874868, 4.868522, 4.85693, 
    4.843543, 4.825792, 4.805592, 4.785332, 4.766533, 4.751252, 4.741336, 
    4.738557, 4.742521, 4.752098, 4.770198, 4.793586, 4.820644, 4.849438, 
    4.87777, 4.90328, 4.923584, 4.936518, 4.940488, 4.934902, 4.920564, 
    4.899837, 4.876399, 4.854555, 4.838321, 4.830633, 4.832978, 4.845473, 
    4.86724,
  // momentumY(13,36, 0-49)
    5.051935, 5.022963, 4.994163, 4.966357, 4.940342, 4.916883, 4.896673, 
    4.880292, 4.868145, 4.860397, 4.856926, 4.857306, 4.860819, 4.866513, 
    4.873233, 4.864482, 4.860516, 4.863798, 4.861239, 4.853672, 4.841947, 
    4.830064, 4.814686, 4.797793, 4.781472, 4.767046, 4.756203, 4.750443, 
    4.751133, 4.757798, 4.76908, 4.788637, 4.812456, 4.838905, 4.86604, 
    4.891673, 4.9135, 4.929286, 4.937158, 4.935996, 4.925839, 4.908185, 
    4.885969, 4.863123, 4.843789, 4.831448, 4.828336, 4.835277, 4.851907, 
    4.87708,
  // momentumY(13,37, 0-49)
    5.048712, 5.019714, 4.990895, 4.963061, 4.936992, 4.91342, 4.893018, 
    4.876333, 4.863755, 4.855429, 4.851202, 4.850588, 4.852764, 4.856591, 
    4.860627, 4.853176, 4.852786, 4.853034, 4.848742, 4.840593, 4.829271, 
    4.819106, 4.806266, 4.79274, 4.780269, 4.769989, 4.763242, 4.761208, 
    4.764874, 4.773776, 4.78642, 4.806883, 4.830554, 4.855775, 4.880613, 
    4.902925, 4.920528, 4.931437, 4.934191, 4.928248, 4.914334, 4.894584, 
    4.87234, 4.851547, 4.83594, 4.828331, 4.830231, 4.841869, 4.862504, 
    4.890805,
  // momentumY(13,38, 0-49)
    5.046463, 5.017363, 4.988382, 4.960333, 4.933984, 4.910048, 4.889175, 
    4.871894, 4.858581, 4.849375, 4.84412, 4.842312, 4.843084, 4.84521, 
    4.847122, 4.841239, 4.84439, 4.842373, 4.837064, 4.828948, 4.818515, 
    4.810253, 4.800081, 4.789934, 4.781161, 4.774736, 4.771679, 4.772884, 
    4.778982, 4.789603, 4.803183, 4.82395, 4.846866, 4.87026, 4.892232, 
    4.910744, 4.923823, 4.92984, 4.927855, 4.917969, 4.901567, 4.881282, 
    4.860622, 4.843279, 4.832405, 4.830073, 4.83712, 4.853296, 4.877594, 
    4.908586,
  // momentumY(13,39, 0-49)
    5.046107, 5.016935, 4.987735, 4.959342, 4.932527, 4.907993, 4.886375, 
    4.86819, 4.853814, 4.843393, 4.836789, 4.833525, 4.832754, 4.833261, 
    4.833495, 4.82901, 4.835154, 4.83167, 4.826, 4.818432, 4.809279, 
    4.803062, 4.795628, 4.788808, 4.783522, 4.780604, 4.780778, 4.78469, 
    4.79264, 4.804419, 4.818454, 4.838909, 4.860484, 4.881526, 4.900217, 
    4.914691, 4.92329, 4.924838, 4.918981, 4.90646, 4.889201, 4.870115, 
    4.852602, 4.839882, 4.834409, 4.837548, 4.849568, 4.869874, 4.897309, 
    4.930414,
  // momentumY(13,40, 0-49)
    5.048494, 5.019421, 4.990073, 4.961317, 4.933938, 4.90864, 4.886052, 
    4.866689, 4.850931, 4.838945, 4.830641, 4.8256, 4.823055, 4.82189, 
    4.82068, 4.817156, 4.825377, 4.821116, 4.815586, 4.808927, 4.801313, 
    4.797197, 4.792489, 4.788867, 4.786796, 4.786984, 4.789888, 4.795939, 
    4.805148, 4.817516, 4.831503, 4.85106, 4.870792, 4.889106, 4.904329, 
    4.914861, 4.919432, 4.917396, 4.908987, 4.895493, 4.879183, 4.862983, 
    4.84994, 4.842655, 4.842869, 4.851325, 4.86787, 4.891695, 4.921583, 
    4.956109,
  // momentumY(13,41, 0-49)
    5.05427, 5.025635, 4.996369, 4.967378, 4.939467, 4.913352, 4.889659, 
    4.868913, 4.851506, 4.837645, 4.827295, 4.820136, 4.815523, 4.812502, 
    4.809849, 4.806692, 4.81588, 4.811314, 4.806209, 4.800623, 4.794641, 
    4.79257, 4.790468, 4.789821, 4.790624, 4.793467, 4.798572, 4.806185, 
    4.816072, 4.828482, 4.841944, 4.860108, 4.877642, 4.893072, 4.90494, 
    4.911988, 4.913404, 4.909066, 4.899735, 4.887073, 4.87345, 4.861562, 
    4.85393, 4.852476, 4.858293, 4.871628, 4.892047, 4.918634, 4.950186, 
    4.985343,
  // momentumY(13,42, 0-49)
    5.063781, 5.036088, 5.007306, 4.978371, 4.950112, 4.923259, 4.898448, 
    4.876221, 4.856994, 4.841022, 4.828345, 4.818758, 4.811777, 4.806639, 
    4.802362, 4.798909, 4.80793, 4.803259, 4.798624, 4.794068, 4.789628, 
    4.789413, 4.789672, 4.791672, 4.794939, 4.799946, 4.806708, 4.815324, 
    4.825358, 4.837329, 4.84987, 4.866296, 4.881484, 4.894133, 4.903078, 
    4.907446, 4.906895, 4.90178, 4.893241, 4.883102, 4.873612, 4.867048, 
    4.865321, 4.869707, 4.880752, 4.898339, 4.921859, 4.950371, 4.982732, 
    5.017666,
  // momentumY(13,43, 0-49)
    5.077024, 5.050926, 5.02318, 4.994742, 4.966463, 4.939089, 4.913278, 
    4.889596, 4.868496, 4.850291, 4.835114, 4.822883, 4.813281, 4.80576, 
    4.799586, 4.79519, 4.80303, 4.798201, 4.793865, 4.790109, 4.786953, 
    4.788271, 4.790523, 4.794739, 4.799999, 4.80666, 4.814556, 4.823662, 
    4.8334, 4.84456, 4.855913, 4.87045, 4.883365, 4.893603, 4.900323, 
    4.903059, 4.901888, 4.897532, 4.891333, 4.885078, 4.880715, 4.880008, 
    4.884263, 4.894188, 4.909894, 4.931011, 4.956826, 4.986413, 5.018707, 
    5.052526,
  // momentumY(13,44, 0-49)
    5.09363, 5.069897, 5.04386, 5.016483, 4.988629, 4.96107, 4.934496, 
    4.909508, 4.886611, 4.866188, 4.848468, 4.833498, 4.82113, 4.811025, 
    4.802682, 4.796786, 4.802666, 4.797429, 4.793074, 4.789756, 4.787496, 
    4.789924, 4.7937, 4.79963, 4.806377, 4.814182, 4.822727, 4.831895, 
    4.841009, 4.85113, 4.861181, 4.873878, 4.884815, 4.893214, 4.898576, 
    4.900804, 4.900312, 4.898042, 4.895368, 4.893885, 4.895139, 4.900371, 
    4.910341, 4.925292, 4.945001, 4.968908, 4.996238, 5.026088, 5.057459, 
    5.089253,
  // momentumY(13,45, 0-49)
    5.112896, 5.092362, 5.068785, 5.043111, 5.016217, 4.988903, 4.961903, 
    4.935873, 4.911382, 4.88889, 4.868727, 4.851068, 4.835922, 4.823139, 
    4.812431, 4.804618, 4.808037, 4.802051, 4.79729, 4.793986, 4.792167, 
    4.79523, 4.800014, 4.807119, 4.814841, 4.823317, 4.832101, 4.841004, 
    4.8493, 4.858297, 4.867085, 4.878168, 4.887572, 4.894811, 4.899705, 
    4.902462, 4.903721, 4.904501, 4.906074, 4.909746, 4.916643, 4.927522, 
    4.942692, 4.962025, 4.985044, 5.011038, 5.039169, 5.068532, 5.098169, 
    5.127051,
  // momentumY(13,46, 0-49)
    5.133814, 5.117327, 5.096988, 5.073705, 5.048361, 5.021798, 4.994802, 
    4.968101, 4.942336, 4.918055, 4.895684, 4.87552, 4.857718, 4.842292, 
    4.829139, 4.81916, 4.819887, 4.812812, 4.807271, 4.803571, 4.801742, 
    4.80497, 4.81025, 4.818002, 4.826226, 4.834962, 4.843659, 4.852087, 
    4.859497, 4.867418, 4.875102, 4.884908, 4.893291, 4.900041, 4.905254, 
    4.909355, 4.913095, 4.917461, 4.923537, 4.932306, 4.944498, 4.960462, 
    4.980148, 5.003146, 5.028774, 5.056185, 5.084462, 5.112659, 5.139817, 
    5.164942,
  // momentumY(13,47, 0-49)
    5.155118, 5.143477, 5.127144, 5.10696, 5.083807, 5.058568, 5.032099, 
    5.005201, 4.978597, 4.952922, 4.928703, 4.906341, 4.886123, 4.868207, 
    4.85265, 4.840416, 4.838448, 4.830011, 4.823393, 4.818952, 4.816723, 
    4.819705, 4.825018, 4.832941, 4.841257, 4.849924, 4.85831, 4.866159, 
    4.872729, 4.879717, 4.886525, 4.895436, 4.903288, 4.910117, 4.91623, 
    4.922192, 4.928778, 4.936869, 4.947312, 4.960783, 4.977658, 4.997964, 
    5.021375, 5.047264, 5.074781, 5.102951, 5.130748, 5.157147, 5.181139, 
    5.201734,
  // momentumY(13,48, 0-49)
    5.17534, 5.169244, 5.157641, 5.141272, 5.120998, 5.09774, 5.072417, 
    5.045903, 5.019007, 4.992444, 4.966833, 4.942678, 4.920383, 4.900235, 
    4.882427, 4.867987, 4.863477, 4.85351, 4.845624, 4.840209, 4.837288, 
    4.839696, 4.844657, 4.852349, 4.860429, 4.868786, 4.876736, 4.884, 
    4.889857, 4.896114, 4.9023, 4.910675, 4.918396, 4.925701, 4.933056, 
    4.941097, 4.950563, 4.962187, 4.976577, 4.994122, 5.014909, 5.038708, 
    5.064978, 5.092928, 5.121566, 5.149796, 5.176466, 5.200438, 5.22062, 5.236,
  // momentumY(13,49, 0-49)
    5.18919, 5.190837, 5.186273, 5.175988, 5.160712, 5.141308, 5.11869, 
    5.09377, 5.067405, 5.04039, 5.013444, 4.987204, 4.962228, 4.938995, 
    4.917903, 4.901022, 4.900822, 4.888001, 4.877112, 4.869137, 4.864331, 
    4.86836, 4.875689, 4.886596, 4.896372, 4.905116, 4.911828, 4.916348, 
    4.917615, 4.919777, 4.922395, 4.930235, 4.938002, 4.946137, 4.955254, 
    4.966011, 4.979034, 4.994824, 5.013668, 5.035591, 5.060346, 5.087408, 
    5.116018, 5.145223, 5.173903, 5.200845, 5.22479, 5.244488, 5.258783, 
    5.266685,
  // momentumY(14,0, 0-49)
    5.229131, 5.206501, 5.178502, 5.14638, 5.111412, 5.074858, 5.037918, 
    5.001689, 4.967128, 4.935019, 4.905952, 4.880305, 4.858244, 4.839743, 
    4.824595, 4.812624, 4.804584, 4.797328, 4.792109, 4.788625, 4.78663, 
    4.786323, 4.787329, 4.789779, 4.793612, 4.798909, 4.805624, 4.813658, 
    4.822749, 4.832749, 4.84324, 4.854219, 4.865003, 4.875406, 4.885445, 
    4.89538, 4.905724, 4.917185, 4.930576, 4.94668, 4.966119, 4.989237, 
    5.016041, 5.046188, 5.079033, 5.113686, 5.149096, 5.184103, 5.21749, 
    5.247988,
  // momentumY(14,1, 0-49)
    5.207026, 5.182279, 5.152763, 5.119683, 5.084245, 5.047626, 5.010942, 
    4.975212, 4.941328, 4.910021, 4.881835, 4.857101, 4.835941, 4.818269, 
    4.80382, 4.79253, 4.786399, 4.779195, 4.773937, 4.770339, 4.768142, 
    4.767947, 4.769014, 4.771609, 4.775563, 4.781028, 4.787959, 4.796264, 
    4.805616, 4.816019, 4.826934, 4.838686, 4.850087, 4.860837, 4.870841, 
    4.880264, 4.889561, 4.899436, 4.910755, 4.924414, 4.941188, 4.961601, 
    4.985838, 5.013726, 5.044766, 5.078192, 5.113054, 5.148269, 5.182673, 
    5.215027,
  // momentumY(14,2, 0-49)
    5.183304, 5.15703, 5.12666, 5.093325, 5.058139, 5.022183, 4.986475, 
    4.951942, 4.919401, 4.889516, 4.862769, 4.839439, 4.819584, 4.803053, 
    4.789515, 4.779003, 4.774808, 4.767579, 4.762142, 4.758224, 4.755566, 
    4.755175, 4.755948, 4.758294, 4.761974, 4.767229, 4.774033, 4.782334, 
    4.791769, 4.802477, 4.813826, 4.826488, 4.838775, 4.850249, 4.860665, 
    4.870028, 4.878657, 4.887173, 4.896429, 4.907394, 4.921, 4.937978, 
    4.958755, 4.983394, 5.011603, 5.042788, 5.076122, 5.110613, 5.14515, 
    5.178529,
  // momentumY(14,3, 0-49)
    5.159269, 5.132011, 5.101366, 5.068372, 5.034046, 4.999361, 4.965226, 
    4.932481, 4.901851, 4.873924, 4.849108, 4.82761, 4.809415, 4.794293, 
    4.781828, 4.772121, 4.769814, 4.762452, 4.756672, 4.752212, 4.748813, 
    4.747893, 4.747982, 4.749643, 4.752614, 4.757233, 4.763523, 4.771494, 
    4.780782, 4.791656, 4.803401, 4.817072, 4.830497, 4.84309, 4.854418, 
    4.864275, 4.872768, 4.880341, 4.887757, 4.896002, 4.906137, 4.919126, 
    4.935688, 4.956191, 4.980619, 5.008601, 5.039472, 5.072342, 5.106161, 
    5.139763,
  // momentumY(14,4, 0-49)
    5.136073, 5.108289, 5.077836, 5.045656, 5.012658, 4.979708, 4.947617, 
    4.91712, 4.888855, 4.863318, 4.840836, 4.821526, 4.805284, 4.791785, 
    4.780509, 4.771574, 4.771007, 4.763416, 4.75714, 4.751925, 4.747519, 
    4.745743, 4.744758, 4.745288, 4.747094, 4.75062, 4.755964, 4.763226, 
    4.772083, 4.782914, 4.794947, 4.809652, 4.824399, 4.838461, 4.851204, 
    4.862165, 4.871171, 4.878408, 4.884452, 4.890225, 4.896865, 4.905565, 
    4.917366, 4.933001, 4.952807, 4.976699, 5.004219, 5.034612, 5.066907, 
    5.099984,
  // momentumY(14,5, 0-49)
    5.114647, 5.08669, 5.056768, 5.025724, 4.994371, 4.96347, 4.933736, 
    4.905807, 4.880225, 4.857395, 4.837543, 4.82069, 4.806624, 4.794909, 
    4.784913, 4.776653, 4.77757, 4.769712, 4.76284, 4.756712, 4.751087, 
    4.748175, 4.745767, 4.744746, 4.744943, 4.746911, 4.750852, 4.756979, 
    4.765056, 4.775557, 4.787667, 4.803314, 4.819453, 4.835233, 4.849818, 
    4.862471, 4.872696, 4.88035, 4.885726, 4.889578, 4.893041, 4.89748, 
    4.90426, 4.914527, 4.929033, 4.948059, 4.97142, 4.998543, 5.028562, 
    5.060421,
  // momentumY(14,6, 0-49)
    5.095639, 5.06775, 5.038558, 5.008825, 4.979269, 4.950567, 4.923344, 
    4.898149, 4.875429, 4.855488, 4.838451, 4.824225, 4.812485, 4.802677, 
    4.79404, 4.786319, 4.788359, 4.780312, 4.772842, 4.76574, 4.758781, 
    4.754543, 4.750437, 4.747506, 4.745694, 4.74566, 4.747729, 4.752261, 
    4.759154, 4.768952, 4.780826, 4.797183, 4.814626, 4.832209, 4.848913, 
    4.86374, 4.875854, 4.884737, 4.890322, 4.893084, 4.894041, 4.894635, 
    4.896505, 4.901212, 4.909982, 4.923539, 4.942053, 4.9652, 4.992265, 
    5.022275,
  // momentumY(14,7, 0-49)
    5.079382, 5.051685, 5.023293, 4.994893, 4.967136, 4.940629, 4.915915, 
    4.893468, 4.873641, 4.856643, 4.842487, 4.830967, 4.821641, 4.813837, 
    4.806674, 4.799337, 4.802044, 4.794051, 4.786124, 4.778114, 4.769837, 
    4.764191, 4.758224, 4.753119, 4.748968, 4.746531, 4.746279, 4.748741, 
    4.754, 4.762649, 4.773867, 4.790557, 4.809045, 4.82832, 4.847221, 
    4.864514, 4.879047, 4.889917, 4.896648, 4.899345, 4.898779, 4.896335, 
    4.893821, 4.893167, 4.896089, 4.903821, 4.916978, 4.935566, 4.959084, 
    4.986681,
  // momentumY(14,8, 0-49)
    5.065872, 5.038401, 5.01076, 4.983597, 4.95751, 4.933054, 4.910717, 
    4.890898, 4.87387, 4.859747, 4.848433, 4.839616, 4.832747, 4.827052, 
    4.821545, 4.814451, 4.817304, 4.809798, 4.801712, 4.793008, 4.783563, 
    4.776557, 4.76869, 4.761254, 4.754529, 4.749352, 4.746367, 4.746292, 
    4.749443, 4.756443, 4.766504, 4.783024, 4.80213, 4.822789, 4.843732, 
    4.863547, 4.880808, 4.894256, 4.903001, 4.906718, 4.905815, 4.901471, 
    4.895508, 4.890118, 4.887469, 4.889338, 4.896865, 4.91048, 4.92997, 
    4.954655,
  // momentumY(14,9, 0-49)
    5.054821, 5.027532, 5.000518, 4.974404, 4.949765, 4.927123, 4.906926, 
    4.889516, 4.875094, 4.863682, 4.855093, 4.848915, 4.84452, 4.841063, 
    4.837492, 4.83054, 4.83301, 4.826586, 4.818791, 4.809748, 4.799422, 
    4.791223, 4.781535, 4.77173, 4.762289, 4.754117, 4.748044, 4.744996, 
    4.74556, 4.750387, 4.75874, 4.774489, 4.79366, 4.815218, 4.837843, 
    4.859991, 4.880027, 4.896397, 4.907828, 4.913559, 4.913555, 4.908646, 
    4.9005, 4.891405, 4.883876, 4.880214, 4.88213, 4.890561, 4.905677, 
    4.927028,
  // momentumY(14,10, 0-49)
    5.04573, 5.018534, 4.991975, 4.96668, 4.943219, 4.922101, 4.903752, 
    4.888469, 4.876389, 4.867462, 4.861423, 4.857787, 4.855875, 4.854819, 
    4.85357, 4.846726, 4.848333, 4.843694, 4.836761, 4.827849, 4.817042, 
    4.807907, 4.796583, 4.784479, 4.772281, 4.760951, 4.751504, 4.745098, 
    4.742626, 4.744754, 4.750842, 4.765165, 4.783755, 4.805612, 4.829389, 
    4.853467, 4.876074, 4.895433, 4.909956, 4.918473, 4.920488, 4.916383, 
    4.907503, 4.896041, 4.8847, 4.876213, 4.872857, 4.876142, 4.886695, 
    4.904379,
  // momentumY(14,11, 0-49)
    5.038, 5.010782, 4.984499, 4.959789, 4.937232, 4.917344, 4.900531, 
    4.887064, 4.877037, 4.870335, 4.866637, 4.86542, 4.865989, 4.867517, 
    4.869044, 4.862404, 4.862796, 4.860651, 4.855209, 4.846973, 4.836166, 
    4.826419, 4.813724, 4.799486, 4.784587, 4.770025, 4.757013, 4.746933, 
    4.741017, 4.73996, 4.74325, 4.755486, 4.772819, 4.794303, 4.818602, 
    4.844064, 4.868836, 4.890996, 4.908724, 4.92051, 4.925418, 4.923341, 
    4.915177, 4.902844, 4.889031, 4.87675, 4.86878, 4.867208, 4.873197, 
    4.886992,
  // momentumY(14,12, 0-49)
    5.031034, 5.003688, 4.977518, 4.953181, 4.931284, 4.912348, 4.896778, 
    4.884824, 4.876548, 4.871799, 4.870219, 4.871272, 4.8743, 4.878574, 
    4.883319, 4.877185, 4.876233, 4.87719, 4.873849, 4.866863, 4.856576, 
    4.846573, 4.832829, 4.816703, 4.799254, 4.781491, 4.764815, 4.750834, 
    4.741136, 4.736468, 4.736497, 4.746009, 4.761425, 4.781863, 4.806017, 
    4.832239, 4.858638, 4.883218, 4.904005, 4.919235, 4.927595, 4.928498, 
    4.922335, 4.910599, 4.895769, 4.880947, 4.869279, 4.863392, 4.865007, 
    4.874826,
  // momentumY(14,13, 0-49)
    5.024333, 4.99677, 4.970584, 4.946457, 4.925018, 4.906796, 4.892203, 
    4.881479, 4.874665, 4.87159, 4.871881, 4.875025, 4.880433, 4.887527, 
    4.895803, 4.890821, 4.888721, 4.893181, 4.89245, 4.887251, 4.878012, 
    4.868104, 4.853672, 4.835969, 4.816206, 4.795377, 4.775051, 4.757049, 
    4.743318, 4.734697, 4.731096, 4.73732, 4.750211, 4.768974, 4.792344, 
    4.818688, 4.846123, 4.872623, 4.896131, 4.91471, 4.926751, 4.931248, 
    4.928075, 4.918214, 4.903775, 4.887743, 4.873465, 4.864006, 4.861628, 
    4.867535,
  // momentumY(14,14, 0-49)
    5.017553, 4.989715, 4.963422, 4.939384, 4.918242, 4.90054, 4.88669, 
    4.876932, 4.871295, 4.869604, 4.871495, 4.876493, 4.884107, 4.893934, 
    4.905785, 4.903114, 4.900491, 4.908577, 4.910793, 4.907833, 4.900127, 
    4.890634, 4.875879, 4.856959, 4.835193, 4.811535, 4.787686, 4.765656, 
    4.747746, 4.734937, 4.727468, 4.729933, 4.739788, 4.756329, 4.778342, 
    4.804221, 4.832108, 4.85998, 4.88575, 4.90738, 4.923053, 4.931413, 
    4.931864, 4.92485, 4.912005, 4.896032, 4.880286, 4.868128, 4.8623, 
    4.864512,
  // momentumY(14,15, 0-49)
    5.010522, 4.982379, 4.955929, 4.931895, 4.910927, 4.893575, 4.880256, 
    4.871205, 4.866455, 4.865833, 4.869004, 4.875539, 4.885052, 4.897312, 
    4.912402, 4.913854, 4.911866, 4.923392, 4.928685, 4.928277, 4.922505, 
    4.913686, 4.898948, 4.879184, 4.855774, 4.829604, 4.802463, 4.776515, 
    4.754398, 4.737293, 4.725864, 4.724226, 4.730651, 4.744537, 4.764725, 
    4.789639, 4.817448, 4.846156, 4.873679, 4.897934, 4.916968, 4.929162, 
    4.933515, 4.929967, 4.919626, 4.90479, 4.888655, 4.874717, 4.866093, 
    4.864969,
  // momentumY(14,16, 0-49)
    5.003232, 4.974789, 4.948159, 4.924067, 4.903166, 4.886005, 4.872997, 
    4.864381, 4.860195, 4.860283, 4.864339, 4.872, 4.882958, 4.897115, 
    4.91473, 4.922801, 4.923217, 4.937708, 4.946001, 4.948301, 4.94475, 
    4.936777, 4.92233, 4.902053, 4.877351, 4.849022, 4.818892, 4.789238, 
    4.76301, 4.74164, 4.726334, 4.720396, 4.723143, 4.734078, 4.752094, 
    4.775647, 4.802935, 4.831992, 4.860762, 4.887154, 4.909132, 4.924897, 
    4.93313, 4.933318, 4.926054, 4.91317, 4.897569, 4.882729, 4.872013, 
    4.868022,
  // momentumY(14,17, 0-49)
    4.995819, 4.967114, 4.940305, 4.916105, 4.895159, 4.878008, 4.865059, 
    4.856553, 4.85254, 4.852895, 4.857356, 4.865614, 4.877438, 4.892803, 
    4.912023, 4.929695, 4.934912, 4.951701, 4.962767, 4.967796, 4.966612, 
    4.959546, 4.945543, 4.924974, 4.899243, 4.869065, 4.836262, 4.803187, 
    4.773059, 4.747612, 4.728692, 4.718437, 4.717418, 4.725255, 4.740889, 
    4.762807, 4.789228, 4.818224, 4.84777, 4.875792, 4.900223, 4.919144, 
    4.930996, 4.934896, 4.930968, 4.920557, 4.906198, 4.891222, 4.879112, 
    4.872787,
  // momentumY(14,18, 0-49)
    4.988537, 4.959641, 4.932666, 4.9083, 4.887167, 4.869789, 4.856569, 
    4.847752, 4.843416, 4.843479, 4.847744, 4.855983, 4.868048, 4.88397, 
    4.904027, 4.934335, 4.947203, 4.965634, 4.979208, 4.98692, 4.988139, 
    4.981914, 4.968329, 4.947478, 4.920774, 4.888891, 4.85365, 4.81746, 
    4.783762, 4.754593, 4.73253, 4.71814, 4.713455, 4.718208, 4.731387, 
    4.75151, 4.776821, 4.805424, 4.835332, 4.864502, 4.890868, 4.912439, 
    4.927494, 4.934857, 4.934252, 4.926565, 4.913923, 4.899424, 4.88655, 
    4.878451,
  // momentumY(14,19, 0-49)
    4.981731, 4.952747, 4.925626, 4.901007, 4.879478, 4.86154, 4.847589, 
    4.837891, 4.832567, 4.831611, 4.834948, 4.842501, 4.854297, 4.870481, 
    4.891221, 4.936656, 4.959976, 4.979749, 4.995747, 5.00617, 5.009804, 
    5.004245, 4.990828, 4.969369, 4.941361, 4.907585, 4.869937, 4.830897, 
    4.794071, 4.761743, 4.73723, 4.719127, 4.711077, 4.712924, 4.723711, 
    4.741991, 4.766041, 4.793996, 4.823914, 4.853789, 4.881576, 4.90526, 
    4.923007, 4.933437, 4.93594, 4.930997, 4.920331, 4.906754, 4.893658, 
    4.88432,
  // momentumY(14,20, 0-49)
    4.975356, 4.946013, 4.918895, 4.894783, 4.874384, 4.858284, 4.846906, 
    4.840438, 4.838765, 4.841401, 4.847481, 4.8558, 4.864954, 4.87357, 
    4.880587, 0, 4.989855, 4.995119, 5.000073, 5.003455, 5.004048, 4.997201, 
    4.985688, 4.96794, 4.944427, 4.914887, 4.880343, 4.842763, 4.805717, 
    4.771926, 4.745841, 4.724278, 4.712812, 4.711535, 4.719627, 4.735713, 
    4.758105, 4.784973, 4.814407, 4.844437, 4.873043, 4.898208, 4.918039, 
    4.931002, 4.936229, 4.933856, 4.92523, 4.912845, 4.899946, 4.889857,
  // momentumY(14,21, 0-49)
    4.970289, 4.941153, 4.914182, 4.890114, 4.869606, 4.853193, 4.841239, 
    4.833877, 4.830952, 4.831978, 4.836136, 4.842323, 4.849247, 4.85558, 
    4.860119, 0, 5.006929, 5.011988, 5.017016, 5.020457, 5.020889, 5.011185, 
    4.997466, 4.977767, 4.952747, 4.922137, 4.886837, 4.848618, 4.81087, 
    4.776311, 4.749987, 4.726534, 4.71325, 4.710298, 4.716912, 4.731764, 
    4.753213, 4.779468, 4.808661, 4.838869, 4.868112, 4.894393, 4.915797, 
    4.930689, 4.938019, 4.937646, 4.930596, 4.919082, 4.906178, 4.895215,
  // momentumY(14,22, 0-49)
    4.96617, 4.937153, 4.910255, 4.886184, 4.865558, 4.848874, 4.83646, 
    4.828418, 4.824572, 4.824438, 4.827231, 4.831902, 4.837212, 4.841824, 
    4.844385, 0, 5.018405, 5.023205, 5.02841, 5.032224, 5.033048, 5.021325, 
    5.00638, 4.985718, 4.960042, 4.928993, 4.893322, 4.85464, 4.816243, 
    4.780902, 4.754295, 4.728978, 4.713942, 4.709406, 4.71464, 4.728346, 
    4.748909, 4.774562, 4.803468, 4.833735, 4.863416, 4.890533, 4.913163, 
    4.929612, 4.938688, 4.940041, 4.934431, 4.923813, 4.911096, 4.899575,
  // momentumY(14,23, 0-49)
    4.96328, 4.934348, 4.907502, 4.883425, 4.862714, 4.845841, 4.833112, 
    4.824607, 4.820145, 4.819244, 4.821142, 4.824821, 4.829068, 4.832527, 
    4.833734, 0, 5.025937, 5.030453, 5.035746, 5.039857, 5.041064, 5.027761, 
    5.011934, 4.990608, 4.964503, 4.9332, 4.897349, 4.85845, 4.819719, 
    4.783957, 4.757343, 4.730652, 4.714336, 4.708647, 4.712873, 4.725742, 
    4.745659, 4.770877, 4.799579, 4.829896, 4.859901, 4.887634, 4.911168, 
    4.928766, 4.939146, 4.941798, 4.937283, 4.927362, 4.914799, 4.902847,
  // momentumY(14,24, 0-49)
    4.961791, 4.932945, 4.906162, 4.882113, 4.861383, 4.844429, 4.831546, 
    4.822805, 4.81802, 4.816717, 4.818145, 4.821302, 4.824994, 4.827858, 
    4.828371, 0, 5.029955, 5.034287, 5.039621, 5.043921, 5.045398, 5.031094, 
    5.014718, 4.992973, 4.966591, 4.935138, 4.899226, 4.8603, 4.821521, 
    4.785698, 4.759323, 4.731932, 4.714949, 4.708636, 4.712295, 4.724666, 
    4.744171, 4.76908, 4.797589, 4.827847, 4.857946, 4.88594, 4.909908, 
    4.928101, 4.939186, 4.942573, 4.93871, 4.929234, 4.916815, 4.904671,
  // momentumY(14,25, 0-49)
    4.961771, 4.933026, 4.906334, 4.882361, 4.86169, 4.844777, 4.831912, 
    4.823165, 4.818351, 4.816997, 4.818359, 4.821449, 4.825079, 4.827899, 
    4.828384, 0, 5.03003, 5.034381, 5.039783, 5.044186, 5.045787, 5.031203, 
    5.014672, 4.992793, 4.966319, 4.934835, 4.89897, 4.860161, 4.821557, 
    4.785944, 4.759897, 4.732482, 4.715449, 4.709057, 4.712609, 4.724858, 
    4.744236, 4.769025, 4.797433, 4.827615, 4.857674, 4.88567, 4.909687, 
    4.927975, 4.939195, 4.942734, 4.939016, 4.929639, 4.917246, 4.905041,
  // momentumY(14,26, 0-49)
    4.963167, 4.93454, 4.907962, 4.884112, 4.863579, 4.846827, 4.834151, 
    4.825628, 4.821076, 4.820027, 4.821736, 4.825215, 4.829287, 4.832619, 
    4.833757, 0, 5.026039, 5.030636, 5.036156, 5.040594, 5.042174, 5.028095, 
    5.011848, 4.990179, 4.963848, 4.932496, 4.896807, 4.858271, 4.820046, 
    4.784883, 4.759194, 4.73243, 4.715955, 4.710011, 4.713904, 4.726387, 
    4.745905, 4.770749, 4.799131, 4.829207, 4.85908, 4.886809, 4.91048, 
    4.928358, 4.939132, 4.942234, 4.938139, 4.928508, 4.91602, 4.903892,
  // momentumY(14,27, 0-49)
    4.965813, 4.937301, 4.910845, 4.887145, 4.866809, 4.850321, 4.837995, 
    4.829924, 4.825934, 4.825562, 4.828056, 4.832419, 4.837465, 4.841897, 
    4.844372, 0, 5.018102, 5.023104, 5.028753, 5.033145, 5.034584, 5.021748, 
    5.006234, 4.985136, 4.959219, 4.928194, 4.892848, 4.854764, 4.817146, 
    4.782689, 4.757411, 4.731923, 4.71657, 4.711563, 4.716202, 4.729245, 
    4.749143, 4.774192, 4.802603, 4.832528, 4.862057, 4.88924, 4.912171, 
    4.929139, 4.938899, 4.940991, 4.93603, 4.925817, 4.913135, 4.901226,
  // momentumY(14,28, 0-49)
    4.969423, 4.940984, 4.914621, 4.891065, 4.870954, 4.854809, 4.842978, 
    4.835584, 4.832475, 4.833191, 4.836968, 4.842775, 4.849395, 4.855551, 
    4.860049, 0, 5.006672, 5.0121, 5.017801, 5.022041, 5.023263, 5.01228, 
    4.997938, 4.977812, 4.952632, 4.922198, 4.887433, 4.850056, 4.81334, 
    4.779905, 4.755203, 4.731562, 4.717834, 4.714186, 4.719908, 4.733754, 
    4.754178, 4.779477, 4.80786, 4.837467, 4.866374, 4.892624, 4.914323, 
    4.929817, 4.937974, 4.938513, 4.932271, 4.921261, 4.908408, 4.896985,
  // momentumY(14,29, 0-49)
    4.973598, 4.945132, 4.91878, 4.895313, 4.875417, 4.859663, 4.848455, 
    4.841969, 4.840096, 4.842386, 4.848045, 4.855969, 4.864852, 4.873392, 
    4.88053, 0, 4.991336, 4.997087, 5.002714, 5.006726, 5.007765, 4.999115, 
    4.986455, 4.96784, 4.943899, 4.91449, 4.880672, 4.844324, 4.808808, 
    4.776659, 4.752664, 4.731198, 4.719398, 4.717382, 4.724414, 4.739241, 
    4.760315, 4.785926, 4.81427, 4.84347, 4.871576, 4.896624, 4.916734, 
    4.930334, 4.936449, 4.935032, 4.927205, 4.915243, 4.902236, 4.891462,
  // momentumY(14,30, 0-49)
    4.978459, 4.950448, 4.924171, 4.90026, 4.879285, 4.861737, 4.848003, 
    4.838342, 4.832888, 4.831677, 4.83469, 4.841944, 4.853562, 4.869802, 
    4.890952, 4.937116, 4.960141, 4.981357, 4.999086, 5.011297, 5.016665, 
    5.010939, 4.99806, 4.977265, 4.949973, 4.916874, 4.879813, 4.841241, 
    4.804756, 4.772696, 4.748902, 4.729621, 4.719982, 4.719895, 4.728523, 
    4.744562, 4.766439, 4.792431, 4.820715, 4.84939, 4.876489, 4.900041, 
    4.918213, 4.929551, 4.93329, 4.929682, 4.920183, 4.907356, 4.894434, 
    4.88467,
  // momentumY(14,31, 0-49)
    4.983125, 4.955338, 4.929348, 4.905835, 4.885411, 4.868597, 4.85578, 
    4.847207, 4.842966, 4.843014, 4.847225, 4.855464, 4.867691, 4.884041, 
    4.904872, 4.935839, 4.949141, 4.969279, 4.984799, 4.994443, 4.997485, 
    4.991339, 4.978379, 4.958244, 4.932343, 4.901263, 4.86675, 4.83112, 
    4.797772, 4.768725, 4.747015, 4.731064, 4.72435, 4.726704, 4.737257, 
    4.754694, 4.777433, 4.803735, 4.831755, 4.85956, 4.885167, 4.906618, 
    4.922161, 4.930507, 4.931175, 4.92478, 4.913159, 4.899173, 4.886178, 
    4.877337,
  // momentumY(14,32, 0-49)
    4.987358, 4.959856, 4.934148, 4.91095, 4.890905, 4.874556, 4.862307, 
    4.854393, 4.850876, 4.851655, 4.85653, 4.865274, 4.877754, 4.894031, 
    4.914469, 4.932961, 4.939357, 4.958105, 4.971329, 4.978452, 4.979202, 
    4.972534, 4.959299, 4.939528, 4.914677, 4.885373, 4.853353, 4.820845, 
    4.790998, 4.765457, 4.746442, 4.73423, 4.730731, 4.735687, 4.748199, 
    4.766947, 4.790341, 4.816634, 4.843962, 4.870373, 4.893885, 4.912594, 
    4.924883, 4.929708, 4.926944, 4.917631, 4.904008, 4.889196, 4.876601, 
    4.869208,
  // momentumY(14,33, 0-49)
    4.99063, 4.963439, 4.938015, 4.915095, 4.895347, 4.879332, 4.867464, 
    4.859974, 4.856893, 4.858074, 4.863241, 4.872085, 4.88437, 4.900063, 
    4.919447, 4.928698, 4.931004, 4.947732, 4.958413, 4.962972, 4.961474, 
    4.954248, 4.940749, 4.921361, 4.897592, 4.870147, 4.840767, 4.811585, 
    4.785475, 4.763719, 4.747799, 4.739508, 4.739332, 4.746913, 4.761318, 
    4.78121, 4.804995, 4.83091, 4.85707, 4.88152, 4.902306, 4.917626, 
    4.926063, 4.926908, 4.920468, 4.908258, 4.892908, 4.877741, 4.866107, 
    4.860717,
  // momentumY(14,34, 0-49)
    4.992525, 4.96564, 4.940499, 4.917854, 4.898386, 4.882666, 4.871113, 
    4.863943, 4.86116, 4.862561, 4.867793, 4.876443, 4.888147, 4.902713, 
    4.920231, 4.923387, 4.923928, 4.937998, 4.945892, 4.947875, 4.944241, 
    4.936496, 4.92287, 4.90407, 4.881607, 4.856267, 4.829761, 4.804101, 
    4.781861, 4.764022, 4.751439, 4.747082, 4.750193, 4.760307, 4.776446, 
    4.797251, 4.821106, 4.846224, 4.870707, 4.892605, 4.910032, 4.921345, 
    4.92542, 4.921961, 4.911783, 4.896895, 4.880278, 4.865354, 4.855299, 
    4.852454,
  // momentumY(14,35, 0-49)
    4.99278, 4.96617, 4.941314, 4.91896, 4.899793, 4.884388, 4.873153, 
    4.866287, 4.863753, 4.865289, 4.87046, 4.87873, 4.889587, 4.902627, 
    4.917654, 4.917314, 4.917788, 4.928729, 4.933709, 4.933207, 4.927653, 
    4.919489, 4.905965, 4.888046, 4.867195, 4.844253, 4.820849, 4.798853, 
    4.780519, 4.766601, 4.757459, 4.756906, 4.763144, 4.775598, 4.793231, 
    4.814648, 4.838199, 4.862067, 4.884343, 4.903111, 4.916597, 4.923395, 
    4.922756, 4.914888, 4.901155, 4.884047, 4.866805, 4.85282, 4.844973, 
    4.84515,
  // momentumY(14,36, 0-49)
    4.991346, 4.964972, 4.940395, 4.918357, 4.899533, 4.884483, 4.873598, 
    4.867045, 4.864746, 4.866374, 4.871405, 4.879189, 4.889049, 4.900362, 
    4.912611, 4.910634, 4.912133, 4.919724, 4.921842, 4.919075, 4.911914, 
    4.903495, 4.890347, 4.873635, 4.854704, 4.834425, 4.814302, 4.79603, 
    4.781533, 4.77143, 4.765703, 4.768709, 4.777803, 4.792308, 4.811116, 
    4.832782, 4.855612, 4.877761, 4.897319, 4.912441, 4.921529, 4.923491, 
    4.918043, 4.905955, 4.889152, 4.870528, 4.853456, 4.841154, 4.836089, 
    4.839647,
  // momentumY(14,37, 0-49)
    4.988453, 4.962273, 4.937971, 4.916267, 4.897817, 4.883152, 4.872628, 
    4.866377, 4.864271, 4.865924, 4.870734, 4.877946, 4.88674, 4.896296, 
    4.905811, 4.903345, 4.906444, 4.910737, 4.910229, 4.90555, 4.897175, 
    4.888714, 4.876239, 4.86105, 4.844311, 4.826896, 4.810146, 4.795563, 
    4.784745, 4.778251, 4.77579, 4.782004, 4.793592, 4.809768, 4.829356, 
    4.850853, 4.87252, 4.892492, 4.908888, 4.919978, 4.924416, 4.921508, 
    4.911499, 4.895743, 4.87667, 4.857455, 4.841446, 4.831538, 4.829711, 
    4.836845,
  // momentumY(14,38, 0-49)
    4.984639, 4.958626, 4.934591, 4.913228, 4.895154, 4.880854, 4.870646, 
    4.86461, 4.862578, 4.864117, 4.868563, 4.875087, 4.882763, 4.890626, 
    4.897676, 4.89531, 4.900163, 4.901466, 4.898746, 4.892606, 4.88346, 
    4.875215, 4.863713, 4.850336, 4.836003, 4.821574, 4.808197, 4.797181, 
    4.789793, 4.786611, 4.787156, 4.796136, 4.809761, 4.82715, 4.84706, 
    4.867931, 4.887993, 4.905383, 4.918293, 4.92518, 4.925019, 4.917578, 
    4.903661, 4.885168, 4.864916, 4.846192, 4.832146, 4.825239, 4.826932, 
    4.837641,
  // momentumY(14,39, 0-49)
    4.980752, 4.95491, 4.931138, 4.910096, 4.892348, 4.878327, 4.868291, 
    4.862281, 4.86009, 4.861258, 4.865097, 4.870739, 4.877207, 4.88346, 
    4.888396, 4.886341, 4.892785, 4.891613, 4.887215, 4.88012, 4.87067, 
    4.862928, 4.852697, 4.841382, 4.829606, 4.818201, 4.808114, 4.800452, 
    4.796173, 4.795929, 4.799117, 4.810341, 4.825474, 4.843554, 4.863278, 
    4.883053, 4.901103, 4.915614, 4.924913, 4.927712, 4.92337, 4.912158, 
    4.895406, 4.875451, 4.855321, 4.838219, 4.826949, 4.82348, 4.828774, 
    4.842854,
  // momentumY(14,40, 0-49)
    4.977879, 4.952263, 4.928766, 4.908001, 4.890475, 4.876557, 4.866449, 
    4.860152, 4.857441, 4.857857, 4.860724, 4.86519, 4.87028, 4.874952, 
    4.878095, 4.876329, 4.883979, 4.880965, 4.875467, 4.867936, 4.858642, 
    4.851704, 4.843017, 4.833961, 4.824832, 4.816414, 4.809454, 4.804865, 
    4.80331, 4.805566, 4.810947, 4.823834, 4.839893, 4.8581, 4.87712, 
    4.895356, 4.911077, 4.92258, 4.928399, 4.927567, 4.919873, 4.906066, 
    4.88791, 4.868001, 4.849374, 4.834966, 4.827127, 4.827327, 4.836097, 
    4.853168,
  // momentumY(14,41, 0-49)
    4.977243, 4.951975, 4.928784, 4.908237, 4.890777, 4.876709, 4.866188, 
    4.859186, 4.855484, 4.854657, 4.856086, 4.858981, 4.862435, 4.865462, 
    4.867022, 4.865379, 4.873715, 4.869505, 4.863459, 4.855964, 4.84724, 
    4.841386, 4.834473, 4.827814, 4.821355, 4.81582, 4.811758, 4.8099, 
    4.810643, 4.814913, 4.82198, 4.835919, 4.852301, 4.870073, 4.8879, 
    4.904237, 4.91746, 4.92605, 4.928823, 4.925181, 4.915336, 4.900439, 
    4.882529, 4.864255, 4.848449, 4.837637, 4.833674, 4.837571, 4.849523, 
    4.869064,
  // momentumY(14,42, 0-49)
    4.980048, 4.955317, 4.932497, 4.912102, 4.894521, 4.880002, 4.868662, 
    4.860474, 4.855247, 4.852629, 4.852093, 4.852965, 4.854447, 4.855668, 
    4.855711, 4.853931, 4.862373, 4.857519, 4.851374, 4.844295, 4.836475, 
    4.831925, 4.826941, 4.822737, 4.818897, 4.816074, 4.814629, 4.815122, 
    4.817711, 4.823489, 4.831711, 4.846095, 4.862226, 4.879052, 4.895293, 
    4.909513, 4.92027, 4.926304, 4.926771, 4.921447, 4.910919, 4.896608, 
    4.88063, 4.865476, 4.85361, 4.847065, 4.847208, 4.854662, 4.869378, 
    4.89079,
  // momentumY(14,43, 0-49)
    4.987293, 4.963366, 4.941016, 4.920723, 4.902826, 4.887541, 4.874972, 
    4.865113, 4.857836, 4.852889, 4.849873, 4.848258, 4.847405, 4.846586, 
    4.845038, 4.842797, 4.850761, 4.845643, 4.839696, 4.833277, 4.826568, 
    4.82345, 4.820451, 4.818665, 4.817314, 4.816969, 4.817812, 4.820253, 
    4.824242, 4.831039, 4.839899, 4.854184, 4.869569, 4.885051, 4.89946, 
    4.911537, 4.920093, 4.924184, 4.923324, 4.917646, 4.908003, 4.895916, 
    4.88339, 4.872587, 4.865491, 4.863626, 4.867915, 4.878666, 4.895671, 
    4.918324,
  // momentumY(14,44, 0-49)
    4.999643, 4.97684, 4.955107, 4.934894, 4.916515, 4.900183, 4.886018, 
    4.874065, 4.864291, 4.85656, 4.850628, 4.846134, 4.842605, 4.839487, 
    4.83618, 4.833108, 4.840065, 4.83484, 4.82921, 4.823539, 4.818005, 
    4.81632, 4.815243, 4.815725, 4.816647, 4.818492, 4.821272, 4.825261, 
    4.830235, 4.837609, 4.846658, 4.8604, 4.874674, 4.888574, 4.901094, 
    4.911215, 4.918052, 4.921008, 4.91994, 4.915264, 4.907966, 4.899511, 
    4.891633, 4.886055, 4.884239, 4.887223, 4.895544, 4.909267, 4.928077, 
    4.951357,
  // momentumY(14,45, 0-49)
    5.017312, 4.996, 4.97507, 4.95496, 4.935992, 4.918405, 4.902376, 4.88803, 
    4.875444, 4.864624, 4.855481, 4.847826, 4.841365, 4.835716, 4.83044, 
    4.826169, 4.831665, 4.826299, 4.820926, 4.815934, 4.811489, 4.81111, 
    4.811764, 4.814254, 4.81716, 4.820862, 4.825219, 4.830384, 4.835991, 
    4.843586, 4.852475, 4.865373, 4.878339, 4.890605, 4.901376, 4.909918, 
    4.915675, 4.918389, 4.918215, 4.915745, 4.911979, 4.908191, 4.905741, 
    4.90587, 4.909535, 4.917328, 4.92946, 4.945801, 4.965949, 4.989285,
  // momentumY(14,46, 0-49)
    5.040022, 5.0206, 5.000702, 4.98078, 4.9612, 4.942265, 4.924236, 
    4.907354, 4.891817, 4.877773, 4.865296, 4.854357, 4.84483, 4.83649, 
    4.829052, 4.823248, 4.82694, 4.821243, 4.81594, 4.811431, 4.807864, 
    4.808546, 4.810627, 4.814773, 4.819308, 4.82451, 4.8301, 4.836121, 
    4.842098, 4.849669, 4.858179, 4.870093, 4.881728, 4.892483, 4.901812, 
    4.909278, 4.914648, 4.917972, 4.919623, 4.920277, 4.920839, 4.922309, 
    4.92564, 4.931595, 4.94067, 4.953065, 4.968709, 4.987298, 5.008345, 
    5.031216,
  // momentumY(14,47, 0-49)
    5.067022, 5.049904, 5.031317, 5.011751, 4.991643, 4.971396, 4.951393, 
    4.931998, 4.913552, 4.896341, 4.880581, 4.866395, 4.853802, 4.842718, 
    4.832986, 4.825392, 4.827056, 4.820758, 4.815261, 4.810961, 4.807976, 
    4.809393, 4.812525, 4.817905, 4.823682, 4.830026, 4.836539, 4.843167, 
    4.849349, 4.856772, 4.86482, 4.875768, 4.8862, 4.89571, 4.904, 4.910928, 
    4.916553, 4.921173, 4.925306, 4.929629, 4.934891, 4.941786, 4.950864, 
    4.962459, 4.976653, 4.993308, 5.012097, 5.032546, 5.05407, 5.075994,
  // momentumY(14,48, 0-49)
    5.097138, 5.082759, 5.065822, 5.046871, 5.026447, 5.005077, 4.983285, 
    4.961578, 4.940433, 4.920274, 4.901444, 4.884194, 4.868665, 4.854891, 
    4.842824, 4.833281, 4.832807, 4.825633, 4.819666, 4.81528, 4.812549, 
    4.814342, 4.818109, 4.824279, 4.830903, 4.838052, 4.845232, 4.852296, 
    4.858621, 4.86589, 4.873518, 4.883643, 4.893113, 4.901714, 4.90939, 
    4.916262, 4.922637, 4.928999, 4.935947, 4.944109, 4.954046, 4.966163, 
    4.980648, 4.997454, 5.016309, 5.036768, 5.058268, 5.080154, 5.101726, 
    5.122242,
  // momentumY(14,49, 0-49)
    5.131782, 5.121768, 5.107812, 5.090503, 5.070491, 5.048445, 5.025044, 
    5.000954, 4.976798, 4.953141, 4.93047, 4.909184, 4.889575, 4.87183, 
    4.856054, 4.844022, 4.848143, 4.838534, 4.83033, 4.824347, 4.820787, 
    4.825149, 4.832235, 4.842608, 4.852149, 4.861037, 4.868387, 4.874065, 
    4.877024, 4.881012, 4.885324, 4.894529, 4.902976, 4.910685, 4.917894, 
    4.925021, 4.93263, 4.941376, 4.951897, 4.964715, 4.980152, 4.99826, 
    5.018826, 5.04138, 5.065258, 5.08966, 5.113735, 5.1366, 5.15739, 5.175267,
  // momentumY(15,0, 0-49)
    5.116331, 5.087602, 5.057508, 5.02688, 4.99647, 4.966957, 4.938937, 
    4.912934, 4.889373, 4.86856, 4.850661, 4.835689, 4.823497, 4.813806, 
    4.806232, 4.800476, 4.797285, 4.793497, 4.79044, 4.787902, 4.785748, 
    4.784293, 4.783263, 4.78291, 4.783345, 4.784853, 4.787655, 4.791958, 
    4.797826, 4.805394, 4.814459, 4.825126, 4.83667, 4.848646, 4.860583, 
    4.872067, 4.882796, 4.892663, 4.901782, 4.910505, 4.919398, 4.929152, 
    4.940503, 4.954107, 4.970463, 4.989839, 5.012252, 5.037459, 5.064975, 
    5.094105,
  // momentumY(15,1, 0-49)
    5.096625, 5.067094, 5.036662, 5.006133, 4.976219, 4.94755, 4.920673, 
    4.896048, 4.874031, 4.854852, 4.838602, 4.825209, 4.81445, 4.805967, 
    4.799304, 4.794245, 4.792803, 4.788857, 4.785463, 4.782435, 4.779634, 
    4.777761, 4.776192, 4.775315, 4.77516, 4.776093, 4.778361, 4.782217, 
    4.787709, 4.795141, 4.804237, 4.815469, 4.827672, 4.840302, 4.852779, 
    4.864544, 4.87516, 4.884389, 4.892262, 4.899111, 4.905552, 4.912408, 
    4.920602, 4.931015, 4.944372, 4.961137, 4.981477, 5.005255, 5.032047, 
    5.061183,
  // momentumY(15,2, 0-49)
    5.078791, 5.048922, 5.018562, 4.988491, 4.95939, 4.931859, 4.906399, 
    4.883417, 4.863198, 4.845896, 4.831511, 4.819883, 4.810696, 4.803508, 
    4.797784, 4.793371, 4.793595, 4.789402, 4.78556, 4.781904, 4.778296, 
    4.775818, 4.773477, 4.771796, 4.770742, 4.770769, 4.772155, 4.775218, 
    4.780015, 4.787013, 4.795884, 4.807501, 4.820284, 4.833621, 4.846819, 
    4.859183, 4.870113, 4.879212, 4.886373, 4.891838, 4.89621, 4.900389, 
    4.905457, 4.912516, 4.922533, 4.936205, 4.953891, 4.975585, 5.000948, 
    5.029352,
  // momentumY(15,3, 0-49)
    5.06324, 5.033447, 5.003518, 4.974208, 4.946181, 4.920012, 4.896168, 
    4.875008, 4.856752, 4.841472, 4.829074, 4.819304, 4.811752, 4.805884, 
    4.801088, 4.797221, 4.798965, 4.794469, 4.790111, 4.78574, 4.781212, 
    4.777983, 4.774674, 4.771935, 4.769695, 4.768483, 4.768632, 4.770534, 
    4.774281, 4.780493, 4.788819, 4.800562, 4.81377, 4.827785, 4.841828, 
    4.855076, 4.866765, 4.876311, 4.883421, 4.888182, 4.891104, 4.893085, 
    4.895307, 4.899062, 4.905564, 4.915772, 4.93028, 4.949261, 4.972499, 
    4.999438,
  // momentumY(15,4, 0-49)
    5.050073, 5.020701, 4.9915, 4.963202, 4.936454, 4.911811, 4.889717, 
    4.87048, 4.854262, 4.841056, 4.830678, 4.822776, 4.81685, 4.812282, 
    4.808378, 4.804924, 4.807982, 4.803201, 4.798327, 4.79323, 4.787751, 
    4.783697, 4.779289, 4.77529, 4.771614, 4.768863, 4.767426, 4.767785, 
    4.770104, 4.775139, 4.782532, 4.794057, 4.807438, 4.822003, 4.836916, 
    4.851248, 4.864085, 4.874649, 4.88243, 4.887299, 4.88959, 4.890103, 
    4.890029, 4.890785, 4.89381, 4.900341, 4.911246, 4.92694, 4.947388, 
    4.972149,
  // momentumY(15,5, 0-49)
    5.039103, 5.010417, 4.982175, 4.95508, 4.929761, 4.906757, 4.886483, 
    4.869208, 4.855032, 4.843874, 4.835467, 4.829376, 4.825019, 4.821709, 
    4.818674, 4.815492, 4.819603, 4.814657, 4.809369, 4.803624, 4.797256, 
    4.792387, 4.786834, 4.781446, 4.776152, 4.771607, 4.768267, 4.766716, 
    4.767217, 4.770647, 4.77667, 4.787555, 4.800759, 4.81563, 4.831312, 
    4.846801, 4.861059, 4.873127, 4.882268, 4.888099, 4.8907, 4.89067, 
    4.889099, 4.887434, 4.887277, 4.890124, 4.89716, 4.909099, 4.926156, 
    4.948071,
  // momentumY(15,6, 0-49)
    5.029912, 5.00209, 4.974963, 4.949202, 4.925413, 4.904112, 4.885684, 
    4.870354, 4.85817, 4.848981, 4.84245, 4.838074, 4.835212, 4.833121, 
    4.830979, 4.827941, 4.832795, 4.827935, 4.822438, 4.816226, 4.809129, 
    4.803551, 4.796894, 4.790074, 4.783056, 4.776528, 4.771018, 4.767218, 
    4.765527, 4.766914, 4.771096, 4.780854, 4.793445, 4.80827, 4.824483, 
    4.841054, 4.856845, 4.870752, 4.88182, 4.889394, 4.893252, 4.893704, 
    4.891622, 4.888361, 4.885583, 4.885003, 4.888118, 4.895999, 4.909183, 
    4.927671,
  // momentumY(15,7, 0-49)
    5.021935, 4.99507, 4.96914, 4.944782, 4.922575, 4.902999, 4.886406, 
    4.872977, 4.862704, 4.855379, 4.850611, 4.847847, 4.846417, 4.845552, 
    4.844402, 4.841412, 4.846661, 4.84226, 4.836864, 4.83046, 4.822882, 
    4.816778, 4.809143, 4.800937, 4.792175, 4.783555, 4.775673, 4.769339, 
    4.765112, 4.764037, 4.765896, 4.774005, 4.785484, 4.799817, 4.816212, 
    4.833632, 4.850895, 4.866778, 4.880141, 4.89007, 4.896023, 4.897958, 
    4.896429, 4.892569, 4.887981, 4.884502, 4.88391, 4.887653, 4.896658, 
    4.911267,
  // momentumY(15,8, 0-49)
    5.014567, 4.988669, 4.963949, 4.941008, 4.920386, 4.902526, 4.887734, 
    4.876143, 4.867693, 4.862128, 4.859016, 4.857789, 4.857767, 4.858192, 
    4.858227, 4.855232, 4.860509, 4.857036, 4.852131, 4.845875, 4.838133, 
    4.83175, 4.82334, 4.813871, 4.803432, 4.792694, 4.782328, 4.773249, 
    4.766201, 4.762278, 4.76136, 4.767284, 4.777114, 4.790453, 4.806582, 
    4.824496, 4.842996, 4.860787, 4.876583, 4.889243, 4.897914, 4.902189, 
    4.902226, 4.898835, 4.893422, 4.887823, 4.884019, 4.883815, 4.888562, 
    4.899018,
  // momentumY(15,9, 0-49)
    5.007263, 4.982272, 4.958714, 4.937149, 4.918076, 4.901892, 4.888849, 
    4.879029, 4.872319, 4.868426, 4.866897, 4.867163, 4.868573, 4.870416, 
    4.871912, 4.868925, 4.873866, 4.87183, 4.867853, 4.862131, 4.854586, 
    4.848204, 4.83927, 4.828737, 4.816766, 4.803984, 4.791113, 4.779171, 
    4.76909, 4.762001, 4.7579, 4.761126, 4.768773, 4.780583, 4.795938, 
    4.813896, 4.833264, 4.85271, 4.870847, 4.886352, 4.898101, 4.905329, 
    4.907785, 4.905872, 4.900687, 4.893928, 4.887661, 4.883976, 4.884649, 
    4.890883,
  // momentumY(15,10, 0-49)
    4.999604, 4.975416, 4.952922, 4.932649, 4.915052, 4.900475, 4.889113, 
    4.880991, 4.875949, 4.873662, 4.873672, 4.875424, 4.878328, 4.881759, 
    4.885052, 4.882169, 4.886457, 4.886337, 4.883721, 4.878932, 4.87196, 
    4.865866, 4.856699, 4.845355, 4.832079, 4.817416, 4.802129, 4.787311, 
    4.774088, 4.7636, 4.755988, 4.756044, 4.760993, 4.770745, 4.784802, 
    4.802295, 4.822069, 4.84278, 4.862974, 4.881195, 4.896103, 4.906617, 
    4.912094, 4.912504, 4.908549, 4.901665, 4.893864, 4.887411, 4.884446, 
    4.886625,
  // momentumY(15,11, 0-49)
    4.991342, 4.967822, 4.946262, 4.927166, 4.910937, 4.897869, 4.8881, 
    4.881597, 4.878156, 4.877424, 4.878942, 4.882198, 4.886673, 4.891865, 
    4.897288, 4.89474, 4.898158, 4.900331, 4.899464, 4.895978, 4.889944, 
    4.88441, 4.875308, 4.863452, 4.849164, 4.832879, 4.815373, 4.797784, 
    4.781417, 4.767402, 4.756055, 4.752538, 4.754327, 4.761522, 4.773763, 
    4.790272, 4.809944, 4.831436, 4.853266, 4.873887, 4.891792, 4.905651, 
    4.914472, 4.917807, 4.915928, 4.909914, 4.901585, 4.893248, 4.8873, 
    4.885808,
  // momentumY(15,12, 0-49)
    4.982402, 4.959404, 4.938636, 4.920569, 4.905574, 4.893891, 4.885602, 
    4.880623, 4.878705, 4.879471, 4.882472, 4.887239, 4.893341, 4.900425, 
    4.908225, 4.906451, 4.908953, 4.913633, 4.914804, 4.91294, 4.908176, 
    4.903432, 4.894686, 4.88264, 4.867683, 4.850114, 4.830691, 4.810552, 
    4.791155, 4.773605, 4.758424, 4.751015, 4.749251, 4.753448, 4.763399, 
    4.778428, 4.797483, 4.819242, 4.842208, 4.86478, 4.885344, 4.90237, 
    4.914593, 4.92119, 4.922007, 4.917713, 4.90983, 4.900563, 4.892437, 
    4.887838,
  // momentumY(15,13, 0-49)
    4.972854, 4.950241, 4.930109, 4.912913, 4.898992, 4.888544, 4.881598, 
    4.87802, 4.877524, 4.879713, 4.884143, 4.890391, 4.89812, 4.907125, 
    4.917382, 4.917123, 4.918903, 4.926107, 4.929477, 4.929471, 4.926257, 
    4.922477, 4.914348, 4.90243, 4.887171, 4.868714, 4.847758, 4.825398, 
    4.803198, 4.782228, 4.763248, 4.751732, 4.746114, 4.746946, 4.7542, 
    4.767303, 4.785262, 4.806781, 4.830365, 4.854382, 4.877144, 4.897, 
    4.912463, 4.922406, 4.926286, 4.924352, 4.917756, 4.908478, 4.899033, 
    4.892014,
  // momentumY(15,14, 0-49)
    4.96287, 4.940514, 4.920871, 4.904384, 4.891365, 4.881975, 4.876204, 
    4.873875, 4.874665, 4.878159, 4.883919, 4.89156, 4.900823, 4.911641, 
    4.924194, 4.926576, 4.928138, 4.937673, 4.943261, 4.945259, 4.943804, 
    4.941094, 4.933791, 4.922291, 4.907089, 4.888156, 4.866101, 4.841918, 
    4.817236, 4.793077, 4.770475, 4.754752, 4.745088, 4.742292, 4.746523, 
    4.757329, 4.773777, 4.7946, 4.818307, 4.843254, 4.867715, 4.889956, 
    4.908341, 4.921505, 4.928574, 4.929399, 4.924733, 4.916243, 4.906309, 
    4.897605,
  // momentumY(15,15, 0-49)
    4.952686, 4.930484, 4.911194, 4.895252, 4.88295, 4.874424, 4.869629, 
    4.868354, 4.870248, 4.874878, 4.881808, 4.890677, 4.901279, 4.913642, 
    4.92807, 4.93463, 4.936832, 4.948342, 4.95604, 4.960089, 4.960528, 
    4.958922, 4.952585, 4.941731, 4.926888, 4.907864, 4.885134, 4.85956, 
    4.832775, 4.80575, 4.779841, 4.759933, 4.746149, 4.739574, 4.740567, 
    4.748801, 4.763408, 4.783151, 4.806544, 4.831944, 4.857608, 4.881755, 
    4.90265, 4.918758, 4.928937, 4.932689, 4.930367, 4.923283, 4.913586, 
    4.903914,
  // momentumY(15,16, 0-49)
    4.942564, 4.920435, 4.90138, 4.885822, 4.874048, 4.866168, 4.862118, 
    4.86166, 4.864422, 4.869958, 4.877826, 4.887679, 4.899335, 4.912846, 
    4.92854, 4.941131, 4.945195, 4.958213, 4.967833, 4.973904, 4.976303, 
    4.975766, 4.970457, 4.960384, 4.946107, 4.927279, 4.904236, 4.877665, 
    4.849168, 4.819665, 4.790876, 4.766929, 4.749082, 4.738706, 4.736363, 
    4.741861, 4.7544, 4.77277, 4.795497, 4.820938, 4.847348, 4.872924, 
    4.89588, 4.91456, 4.92762, 4.934264, 4.934485, 4.929224, 4.920336, 
    4.910336,
  // momentumY(15,17, 0-49)
    4.932777, 4.910663, 4.891735, 4.876411, 4.864961, 4.857486, 4.853906, 
    4.853971, 4.857299, 4.863437, 4.871946, 4.88248, 4.894852, 4.909085, 
    4.925418, 4.945959, 4.953385, 4.967457, 4.978798, 4.986842, 4.991218, 
    4.991667, 4.987359, 4.978087, 4.964433, 4.945938, 4.922795, 4.895525, 
    4.865663, 4.834091, 4.80294, 4.77522, 4.753508, 4.739446, 4.733802, 
    4.736515, 4.746866, 4.76367, 4.785466, 4.810616, 4.837379, 4.863954, 
    4.888523, 4.909357, 4.924963, 4.934315, 4.937086, 4.933866, 4.926193, 
    4.916392,
  // momentumY(15,18, 0-49)
    4.923589, 4.901454, 4.882562, 4.867312, 4.855964, 4.848607, 4.845161, 
    4.845378, 4.848886, 4.855247, 4.864042, 4.874938, 4.887739, 4.902402, 
    4.918972, 4.949069, 4.961415, 4.976269, 4.989225, 4.999232, 5.005604, 
    5.006928, 5.003522, 4.994929, 4.981759, 4.963496, 4.940249, 4.9124, 
    4.881422, 4.848179, 4.815248, 4.784146, 4.758912, 4.741425, 4.732646, 
    4.732654, 4.740804, 4.755947, 4.776639, 4.801248, 4.828047, 4.855239, 
    4.881002, 4.903563, 4.921335, 4.933104, 4.938289, 4.93716, 4.930946, 
    4.921741,
  // momentumY(15,19, 0-49)
    4.915263, 4.893085, 4.874133, 4.858778, 4.847258, 4.839663, 4.83592, 
    4.835809, 4.838999, 4.845114, 4.853805, 4.864809, 4.877959, 4.89312, 
    4.910018, 4.950513, 4.968981, 4.984726, 4.999439, 5.011564, 5.02004, 
    5.022157, 5.019508, 5.011316, 4.998226, 4.979774, 4.956087, 4.927523, 
    4.895533, 4.860983, 4.826902, 4.792949, 4.764691, 4.744195, 4.732588, 
    4.730083, 4.736119, 4.749599, 4.769093, 4.792991, 4.819576, 4.847066, 
    4.873648, 4.897533, 4.917068, 4.93091, 4.938273, 4.939157, 4.934505, 
    4.926172,
  // momentumY(15,20, 0-49)
    4.908185, 4.886056, 4.867468, 4.852916, 4.84274, 4.837077, 4.835821, 
    4.838592, 4.844738, 4.853366, 4.863411, 4.873747, 4.883327, 4.89133, 
    4.897302, 0, 4.994577, 4.999668, 5.005548, 5.011305, 5.016126, 5.015633, 
    5.013115, 5.006968, 4.997258, 4.982792, 4.962961, 4.937488, 4.907465, 
    4.873701, 4.839848, 4.803802, 4.772908, 4.749545, 4.735105, 4.72999, 
    4.733762, 4.745383, 4.763453, 4.786373, 4.812434, 4.839869, 4.866875, 
    4.891658, 4.912527, 4.928051, 4.937283, 4.939999, 4.936891, 4.929584,
  // momentumY(15,21, 0-49)
    4.90235, 4.880386, 4.861916, 4.847402, 4.837146, 4.831253, 4.829581, 
    4.831733, 4.837054, 4.844685, 4.853627, 4.862837, 4.871323, 4.878238, 
    4.882979, 0, 5.004196, 5.009486, 5.015777, 5.021951, 5.027033, 5.024549, 
    5.020569, 5.013208, 5.002763, 4.988084, 4.968498, 4.943565, 4.914167, 
    4.880956, 4.847917, 4.810899, 4.778774, 4.753971, 4.737977, 4.73131, 
    4.733636, 4.743992, 4.761029, 4.783178, 4.80876, 4.836029, 4.863201, 
    4.888492, 4.910194, 4.926821, 4.937312, 4.941274, 4.939192, 4.932497,
  // momentumY(15,22, 0-49)
    4.897773, 4.875886, 4.857458, 4.842922, 4.832562, 4.826463, 4.824469, 
    4.826171, 4.830924, 4.837883, 4.846084, 4.854511, 4.862186, 4.868207, 
    4.871812, 0, 5.010537, 5.015932, 5.022656, 5.029411, 5.035066, 5.0311, 
    5.026239, 5.01824, 5.007516, 4.992895, 4.973616, 4.949099, 4.920087, 
    4.887161, 4.854692, 4.816629, 4.78334, 4.757275, 4.739974, 4.732033, 
    4.73318, 4.742507, 4.758702, 4.78022, 4.805398, 4.83251, 4.859784, 
    4.885447, 4.907785, 4.925273, 4.936773, 4.941762, 4.940569, 4.934464,
  // momentumY(15,23, 0-49)
    4.894632, 4.872791, 4.854372, 4.839801, 4.829348, 4.823086, 4.820855, 
    4.822244, 4.826617, 4.833141, 4.840868, 4.848798, 4.855937, 4.861334, 
    4.864092, 0, 5.014832, 5.020237, 5.02725, 5.034447, 5.040577, 5.035399, 
    5.029847, 5.021343, 5.010375, 4.995757, 4.976672, 4.952449, 4.923741, 
    4.891075, 4.859142, 4.82031, 4.786209, 4.75929, 4.741114, 4.732311, 
    4.73266, 4.741292, 4.75692, 4.778018, 4.802937, 4.829955, 4.857316, 
    4.883248, 4.906034, 4.924124, 4.93632, 4.94202, 4.941433, 4.935718,
  // momentumY(15,24, 0-49)
    4.89303, 4.871227, 4.852822, 4.83823, 4.827715, 4.821345, 4.818963, 
    4.820161, 4.824309, 4.830588, 4.838061, 4.845731, 4.8526, 4.857682, 4.86, 
    0, 5.017446, 5.022851, 5.03004, 5.037525, 5.043984, 5.038036, 5.032043, 
    5.023195, 5.012022, 4.997339, 4.978312, 4.954233, 4.925709, 4.893244, 
    4.861749, 4.822506, 4.787988, 4.760626, 4.741983, 4.732702, 4.732585, 
    4.740788, 4.756044, 4.776845, 4.801548, 4.828448, 4.855792, 4.881816, 
    4.904807, 4.9232, 4.935774, 4.941876, 4.941653, 4.936192,
  // momentumY(15,25, 0-49)
    4.892978, 4.871228, 4.852853, 4.838268, 4.827735, 4.821324, 4.818879, 
    4.820003, 4.824073, 4.830282, 4.8377, 4.84534, 4.852205, 4.857303, 
    4.859646, 0, 5.017977, 5.023447, 5.030755, 5.038391, 5.045011, 5.03886, 
    5.032743, 5.023767, 5.012475, 4.997696, 4.978612, 4.954521, 4.926036, 
    4.893661, 4.862384, 4.823091, 4.788538, 4.761134, 4.742421, 4.733041, 
    4.732802, 4.74087, 4.755989, 4.776659, 4.801252, 4.828063, 4.855346, 
    4.881342, 4.904335, 4.922764, 4.935397, 4.941571, 4.941417, 4.935998,
  // momentumY(15,26, 0-49)
    4.894406, 4.87272, 4.854392, 4.839842, 4.829338, 4.822953, 4.820543, 
    4.82172, 4.82587, 4.832198, 4.839781, 4.84764, 4.854785, 4.860251, 
    4.863098, 0, 5.016332, 5.021949, 5.029336, 5.036996, 5.043603, 5.037862, 
    5.031976, 5.023129, 5.011848, 4.996982, 4.977752, 4.953513, 4.924929, 
    4.892527, 4.861219, 4.822248, 4.78804, 4.760976, 4.742573, 4.733451, 
    4.733408, 4.741605, 4.756795, 4.777483, 4.802044, 4.828778, 4.855942, 
    4.881776, 4.904565, 4.922753, 4.935126, 4.941044, 4.940664, 4.935086,
  // momentumY(15,27, 0-49)
    4.89715, 4.875522, 4.857244, 4.842745, 4.83231, 4.826026, 4.823761, 
    4.825141, 4.829566, 4.836245, 4.84426, 4.852632, 4.860379, 4.866575, 
    4.870389, 0, 5.012642, 5.018445, 5.025831, 5.033369, 5.039788, 5.035005, 
    5.029674, 5.021203, 5.01006, 4.995123, 4.97568, 4.951184, 4.922391, 
    4.889878, 4.858337, 4.820057, 4.786572, 4.760231, 4.74251, 4.733994, 
    4.734449, 4.743031, 4.758483, 4.779317, 4.80391, 4.830564, 4.857533, 
    4.883053, 4.905414, 4.923075, 4.934859, 4.940183, 4.939286, 4.933345,
  // momentumY(15,28, 0-49)
    4.900956, 4.87935, 4.861095, 4.846647, 4.83631, 4.830202, 4.828211, 
    4.829986, 4.834939, 4.842281, 4.851081, 4.860333, 4.869051, 4.876345, 
    4.881514, 0, 5.007342, 5.013274, 5.020514, 5.02774, 5.033801, 5.030379, 
    5.02587, 5.017995, 5.00712, 4.992149, 4.972463, 4.947652, 4.918607, 
    4.885978, 4.854132, 4.816909, 4.784528, 4.759285, 4.742601, 4.735004, 
    4.736219, 4.745374, 4.761208, 4.782232, 4.806831, 4.833304, 4.85991, 
    4.884882, 4.906523, 4.923325, 4.934174, 4.938588, 4.936932, 4.93051,
  // momentumY(15,29, 0-49)
    4.905488, 4.883822, 4.865526, 4.851095, 4.840873, 4.835017, 4.833459, 
    4.83588, 4.841707, 4.850139, 4.860193, 4.870795, 4.8809, 4.889626, 
    4.896388, 0, 5.000063, 5.005975, 5.012874, 5.019604, 5.025175, 5.023331, 
    5.019852, 5.012797, 5.002379, 4.987502, 4.967638, 4.942543, 4.913272, 
    4.880569, 4.848407, 4.812506, 4.781537, 4.757733, 4.742431, 4.736076, 
    4.738331, 4.748291, 4.764679, 4.786003, 4.810646, 4.836909, 4.86304, 
    4.887277, 4.907935, 4.923557, 4.933121, 4.936285, 4.933587, 4.926498,
  // momentumY(15,30, 0-49)
    4.910488, 4.888827, 4.870213, 4.855021, 4.843503, 4.83578, 4.831827, 
    4.831496, 4.834548, 4.840704, 4.849711, 4.861379, 4.875586, 4.892223, 
    4.911034, 4.954827, 4.973868, 4.991736, 5.008694, 5.022947, 5.033298, 
    5.035358, 5.033057, 5.025144, 5.012241, 4.993824, 4.97003, 4.941264, 
    4.909084, 4.874454, 4.840883, 4.805935, 4.77645, 4.754404, 4.74091, 
    4.73623, 4.739908, 4.750978, 4.768137, 4.789886, 4.814612, 4.84061, 
    4.866129, 4.889415, 4.908816, 4.922949, 4.930926, 4.932596, 4.928713, 
    4.920949,
  // momentumY(15,31, 0-49)
    4.915942, 4.89447, 4.876083, 4.861194, 4.850078, 4.842865, 4.83952, 
    4.839871, 4.843635, 4.850474, 4.860056, 4.872119, 4.886497, 4.903143, 
    4.922074, 4.95497, 4.968733, 4.986028, 5.00144, 5.013679, 5.021948, 
    5.023351, 5.020294, 5.011942, 4.998954, 4.980783, 4.957542, 4.929637, 
    4.898599, 4.865321, 4.832775, 4.800514, 4.773793, 4.754419, 4.743352, 
    4.740744, 4.746068, 4.758324, 4.776205, 4.798216, 4.822738, 4.848071, 
    4.872464, 4.894181, 4.911629, 4.923537, 4.929198, 4.928702, 4.923073, 
    4.914211,
  // momentumY(15,32, 0-49)
    4.921215, 4.899942, 4.881758, 4.8671, 4.856259, 4.849372, 4.846404, 
    4.847165, 4.851349, 4.858582, 4.868499, 4.880802, 4.895323, 4.912056, 
    4.93118, 4.954336, 4.96384, 4.98057, 4.994486, 5.004793, 5.011045, 
    5.011725, 5.007792, 4.99875, 4.985291, 4.966941, 4.943911, 4.916705, 
    4.886889, 4.855299, 4.824359, 4.795338, 4.771907, 4.755643, 4.747331, 
    4.746997, 4.754054, 4.767476, 4.785954, 4.808, 4.832004, 4.856267, 
    4.879059, 4.898688, 4.913652, 4.922843, 4.925797, 4.9229, 4.91548, 
    4.905674,
  // momentumY(15,33, 0-49)
    4.92593, 4.904881, 4.886914, 4.872478, 4.861875, 4.855245, 4.852547, 
    4.853583, 4.858017, 4.865453, 4.875493, 4.887812, 4.902227, 4.91875, 
    4.937635, 4.952839, 4.959489, 4.975294, 4.98753, 4.995835, 5.000043, 
    4.999904, 4.99502, 4.985198, 4.971148, 4.952522, 4.929667, 4.903242, 
    4.874849, 4.845289, 4.816482, 4.7911, 4.771321, 4.758461, 4.753111, 
    4.755168, 4.763979, 4.778497, 4.797407, 4.819228, 4.842355, 4.865105, 
    4.885779, 4.902761, 4.914688, 4.920676, 4.920567, 4.915102, 4.905936, 
    4.895429,
  // momentumY(15,34, 0-49)
    4.929762, 4.908973, 4.891263, 4.877086, 4.866748, 4.860384, 4.857946, 
    4.859209, 4.863815, 4.871333, 4.881327, 4.893431, 4.907422, 4.923276, 
    4.941233, 4.950496, 4.955647, 4.969988, 4.980257, 4.986433, 4.988561, 
    4.987503, 4.981656, 4.971096, 4.956528, 4.937751, 4.915259, 4.889861, 
    4.86318, 4.836005, 4.809812, 4.788346, 4.772446, 4.763155, 4.760866, 
    4.765345, 4.775867, 4.791358, 4.810493, 4.831789, 4.853648, 4.874407, 
    4.892422, 4.906191, 4.914549, 4.916904, 4.913468, 4.905375, 4.89462, 
    4.883753,
  // momentumY(15,35, 0-49)
    4.932462, 4.911976, 4.894581, 4.880731, 4.870724, 4.864684, 4.862538, 
    4.864038, 4.868792, 4.87632, 4.886137, 4.897826, 4.911088, 4.925822, 
    4.942156, 4.947344, 4.952077, 4.964399, 4.972419, 4.976362, 4.976421, 
    4.974379, 4.967628, 4.95648, 4.941605, 4.922957, 4.901151, 4.877123, 
    4.852477, 4.828023, 4.80485, 4.787461, 4.77554, 4.769867, 4.77063, 
    4.777473, 4.789596, 4.805881, 4.824989, 4.845424, 4.865595, 4.883875, 
    4.898703, 4.908737, 4.913075, 4.911485, 4.904602, 4.893983, 4.881938, 
    4.87114,
  // momentumY(15,36, 0-49)
    4.933903, 4.91376, 4.896746, 4.883297, 4.873699, 4.86805, 4.866251, 
    4.868015, 4.872907, 4.880397, 4.889943, 4.901053, 4.91335, 4.926611, 
    4.940794, 4.943399, 4.948446, 4.958294, 4.963863, 4.965548, 4.963623, 
    4.960588, 4.953065, 4.941565, 4.926686, 4.908533, 4.887803, 4.865521, 
    4.843225, 4.821772, 4.801928, 4.788659, 4.780696, 4.778567, 4.782275, 
    4.791337, 4.804873, 4.821717, 4.840497, 4.85971, 4.87777, 4.893103, 
    4.904272, 4.910153, 4.91017, 4.904511, 4.894277, 4.881431, 4.868542, 
    4.858325,
  // momentumY(15,37, 0-49)
    4.934103, 4.914344, 4.897767, 4.884783, 4.875652, 4.870442, 4.86902, 
    4.871055, 4.876065, 4.883467, 4.892656, 4.903069, 4.914239, 4.925816, 
    4.937567, 4.938635, 4.944391, 4.951484, 4.954533, 4.954038, 4.950295, 
    4.946325, 4.938226, 4.926672, 4.912144, 4.894886, 4.875633, 4.855452, 
    4.83577, 4.817514, 4.801187, 4.791965, 4.787823, 4.789057, 4.795502, 
    4.806548, 4.821237, 4.838345, 4.856464, 4.874076, 4.889618, 4.9016, 
    4.908755, 4.910237, 4.905857, 4.896271, 4.883037, 4.868485, 4.855347, 
    4.846265,
  // momentumY(15,38, 0-49)
    4.933275, 4.913924, 4.897812, 4.885321, 4.876671, 4.871897, 4.870824, 
    4.873085, 4.878146, 4.88538, 4.894122, 4.903744, 4.913695, 4.923514, 
    4.932799, 4.932977, 4.93955, 4.943816, 4.944435, 4.941947, 4.936632, 
    4.93186, 4.923436, 4.912159, 4.898354, 4.882379, 4.864967, 4.847182, 
    4.8303, 4.815341, 4.802587, 4.797229, 4.79666, 4.800972, 4.809848, 
    4.822561, 4.83807, 4.855095, 4.872189, 4.887829, 4.900504, 4.908844, 
    4.911808, 4.908888, 4.900332, 4.88727, 4.871682, 4.85616, 4.843473, 
    4.836088,
  // momentumY(15,39, 0-49)
    4.931844, 4.912904, 4.897245, 4.885211, 4.876986, 4.87256, 4.871725, 
    4.874079, 4.879056, 4.885987, 4.894164, 4.902904, 4.911595, 4.919686, 
    4.926654, 4.926291, 4.933585, 4.935168, 4.933599, 4.929408, 4.922832, 
    4.91746, 4.909001, 4.898345, 4.885618, 4.871275, 4.856004, 4.840826, 
    4.826837, 4.815162, 4.805911, 4.804132, 4.80679, 4.813807, 4.824722, 
    4.838705, 4.85464, 4.871191, 4.88689, 4.900232, 4.909787, 4.914362, 
    4.913201, 4.906186, 4.894016, 4.878262, 4.861233, 4.845648, 4.834178, 
    4.828999,
  // momentumY(15,40, 0-49)
    4.930457, 4.911899, 4.896629, 4.884946, 4.876993, 4.872725, 4.87191, 
    4.874125, 4.878788, 4.885204, 4.892647, 4.900396, 4.907799, 4.914251, 
    4.919162, 4.918425, 4.926207, 4.925446, 4.92205, 4.916519, 4.909047, 
    4.903338, 4.895158, 4.885455, 4.874131, 4.861706, 4.848792, 4.836337, 
    4.825235, 4.816731, 4.810798, 4.812224, 4.817683, 4.826947, 4.839435, 
    4.854232, 4.870153, 4.885829, 4.899788, 4.910583, 4.91692, 4.917839, 
    4.912915, 4.902449, 4.887573, 4.870214, 4.852869, 4.838229, 4.828725, 
    4.826172,
  // momentumY(15,41, 0-49)
    4.929952, 4.911724, 4.896721, 4.885202, 4.877274, 4.872872, 4.871749, 
    4.873485, 4.877499, 4.883104, 4.889571, 4.896175, 4.902244, 4.907153, 
    4.910297, 4.909247, 4.917224, 4.914587, 4.909807, 4.903347, 4.895372, 
    4.889627, 4.882048, 4.873604, 4.863957, 4.853662, 4.843232, 4.833522, 
    4.825214, 4.819678, 4.816773, 4.820962, 4.828731, 4.839725, 4.853273, 
    4.868386, 4.883842, 4.898261, 4.910213, 4.918354, 4.921581, 4.919222, 
    4.911222, 4.898285, 4.881907, 4.864242, 4.847815, 4.835123, 4.828254, 
    4.828617,
  // momentumY(15,42, 0-49)
    4.931294, 4.913325, 4.898424, 4.886817, 4.878589, 4.873669, 4.871818, 
    4.872636, 4.875574, 4.879983, 4.885159, 4.890398, 4.895037, 4.898464, 
    4.900094, 4.898733, 4.906603, 4.902615, 4.896917, 4.88995, 4.881868, 
    4.876405, 4.86973, 4.862811, 4.855051, 4.847018, 4.839118, 4.832088, 
    4.826405, 4.823557, 4.823317, 4.829775, 4.83932, 4.851501, 4.865571, 
    4.880503, 4.89507, 4.907923, 4.917725, 4.923294, 4.923772, 4.918811, 
    4.908726, 4.894571, 4.878089, 4.861507, 4.847205, 4.837363, 4.833653, 
    4.837076,
  // momentumY(15,43, 0-49)
    4.935475, 4.917697, 4.902711, 4.890727, 4.881828, 4.875952, 4.872892, 
    4.872292, 4.873665, 4.876423, 4.879921, 4.883506, 4.886554, 4.888489, 
    4.888772, 4.887052, 4.894532, 4.889695, 4.883519, 4.876438, 4.868618, 
    4.863738, 4.85823, 4.853035, 4.847303, 4.841592, 4.836183, 4.831695, 
    4.828406, 4.827918, 4.829926, 4.83814, 4.84892, 4.86174, 4.875812, 
    4.89011, 4.90344, 4.914546, 4.922236, 4.925542, 4.923896, 4.917282, 
    4.906342, 4.892384, 4.877251, 4.863077, 4.851962, 4.845681, 4.845468, 
    4.851949,
  // momentumY(15,44, 0-49)
    4.943389, 4.925753, 4.910508, 4.897867, 4.887924, 4.880651, 4.875891, 
    4.873359, 4.872651, 4.87327, 4.874662, 4.876251, 4.877479, 4.87783, 
    4.876827, 4.87465, 4.881481, 4.876204, 4.869909, 4.863044, 4.855793, 
    4.851745, 4.847598, 4.844251, 4.840609, 4.837198, 4.834173, 4.832032, 
    4.830871, 4.832383, 4.836201, 4.845671, 4.857166, 4.870117, 4.883736, 
    4.897036, 4.908914, 4.918256, 4.924076, 4.925666, 4.922758, 4.91564, 
    4.905199, 4.892863, 4.880429, 4.869793, 4.862683, 4.860432, 4.863861, 
    4.873267,
  // momentumY(15,45, 0-49)
    4.955724, 4.938224, 4.922591, 4.909056, 4.897744, 4.88868, 4.881776, 
    4.876834, 4.873561, 4.871572, 4.870428, 4.86966, 4.868797, 4.867399, 
    4.865062, 4.862271, 4.868221, 4.862769, 4.856599, 4.850181, 4.843715, 
    4.840663, 4.837982, 4.836504, 4.834927, 4.833717, 4.832911, 4.832884, 
    4.833569, 4.836724, 4.841933, 4.852195, 4.863946, 4.876606, 4.889421, 
    4.901495, 4.911865, 4.919618, 4.924015, 4.924632, 4.921483, 4.915091, 
    4.906478, 4.897058, 4.888436, 4.882178, 4.879595, 4.881592, 4.888622, 
    4.900716,
  // momentumY(15,46, 0-49)
    4.972857, 4.955551, 4.939471, 4.924886, 4.911969, 4.900812, 4.891409, 
    4.883674, 4.877432, 4.872438, 4.868383, 4.864922, 4.861692, 4.858339, 
    4.854538, 4.850924, 4.855777, 4.850251, 4.844319, 4.838459, 4.832879, 
    4.830882, 4.82966, 4.82997, 4.830338, 4.831164, 4.832362, 4.834197, 
    4.836456, 4.840928, 4.847151, 4.857822, 4.869471, 4.881536, 4.893338, 
    4.904113, 4.913095, 4.919608, 4.923187, 4.923685, 4.921351, 4.916856, 
    4.911235, 4.905757, 4.901744, 4.900376, 4.902549, 4.908782, 4.91922, 
    4.933684,
  // momentumY(15,47, 0-49)
    4.994822, 4.977833, 4.961337, 4.945648, 4.931002, 4.917567, 4.905441, 
    4.894656, 4.885172, 4.87689, 4.869647, 4.863233, 4.857401, 4.851891, 
    4.846448, 4.841775, 4.845335, 4.839686, 4.833971, 4.828657, 4.82394, 
    4.822939, 4.823054, 4.824963, 4.827073, 4.829704, 4.832666, 4.836111, 
    4.839708, 4.845225, 4.85217, 4.862968, 4.874279, 4.885587, 4.896322, 
    4.905891, 4.913754, 4.9195, 4.922939, 4.92417, 4.923613, 4.921988, 
    4.920238, 4.919398, 4.920445, 4.924166, 4.931067, 4.941337, 4.954875, 
    4.971336,
  // momentumY(15,48, 0-49)
    5.021287, 5.004817, 4.988027, 4.971284, 4.954903, 4.939142, 4.92421, 
    4.910266, 4.897417, 4.885714, 4.875143, 4.865629, 4.857044, 4.849217, 
    4.841962, 4.835991, 4.838085, 4.832155, 4.826528, 4.821638, 4.817649, 
    4.817477, 4.818703, 4.821928, 4.825503, 4.829668, 4.834137, 4.838961, 
    4.843709, 4.850078, 4.857544, 4.868315, 4.879192, 4.88973, 4.899494, 
    4.908081, 4.915195, 4.920693, 4.92464, 4.927336, 4.929301, 4.931226, 
    4.933884, 4.938024, 4.944261, 4.953, 4.964405, 4.978386, 4.994637, 5.01268,
  // momentumY(15,49, 0-49)
    5.058356, 5.043217, 5.026606, 5.00895, 4.990648, 4.972076, 4.953585, 
    4.935503, 4.918123, 4.901687, 4.886375, 4.872292, 4.859453, 4.847805, 
    4.837231, 4.829314, 4.83676, 4.82897, 4.82178, 4.815975, 4.811789, 
    4.814678, 4.819662, 4.827548, 4.834721, 4.8415, 4.847211, 4.851875, 
    4.854626, 4.859023, 4.86429, 4.875, 4.885332, 4.89494, 4.903584, 
    4.911133, 4.917612, 4.923219, 4.928326, 4.933444, 4.939155, 4.946041, 
    4.9546, 4.965176, 4.977912, 4.992743, 5.009426, 5.027546, 5.046576, 
    5.065892,
  // momentumY(16,0, 0-49)
    5.010379, 4.983305, 4.957535, 4.933589, 4.911873, 4.89267, 4.876139, 
    4.862313, 4.851107, 4.842322, 4.835676, 4.830809, 4.827321, 4.824801, 
    4.82285, 4.821224, 4.82087, 4.8188, 4.816489, 4.813863, 4.810887, 
    4.80795, 4.804797, 4.801712, 4.798837, 4.796524, 4.795112, 4.794984, 
    4.796442, 4.799865, 4.805302, 4.813079, 4.822648, 4.833603, 4.845372, 
    4.857257, 4.868512, 4.878438, 4.88649, 4.892384, 4.896164, 4.898243, 
    4.899375, 4.90057, 4.90296, 4.907646, 4.915551, 4.92732, 4.943265, 
    4.963357,
  // momentumY(16,1, 0-49)
    4.998121, 4.971027, 4.945522, 4.922115, 4.901196, 4.88303, 4.86775, 
    4.855347, 4.845687, 4.838506, 4.833449, 4.830081, 4.827929, 4.826505, 
    4.825345, 4.824247, 4.825438, 4.823134, 4.820419, 4.817234, 4.813533, 
    4.810053, 4.806176, 4.802295, 4.798471, 4.795121, 4.792607, 4.79137, 
    4.791726, 4.794225, 4.798886, 4.806432, 4.81596, 4.827044, 4.839068, 
    4.851271, 4.86282, 4.87292, 4.880921, 4.886435, 4.889426, 4.890259, 
    4.889693, 4.888795, 4.888814, 4.891007, 4.896475, 4.906033, 4.920139, 
    4.938877,
  // momentumY(16,2, 0-49)
    4.988944, 4.96211, 4.937086, 4.914367, 4.894336, 4.877245, 4.863204, 
    4.852176, 4.84398, 4.838302, 4.834718, 4.832727, 4.831792, 4.831364, 
    4.830914, 4.830249, 4.832897, 4.830378, 4.827298, 4.8236, 4.819216, 
    4.815224, 4.810616, 4.805884, 4.801012, 4.796468, 4.792636, 4.790017, 
    4.788951, 4.790158, 4.793639, 4.800545, 4.809657, 4.82056, 4.832631, 
    4.845079, 4.857021, 4.867584, 4.876018, 4.881814, 4.884809, 4.885249, 
    4.883801, 4.88151, 4.879666, 4.879637, 4.882692, 4.889841, 4.901728, 
    4.918592,
  // momentumY(16,3, 0-49)
    4.98254, 4.95621, 4.931844, 4.90993, 4.890845, 4.874831, 4.861982, 
    4.852237, 4.845376, 4.841043, 4.838762, 4.837986, 4.838121, 4.838571, 
    4.838752, 4.838411, 4.842396, 4.83975, 4.836403, 4.832302, 4.827349, 
    4.822939, 4.817657, 4.812073, 4.806106, 4.800255, 4.794926, 4.790676, 
    4.787887, 4.787426, 4.789301, 4.795124, 4.80339, 4.813739, 4.82558, 
    4.838131, 4.850492, 4.86174, 4.871041, 4.877756, 4.88156, 4.882516, 
    4.881122, 4.878296, 4.87528, 4.873495, 4.874341, 4.879025, 4.888411, 
    4.902944,
  // momentumY(16,4, 0-49)
    4.978348, 4.952726, 4.929165, 4.908149, 4.890049, 4.875096, 4.863371, 
    4.854793, 4.849114, 4.845946, 4.844783, 4.845037, 4.846092, 4.847313, 
    4.848078, 4.847959, 4.853121, 4.85051, 4.847063, 4.842731, 4.837382, 
    4.832712, 4.826875, 4.8205, 4.813451, 4.806242, 4.799288, 4.793202, 
    4.788418, 4.785934, 4.785778, 4.790048, 4.797011, 4.806389, 4.817661, 
    4.830092, 4.842803, 4.854854, 4.865345, 4.873514, 4.878854, 4.881207, 
    4.880831, 4.878424, 4.875085, 4.872192, 4.871225, 4.873564, 4.880309, 
    4.89215,
  // momentumY(16,5, 0-49)
    4.975636, 4.950883, 4.928251, 4.908212, 4.891126, 4.877218, 4.866553, 
    4.859032, 4.85439, 4.852214, 4.851986, 4.853107, 4.85495, 4.856871, 
    4.858217, 4.858232, 4.864367, 4.862026, 4.858702, 4.854363, 4.848849, 
    4.844121, 4.837903, 4.830859, 4.822809, 4.814256, 4.805618, 4.797554, 
    4.790562, 4.785738, 4.78315, 4.785407, 4.790595, 4.798553, 4.808867, 
    4.820886, 4.833784, 4.84663, 4.858483, 4.868478, 4.87593, 4.880437, 
    4.881971, 4.880943, 4.878209, 4.875005, 4.872805, 4.87311, 4.877246, 
    4.886169,
  // momentumY(16,6, 0-49)
    4.97359, 4.949832, 4.92823, 4.909238, 4.893208, 4.880342, 4.870695, 
    4.864148, 4.860424, 4.859102, 4.859666, 4.861528, 4.864074, 4.866668, 
    4.868656, 4.868736, 4.875587, 4.873809, 4.870874, 4.866787, 4.861371, 
    4.856816, 4.85043, 4.842885, 4.83398, 4.824172, 4.81387, 4.803766, 
    4.794423, 4.787009, 4.781643, 4.781456, 4.784411, 4.790498, 4.799439, 
    4.810699, 4.823528, 4.837036, 4.850263, 4.862264, 4.872192, 4.87941, 
    4.883584, 4.884794, 4.883579, 4.880935, 4.878224, 4.876989, 4.878732, 
    4.884682,
  // momentumY(16,7, 0-49)
    4.971429, 4.948754, 4.928265, 4.910394, 4.895467, 4.883669, 4.87503, 
    4.869415, 4.866539, 4.865985, 4.867253, 4.869784, 4.872997, 4.876294, 
    4.879041, 4.879138, 4.8864, 4.885508, 4.883248, 4.879677, 4.874628, 
    4.870487, 4.864169, 4.856335, 4.846771, 4.835867, 4.824009, 4.811897, 
    4.800161, 4.789993, 4.781582, 4.778574, 4.778876, 4.782658, 4.789808, 
    4.799926, 4.812365, 4.826291, 4.840752, 4.85474, 4.86728, 4.877518, 
    4.884831, 4.888952, 4.890053, 4.888813, 4.886382, 4.88424, 4.883992, 
    4.887099,
  // momentumY(16,8, 0-49)
    4.9685, 4.946961, 4.927648, 4.910966, 4.897206, 4.886523, 4.878919, 
    4.874241, 4.872197, 4.872381, 4.874321, 4.877502, 4.881399, 4.885472, 
    4.889145, 4.889234, 4.896564, 4.896873, 4.895561, 4.892765, 4.888341, 
    4.884839, 4.878826, 4.870933, 4.860958, 4.849187, 4.835968, 4.82198, 
    4.807916, 4.794942, 4.783319, 4.777194, 4.774482, 4.775564, 4.780519, 
    4.789104, 4.800787, 4.814806, 4.83023, 4.846014, 4.861082, 4.874398, 
    4.885083, 4.892534, 4.896551, 4.897444, 4.896061, 4.893718, 4.892021, 
    4.892599,
  // momentumY(16,9, 0-49)
    4.964339, 4.943954, 4.92586, 4.910425, 4.897897, 4.888393, 4.88188, 
    4.878181, 4.876997, 4.87794, 4.88057, 4.88443, 4.889064, 4.894015, 
    4.898808, 4.898908, 4.90595, 4.907724, 4.907599, 4.905803, 4.90224, 
    4.89956, 4.894073, 4.886361, 4.876246, 4.863895, 4.849592, 4.833972, 
    4.817759, 4.802047, 4.787168, 4.777723, 4.771718, 4.769764, 4.772158, 
    4.778826, 4.789371, 4.803106, 4.81913, 4.836383, 4.853708, 4.869932, 
    4.883956, 4.894887, 4.902172, 4.905732, 4.906059, 4.904214, 4.901698, 
    4.900219,
  // momentumY(16,10, 0-49)
    4.958708, 4.939458, 4.922597, 4.908445, 4.897206, 4.888947, 4.88359, 
    4.880938, 4.880676, 4.882433, 4.885808, 4.890401, 4.895841, 4.901774, 
    4.907865, 4.908079, 4.914513, 4.917924, 4.919169, 4.918551, 4.916037, 
    4.914315, 4.909543, 4.902239, 4.892272, 4.879665, 4.864626, 4.847709, 
    4.829641, 4.811388, 4.793344, 4.780487, 4.770998, 4.76575, 4.765265, 
    4.769666, 4.77869, 4.791737, 4.807944, 4.826241, 4.845419, 4.864198, 
    4.881311, 4.895623, 4.906263, 4.912791, 4.915321, 4.914591, 4.911907, 
    4.908954,
  // momentumY(16,11, 0-49)
    4.951579, 4.933411, 4.917763, 4.904904, 4.894985, 4.88802, 4.883884, 
    4.882345, 4.883079, 4.88572, 4.889904, 4.895293, 4.901602, 4.9086, 
    4.916114, 4.916668, 4.922263, 4.927371, 4.930091, 4.930777, 4.929453, 
    4.928766, 4.924852, 4.918157, 4.908612, 4.89609, 4.88071, 4.862903, 
    4.84337, 4.822893, 4.801913, 4.785665, 4.77261, 4.763888, 4.760275, 
    4.762101, 4.769247, 4.781209, 4.797158, 4.816027, 4.836568, 4.857426, 
    4.877209, 4.894594, 4.908454, 4.918019, 4.923042, 4.923909, 4.92166, 
    4.917865,
  // momentumY(16,12, 0-49)
    4.94311, 4.925941, 4.911447, 4.899851, 4.89125, 4.885598, 4.882725, 
    4.882352, 4.884141, 4.887729, 4.892781, 4.899015, 4.906228, 4.914317, 
    4.923285, 4.924597, 4.929274, 4.936002, 4.940219, 4.942276, 4.942241, 
    4.942596, 4.939634, 4.933708, 4.924829, 4.912722, 4.897404, 4.879156, 
    4.858614, 4.836325, 4.812768, 4.793261, 4.776662, 4.764382, 4.757468, 
    4.756468, 4.761423, 4.771923, 4.787184, 4.80614, 4.827521, 4.849919, 
    4.871853, 4.891866, 4.908628, 4.921103, 4.928713, 4.931497, 4.930191, 
    4.926173,
  // momentumY(16,13, 0-49)
    4.933587, 4.917305, 4.903876, 4.893475, 4.886146, 4.881787, 4.880175, 
    4.88099, 4.883869, 4.888443, 4.894396, 4.901491, 4.909599, 4.918728, 
    4.929043, 4.931781, 4.935657, 4.943816, 4.94947, 4.952912, 4.954217, 
    4.955572, 4.953596, 4.948547, 4.940525, 4.92912, 4.914241, 4.895998, 
    4.874925, 4.8513, 4.825628, 4.803096, 4.783074, 4.767251, 4.756944, 
    4.752938, 4.755445, 4.764153, 4.778327, 4.796912, 4.81862, 4.842006, 
    4.865535, 4.887653, 4.906889, 4.921998, 4.932122, 4.936985, 4.937004, 
    4.933322,
  // momentumY(16,14, 0-49)
    4.923371, 4.90785, 4.895366, 4.886055, 4.879909, 4.876776, 4.87638, 
    4.87836, 4.882319, 4.887879, 4.894729, 4.902659, 4.9116, 4.921633, 
    4.933037, 4.938135, 4.941565, 4.95087, 4.957839, 4.962636, 4.965298, 
    4.967563, 4.966561, 4.962437, 4.955395, 4.944908, 4.93078, 4.912937, 
    4.891786, 4.867318, 4.84006, 4.814806, 4.791577, 4.772316, 4.758617, 
    4.751506, 4.751376, 4.758027, 4.770776, 4.788579, 4.810141, 4.833998, 
    4.858574, 4.882263, 4.903494, 4.920869, 4.933316, 4.940278, 4.941876, 
    4.938986,
  // momentumY(16,15, 0-49)
    4.912854, 4.897959, 4.88628, 4.877921, 4.87283, 4.870809, 4.871537, 
    4.874606, 4.87959, 4.886088, 4.893784, 4.90248, 4.912133, 4.922858, 
    4.93496, 4.94358, 4.947157, 4.957278, 4.965407, 4.971506, 4.97552, 
    4.978578, 4.978491, 4.975286, 4.969269, 4.959824, 4.946657, 4.929514, 
    4.908661, 4.883808, 4.855515, 4.827887, 4.801735, 4.779232, 4.762231, 
    4.752002, 4.749129, 4.753531, 4.764589, 4.781275, 4.80229, 4.826159, 
    4.851291, 4.876046, 4.898795, 4.918036, 4.932535, 4.941511, 4.944815, 
    4.943059,
  // momentumY(16,16, 0-49)
    4.902413, 4.888007, 4.876982, 4.869414, 4.865215, 4.864151, 4.865855, 
    4.869885, 4.87578, 4.883116, 4.891562, 4.900916, 4.911123, 4.922285, 
    4.934649, 4.948032, 4.952551, 4.96318, 4.972324, 4.979673, 4.985033, 
    4.98876, 4.989505, 4.98716, 4.982129, 4.973736, 4.961613, 4.945337, 
    4.92504, 4.900175, 4.871372, 4.841729, 4.81299, 4.787511, 4.767387, 
    4.75412, 4.748487, 4.750541, 4.759723, 4.775039, 4.795194, 4.818704, 
    4.843974, 4.86935, 4.893178, 4.913892, 4.930142, 4.940972, 4.946005, 
    4.945608,
  // momentumY(16,17, 0-49)
    4.892386, 4.878341, 4.867813, 4.860855, 4.857354, 4.857041, 4.859523, 
    4.864323, 4.870955, 4.878976, 4.88804, 4.897923, 4.908541, 4.919922, 
    4.932185, 4.951418, 4.957764, 4.968699, 4.978784, 4.987378, 4.994099, 
    4.998383, 4.999869, 4.998282, 4.994113, 4.986661, 4.975505, 4.960099, 
    4.940459, 4.915834, 4.886974, 4.855661, 4.824695, 4.796576, 4.773589, 
    4.757456, 4.749144, 4.748833, 4.756054, 4.769843, 4.78891, 4.811782, 
    4.836864, 4.862501, 4.88703, 4.908854, 4.926551, 4.939031, 4.945736, 
    4.946805,
  // momentumY(16,18, 0-49)
    4.883057, 4.86925, 4.859056, 4.852509, 4.849472, 4.849656, 4.852646, 
    4.857956, 4.865088, 4.873597, 4.88313, 4.893447, 4.904416, 4.91596, 
    4.927983, 4.95368, 4.962641, 4.973895, 4.984979, 4.994907, 5.003065, 
    5.007842, 5.009997, 5.009035, 5.005515, 4.998745, 4.988299, 4.973565, 
    4.954499, 4.930216, 4.901648, 4.868981, 4.836173, 4.805798, 4.780288, 
    4.761552, 4.750729, 4.748141, 4.753402, 4.76559, 4.783442, 4.805486, 
    4.83014, 4.855759, 4.880685, 4.903311, 4.922166, 4.936076, 4.944336, 
    4.946891,
  // momentumY(16,19, 0-49)
    4.874649, 4.860956, 4.850918, 4.844546, 4.841686, 4.842038, 4.845186, 
    4.850657, 4.857982, 4.866745, 4.876626, 4.887396, 4.898871, 4.910821, 
    4.922827, 4.954803, 4.966801, 4.978681, 4.991045, 5.002561, 5.012359, 
    5.017647, 5.020454, 5.019977, 5.016799, 5.010279, 5.000051, 4.985547, 
    4.966752, 4.942739, 4.9147, 4.880971, 4.846727, 4.814543, 4.786932, 
    4.765944, 4.752872, 4.748176, 4.751559, 4.76216, 4.778742, 4.799853, 
    4.823924, 4.849325, 4.874414, 4.897583, 4.917346, 4.932465, 4.942127, 
    4.946119,
  // momentumY(16,20, 0-49)
    4.867816, 4.854584, 4.845321, 4.840126, 4.838893, 4.841312, 4.846864, 
    4.85486, 4.864492, 4.874896, 4.885221, 4.894706, 4.902756, 4.909014, 
    4.913389, 0, 4.987489, 4.991956, 4.99765, 5.003873, 5.010102, 5.012218, 
    5.01397, 5.014071, 5.012827, 5.009157, 5.002196, 4.990902, 4.974914, 
    4.953116, 4.927007, 4.893116, 4.858006, 4.824359, 4.79484, 4.771689, 
    4.756392, 4.749557, 4.751001, 4.759923, 4.775121, 4.79516, 4.818483, 
    4.843477, 4.868512, 4.891992, 4.912422, 4.928527, 4.93941, 4.944731,
  // momentumY(16,21, 0-49)
    4.861976, 4.848943, 4.839874, 4.834837, 4.833697, 4.836112, 4.841539, 
    4.849289, 4.858567, 4.868547, 4.878441, 4.887538, 4.895265, 4.901219, 
    4.905196, 0, 4.992397, 4.997305, 5.003582, 5.010384, 5.017054, 5.017688, 
    5.018337, 5.017498, 5.015707, 5.011953, 5.005382, 4.994881, 4.979984, 
    4.959462, 4.935041, 4.90137, 4.866254, 4.832252, 4.801982, 4.777731, 
    4.761089, 4.752796, 4.752783, 4.760341, 4.774326, 4.793342, 4.815856, 
    4.840277, 4.864996, 4.888429, 4.909086, 4.925674, 4.937243, 4.943362,
  // momentumY(16,22, 0-49)
    4.857375, 4.844437, 4.83546, 4.830493, 4.82939, 4.83179, 4.837147, 
    4.844765, 4.853857, 4.863614, 4.873266, 4.882125, 4.889603, 4.895244, 
    4.898731, 0, 4.995681, 5.000916, 5.007755, 5.015225, 5.022527, 5.022017, 
    5.021948, 5.020552, 5.018504, 5.014805, 5.008574, 4.99863, 4.984444, 
    4.964725, 4.941484, 4.907679, 4.872356, 4.837974, 4.807092, 4.781999, 
    4.764341, 4.754937, 4.753801, 4.760295, 4.773324, 4.791523, 4.813382, 
    4.837328, 4.86177, 4.885137, 4.905946, 4.922899, 4.935011, 4.941789,
  // momentumY(16,23, 0-49)
    4.854089, 4.841188, 4.83224, 4.82729, 4.82618, 4.828554, 4.833859, 
    4.841405, 4.850407, 4.860065, 4.869614, 4.878358, 4.885695, 4.891115, 
    4.894202, 0, 4.998227, 5.003655, 5.010888, 5.018858, 5.026659, 5.025187, 
    5.024527, 5.02266, 5.020362, 5.016635, 5.010581, 5.000975, 4.98724, 
    4.968055, 4.945672, 4.911668, 4.876164, 4.841541, 4.810292, 4.784687, 
    4.76639, 4.756265, 4.754383, 4.760154, 4.772521, 4.790148, 4.811541, 
    4.835138, 4.85936, 4.882646, 4.903519, 4.920674, 4.933112, 4.940302,
  // momentumY(16,24, 0-49)
    4.852131, 4.839238, 4.830288, 4.825319, 4.824179, 4.826513, 4.831777, 
    4.839285, 4.848259, 4.8579, 4.867444, 4.876188, 4.88351, 4.888863, 
    4.891764, 0, 5.000336, 5.005877, 5.013352, 5.021645, 5.029784, 5.027698, 
    5.026659, 5.024476, 5.021976, 5.018165, 5.01214, 5.002656, 4.989122, 
    4.970199, 4.948319, 4.914134, 4.878489, 4.843718, 4.812261, 4.786366, 
    4.767694, 4.757131, 4.754774, 4.760069, 4.771986, 4.789208, 4.810258, 
    4.833585, 4.857615, 4.880801, 4.901666, 4.918907, 4.931514, 4.938937,
  // momentumY(16,25, 0-49)
    4.85146, 4.838564, 4.829591, 4.824589, 4.823408, 4.825703, 4.830941, 
    4.838443, 4.847441, 4.857141, 4.866776, 4.875635, 4.883084, 4.888557, 
    4.891555, 0, 5.001617, 5.00724, 5.014842, 5.023288, 5.03158, 5.02933, 
    5.02819, 5.025898, 5.02329, 5.019381, 5.01327, 5.003716, 4.990139, 
    4.971201, 4.949409, 4.915092, 4.87936, 4.844524, 4.813005, 4.787022, 
    4.768224, 4.757499, 4.754951, 4.760036, 4.771738, 4.788752, 4.809611, 
    4.83277, 4.856662, 4.879742, 4.900535, 4.917737, 4.930336, 4.937777,
  // momentumY(16,26, 0-49)
    4.851977, 4.839075, 4.830077, 4.825035, 4.82382, 4.826095, 4.831341, 
    4.838893, 4.847992, 4.857843, 4.867679, 4.876782, 4.884514, 4.890315, 
    4.893711, 0, 5.001983, 5.007671, 5.015292, 5.023718, 5.031972, 5.030043, 
    5.029104, 5.026941, 5.024355, 5.020361, 5.014077, 5.004286, 4.990434, 
    4.971213, 4.949087, 4.914718, 4.878968, 4.844158, 4.812709, 4.786823, 
    4.768129, 4.757494, 4.755009, 4.760123, 4.771822, 4.788801, 4.809599, 
    4.832676, 4.856466, 4.87942, 4.900066, 4.917099, 4.929512, 4.936756,
  // momentumY(16,27, 0-49)
    4.853549, 4.84063, 4.831599, 4.826528, 4.825302, 4.827601, 4.832926, 
    4.840624, 4.849943, 4.860089, 4.870278, 4.879788, 4.887972, 4.894296, 
    4.898354, 0, 5.001553, 5.007257, 5.014753, 5.022965, 5.030978, 5.02979, 
    5.029314, 5.027491, 5.025039, 5.020969, 5.014422, 5.00423, 4.989888, 
    4.970133, 4.947292, 4.912957, 4.877278, 4.842611, 4.811395, 4.785818, 
    4.767478, 4.757198, 4.755036, 4.760416, 4.772312, 4.789418, 4.810269, 
    4.833325, 4.857021, 4.879806, 4.900201, 4.916908, 4.928932, 4.935752,
  // momentumY(16,28, 0-49)
    4.855995, 4.843037, 4.833967, 4.828879, 4.827681, 4.830082, 4.835604, 
    4.843608, 4.853339, 4.863991, 4.874754, 4.884873, 4.89369, 4.900697, 
    4.905574, 0, 5.000744, 5.006339, 5.013515, 5.021286, 5.028846, 5.028683, 
    5.02886, 5.027533, 5.025298, 5.021149, 5.014251, 5.003506, 4.988485, 
    4.967993, 4.944139, 4.909925, 4.874425, 4.840048, 4.809262, 4.78423, 
    4.766501, 4.756835, 4.75523, 4.761073, 4.773315, 4.790642, 4.811593, 
    4.834626, 4.858176, 4.88069, 4.900694, 4.916894, 4.928325, 4.934512,
  // momentumY(16,29, 0-49)
    4.859104, 4.846059, 4.836926, 4.831833, 4.830725, 4.833347, 4.839246, 
    4.847798, 4.858232, 4.869702, 4.881335, 4.892307, 4.901924, 4.909692, 
    4.91538, 0, 4.999225, 5.004516, 5.011139, 5.018236, 5.025145, 5.026101, 
    5.027013, 5.026284, 5.024335, 5.02012, 5.012819, 5.001411, 4.985559, 
    4.964156, 4.939056, 4.904996, 4.869781, 4.835892, 4.805812, 4.781667, 
    4.764914, 4.756218, 4.755496, 4.762076, 4.774881, 4.792583, 4.813718, 
    4.836743, 4.86009, 4.882205, 4.90162, 4.917064, 4.927612, 4.93287,
  // momentumY(16,30, 0-49)
    4.862476, 4.849107, 4.839384, 4.833349, 4.830894, 4.831782, 4.835658, 
    4.842111, 4.850717, 4.861089, 4.872904, 4.885905, 4.899866, 4.914509, 
    4.92938, 4.966947, 4.978901, 4.992922, 5.007429, 5.020907, 5.032383, 
    5.037577, 5.040587, 5.040208, 5.037008, 5.03027, 5.019615, 5.004519, 
    4.98509, 4.960538, 4.932539, 4.897691, 4.862357, 4.828973, 4.799906, 
    4.777106, 4.761838, 4.754601, 4.75519, 4.762854, 4.776481, 4.794729, 
    4.81613, 4.839152, 4.862225, 4.883802, 4.902434, 4.91689, 4.926324, 
    4.930448,
  // momentumY(16,31, 0-49)
    4.866781, 4.853611, 4.844128, 4.83839, 4.836299, 4.837609, 4.84195, 
    4.848881, 4.857934, 4.868675, 4.880737, 4.893844, 4.9078, 4.922468, 
    4.937697, 4.967824, 4.977847, 4.991458, 5.004806, 5.016727, 5.02653, 
    5.031267, 5.033574, 5.032618, 5.028995, 5.021968, 5.011114, 4.995862, 
    4.976276, 4.951561, 4.923069, 4.889333, 4.855425, 4.823767, 4.796635, 
    4.775844, 4.762507, 4.756995, 4.759011, 4.767756, 4.782095, 4.800686, 
    4.822061, 4.844687, 4.867003, 4.887477, 4.904691, 4.917486, 4.925124, 
    4.927476,
  // momentumY(16,32, 0-49)
    4.871303, 4.858335, 4.849073, 4.843582, 4.841766, 4.843366, 4.848002, 
    4.855215, 4.864517, 4.875458, 4.887661, 4.900854, 4.91489, 4.929732, 
    4.945438, 4.968321, 4.976445, 4.989829, 5.002178, 5.012691, 5.02094, 
    5.025236, 5.026824, 5.025161, 5.020825, 5.013091, 5.001563, 4.985727, 
    4.965698, 4.940761, 4.912001, 4.879725, 4.847709, 4.81828, 4.793566, 
    4.775197, 4.764112, 4.760547, 4.764117, 4.773983, 4.788996, 4.807811, 
    4.82897, 4.850946, 4.872193, 4.891208, 4.906636, 4.917415, 4.922964, 
    4.92335,
  // momentumY(16,33, 0-49)
    4.875925, 4.863193, 4.854173, 4.84893, 4.847354, 4.84918, 4.854009, 
    4.861369, 4.870765, 4.881741, 4.893917, 4.907042, 4.921004, 4.935845, 
    4.951768, 4.968263, 4.974986, 4.988035, 4.999339, 5.008449, 5.015163, 
    5.01895, 5.019767, 5.017297, 5.012066, 5.003394, 4.99095, 4.974339, 
    4.95378, 4.928711, 4.900013, 4.869541, 4.839824, 4.813044, 4.791133, 
    4.775503, 4.766909, 4.765444, 4.770644, 4.78163, 4.797239, 4.816132, 
    4.836852, 4.857888, 4.877718, 4.894889, 4.908136, 4.916543, 4.919724, 
    4.917984,
  // momentumY(16,34, 0-49)
    4.880545, 4.868095, 4.859358, 4.854384, 4.85305, 4.855068, 4.860024, 
    4.867435, 4.876794, 4.887642, 4.899608, 4.912449, 4.926073, 4.940565, 
    4.956202, 4.967526, 4.973517, 4.985917, 4.996002, 5.003626, 5.008771, 
    5.011938, 5.011914, 5.00858, 5.002374, 4.992685, 4.979272, 4.961896, 
    4.940898, 4.915932, 4.887727, 4.859404, 4.832354, 4.80857, 4.789754, 
    4.777088, 4.771133, 4.771847, 4.778687, 4.790736, 4.806821, 4.825599, 
    4.845624, 4.865399, 4.883441, 4.89837, 4.909048, 4.914743, 4.915324, 
    4.911375,
  // momentumY(16,35, 0-49)
    4.885081, 4.87296, 4.864542, 4.85986, 4.858766, 4.86095, 4.865981, 
    4.873355, 4.882562, 4.893137, 4.904713, 4.917045, 4.930042, 4.943787, 
    4.95856, 4.96601, 4.971895, 4.98324, 4.991876, 4.997907, 5.001445, 
    5.003863, 5.002946, 4.998738, 4.991569, 4.980916, 4.966636, 4.948666, 
    4.927465, 4.902946, 4.87573, 4.849896, 4.825834, 4.805314, 4.78979, 
    4.780211, 4.776949, 4.779835, 4.788252, 4.801247, 4.817632, 4.836062, 
    4.855099, 4.87327, 4.889144, 4.901443, 4.909194, 4.911911, 4.909752, 
    4.903614,
  // momentumY(16,36, 0-49)
    4.889462, 4.877706, 4.869629, 4.86524, 4.864367, 4.866679, 4.871722, 
    4.878978, 4.887927, 4.898099, 4.909123, 4.920747, 4.932858, 4.9455, 
    4.958887, 4.963627, 4.969875, 4.979753, 4.986724, 4.99107, 4.992982, 
    4.994537, 4.992704, 4.987673, 4.979637, 4.968187, 4.95327, 4.935, 
    4.913944, 4.890288, 4.86458, 4.841549, 4.820729, 4.803648, 4.791512, 
    4.78504, 4.784429, 4.789392, 4.799244, 4.812998, 4.82945, 4.847256, 
    4.864984, 4.881196, 4.894536, 4.903861, 4.908413, 4.907989, 4.90308, 
    4.894912,
  // momentumY(16,37, 0-49)
    4.893633, 4.882252, 4.874506, 4.870379, 4.869679, 4.872052, 4.877029, 
    4.88408, 4.892673, 4.902333, 4.912676, 4.923434, 4.934464, 4.94574, 
    4.957366, 4.960308, 4.967186, 4.975255, 4.980393, 4.983005, 4.983312, 
    4.983918, 4.981193, 4.975446, 4.966719, 4.954725, 4.939501, 4.921314, 
    4.900814, 4.878473, 4.854766, 4.834799, 4.817393, 4.803834, 4.79508, 
    4.791636, 4.793539, 4.800397, 4.811465, 4.825723, 4.841955, 4.858814, 
    4.87489, 4.888796, 4.899277, 4.905368, 4.906568, 4.902996, 4.895502, 
    4.885627,
  // momentumY(16,38, 0-49)
    4.897552, 4.886523, 4.879058, 4.875122, 4.874506, 4.876844, 4.881657, 
    4.888404, 4.896548, 4.905604, 4.915175, 4.924968, 4.934794, 4.944555, 
    4.954224, 4.956, 4.963574, 4.969604, 4.972828, 4.973719, 4.972487, 
    4.972108, 4.968562, 4.962262, 4.953082, 4.940866, 4.925722, 4.908052, 
    4.888546, 4.867952, 4.846678, 4.82996, 4.816054, 4.805999, 4.800521, 
    4.799932, 4.804125, 4.812616, 4.824606, 4.83905, 4.854722, 4.870285, 
    4.884364, 4.895648, 4.903024, 4.905744, 4.903603, 4.897072, 4.887355, 
    4.876265,
  // momentumY(16,39, 0-49)
    4.901218, 4.89047, 4.88319, 4.879328, 4.878665, 4.880836, 4.885359, 
    4.891698, 4.899304, 4.907685, 4.916423, 4.925197, 4.933774, 4.94198, 
    4.94967, 4.950666, 4.958837, 4.962734, 4.964062, 4.96331, 4.960653, 
    4.959311, 4.955066, 4.948422, 4.939073, 4.926993, 4.912344, 4.89563, 
    4.877538, 4.859074, 4.840569, 4.827199, 4.81678, 4.810116, 4.807721, 
    4.809731, 4.815915, 4.825707, 4.838266, 4.852526, 4.867264, 4.881167, 
    4.892925, 4.901339, 4.905478, 4.904854, 4.89959, 4.890512, 4.879136, 
    4.86748,
  // momentumY(16,40, 0-49)
    4.904684, 4.894101, 4.886861, 4.882905, 4.882024, 4.883858, 4.887946, 
    4.893749, 4.900727, 4.90837, 4.916239, 4.923985, 4.931323, 4.938021, 
    4.943837, 4.94427, 4.952819, 4.954637, 4.954183, 4.951932, 4.948014, 
    4.94579, 4.941018, 4.934273, 4.925064, 4.913489, 4.89974, 4.884389, 
    4.868077, 4.852043, 4.83653, 4.826512, 4.819475, 4.816006, 4.816424, 
    4.820711, 4.828525, 4.839235, 4.851963, 4.865639, 4.879057, 4.89096, 
    4.900132, 4.905531, 4.906458, 4.902721, 4.89478, 4.883789, 4.871507, 
    4.860053,
  // momentumY(16,41, 0-49)
    4.908092, 4.897519, 4.89013, 4.885876, 4.884562, 4.88586, 4.889328, 
    4.894451, 4.90069, 4.907524, 4.914495, 4.921216, 4.927366, 4.932658, 
    4.93679, 4.93676, 4.945415, 4.945338, 4.943303, 4.939752, 4.934779, 
    4.93182, 4.926731, 4.920149, 4.911396, 4.900678, 4.888195, 4.874551, 
    4.86031, 4.846904, 4.834485, 4.827735, 4.823891, 4.823347, 4.826247, 
    4.832436, 4.841479, 4.852689, 4.86517, 4.87786, 4.889602, 4.899222, 
    4.905647, 4.908044, 4.905981, 4.899584, 4.889641, 4.877569, 4.865269, 
    4.854838,
  // momentumY(16,42, 0-49)
    4.911717, 4.900965, 4.893209, 4.888418, 4.886428, 4.886953, 4.889586, 
    4.893843, 4.899196, 4.905123, 4.911144, 4.91684, 4.921854, 4.925863, 
    4.928534, 4.928086, 4.936563, 4.934877, 4.931522, 4.926918, 4.92114, 
    4.917643, 4.912477, 4.906325, 4.89833, 4.888782, 4.877871, 4.866199, 
    4.854226, 4.843546, 4.834213, 4.830557, 4.829648, 4.831701, 4.836706, 
    4.84439, 4.854242, 4.865532, 4.877361, 4.888703, 4.898479, 4.905645, 
    4.909317, 4.908913, 4.904303, 4.895933, 4.88486, 4.872675, 4.861303, 
    4.852696,
  // momentumY(16,43, 0-49)
    4.915979, 4.904849, 4.896491, 4.890907, 4.887977, 4.887463, 4.889009, 
    4.892169, 4.896441, 4.901309, 4.90628, 4.910909, 4.914815, 4.91765, 
    4.919073, 4.918221, 4.926271, 4.923316, 4.918942, 4.91356, 4.907251, 
    4.903452, 4.898461, 4.892997, 4.886028, 4.877912, 4.868806, 4.859283, 
    4.849682, 4.841722, 4.835365, 4.834563, 4.836274, 4.840557, 4.847266, 
    4.856031, 4.866275, 4.877251, 4.888074, 4.897788, 4.905428, 4.910126, 
    4.911233, 4.908454, 4.901965, 4.892494, 4.881298, 4.870026, 4.860497, 
    4.854419,
  // momentumY(16,44, 0-49)
    4.921442, 4.909743, 4.900558, 4.893926, 4.889781, 4.887942, 4.888114, 
    4.889902, 4.892839, 4.89643, 4.900186, 4.903648, 4.906418, 4.90814, 
    4.908477, 4.907215, 4.914638, 4.910761, 4.905677, 4.899805, 4.89325, 
    4.8894, 4.884832, 4.880281, 4.874562, 4.868074, 4.860928, 4.853642, 
    4.846432, 4.841105, 4.837529, 4.839285, 4.843264, 4.849389, 4.857398, 
    4.866843, 4.877102, 4.887429, 4.896988, 4.90492, 4.910418, 4.912833, 
    4.911785, 4.907272, 4.89976, 4.890192, 4.879921, 4.87054, 4.863652, 
    4.860648,
  // momentumY(16,45, 0-49)
    4.928774, 4.916354, 4.906143, 4.89823, 4.892606, 4.889152, 4.887639, 
    4.887737, 4.889032, 4.891066, 4.893369, 4.895489, 4.897025, 4.897626, 
    4.89697, 4.895264, 4.901911, 4.897421, 4.891912, 4.885824, 4.879295, 
    4.875637, 4.871709, 4.868249, 4.863946, 4.85921, 4.854095, 4.849058, 
    4.844183, 4.84133, 4.840287, 4.844272, 4.850154, 4.857734, 4.866662, 
    4.876428, 4.886393, 4.895836, 4.903998, 4.910158, 4.913705, 4.914233, 
    4.911644, 4.906223, 4.898661, 4.890035, 4.881682, 4.875031, 4.871395, 
    4.871812,
  // momentumY(16,46, 0-49)
    4.93868, 4.925437, 4.914054, 4.904667, 4.897326, 4.891982, 4.888477, 
    4.886553, 4.885867, 4.886013, 4.886566, 4.887105, 4.88724, 4.886635, 
    4.884993, 4.88277, 4.888525, 4.883657, 4.877955, 4.871884, 4.865617, 
    4.862357, 4.859235, 4.856978, 4.854181, 4.851244, 4.848159, 4.845309, 
    4.842661, 4.842082, 4.843284, 4.849162, 4.856587, 4.865265, 4.874779, 
    4.88458, 4.894042, 4.902493, 4.909286, 4.913868, 4.915846, 4.915076, 
    4.911729, 4.906325, 4.899712, 4.892994, 4.887399, 4.884111, 4.884117, 
    4.888099,
  // momentumY(16,47, 0-49)
    4.951799, 4.937706, 4.925067, 4.914071, 4.904827, 4.897355, 4.891575, 
    4.887312, 4.884302, 4.88222, 4.880702, 4.879376, 4.87789, 4.875928, 
    4.873226, 4.870365, 4.875134, 4.870023, 4.864284, 4.858397, 4.852556, 
    4.849838, 4.847615, 4.846592, 4.845309, 4.844142, 4.843019, 4.842241, 
    4.841671, 4.843141, 4.846299, 4.853746, 4.862389, 4.871863, 4.881702, 
    4.891355, 4.900224, 4.907723, 4.913341, 4.916712, 4.917672, 4.916331, 
    4.913086, 4.908631, 4.903881, 4.899878, 4.897662, 4.89813, 4.901938, 
    4.909441,
  // momentumY(16,48, 0-49)
    4.968619, 4.953721, 4.939814, 4.927141, 4.915872, 4.906098, 4.897817, 
    4.890945, 4.885314, 4.880691, 4.876794, 4.873322, 4.869973, 4.866468, 
    4.862566, 4.858901, 4.862593, 4.857264, 4.85155, 4.845926, 4.840598, 
    4.838478, 4.837162, 4.837315, 4.837472, 4.837968, 4.838675, 4.839813, 
    4.841158, 4.844455, 4.849295, 4.858031, 4.867624, 4.877662, 4.887666, 
    4.897097, 4.905418, 4.912148, 4.916932, 4.919597, 4.920197, 4.91906, 
    4.916761, 4.914085, 4.911936, 4.911226, 4.912759, 4.917141, 4.92471, 
    4.935537,
  // momentumY(16,49, 0-49)
    4.997341, 4.981748, 4.96641, 4.95162, 4.937616, 4.924573, 4.9126, 
    4.901742, 4.89198, 4.883229, 4.875348, 4.868152, 4.861418, 4.854907, 
    4.848384, 4.843278, 4.852906, 4.845834, 4.83861, 4.832042, 4.8264, 
    4.827126, 4.82929, 4.833854, 4.837558, 4.840845, 4.843235, 4.844953, 
    4.845376, 4.847987, 4.852074, 4.862319, 4.872993, 4.88364, 4.893794, 
    4.902972, 4.910752, 4.916822, 4.921046, 4.923507, 4.924527, 4.92465, 
    4.9246, 4.925184, 4.927189, 4.931278, 4.93792, 4.947337, 4.959503, 
    4.974175,
  // momentumY(17,0, 0-49)
    4.932086, 4.910845, 4.892358, 4.876889, 4.864563, 4.855368, 4.849143, 
    4.845583, 4.844279, 4.84473, 4.846404, 4.84877, 4.851345, 4.853716, 
    4.855547, 4.85666, 4.858193, 4.857396, 4.855773, 4.853347, 4.850139, 
    4.846555, 4.84232, 4.837674, 4.832701, 4.827689, 4.822936, 4.818818, 
    4.815685, 4.813998, 4.813952, 4.81605, 4.819995, 4.825649, 4.832704, 
    4.840699, 4.849057, 4.857137, 4.864295, 4.869975, 4.873768, 4.8755, 
    4.875279, 4.87353, 4.870981, 4.868604, 4.867512, 4.868828, 4.873548, 
    4.882422,
  // momentumY(17,1, 0-49)
    4.927293, 4.906449, 4.888511, 4.873724, 4.862199, 4.853904, 4.848652, 
    4.846119, 4.845862, 4.847353, 4.850029, 4.853331, 4.856744, 4.859819, 
    4.862175, 4.863629, 4.866576, 4.865678, 4.863865, 4.861151, 4.857523, 
    4.853695, 4.849001, 4.843752, 4.837935, 4.831862, 4.825829, 4.820256, 
    4.815511, 4.812222, 4.810579, 4.811505, 4.814435, 4.819283, 4.825787, 
    4.83351, 4.841879, 4.850229, 4.85787, 4.864164, 4.868599, 4.870879, 
    4.870985, 4.869229, 4.866257, 4.863015, 4.860652, 4.860381, 4.863338, 
    4.87043,
  // momentumY(17,2, 0-49)
    4.925047, 4.904743, 4.887443, 4.873371, 4.862625, 4.855145, 4.85073, 
    4.849032, 4.849593, 4.851871, 4.855292, 4.859291, 4.863336, 4.866961, 
    4.86975, 4.871462, 4.875763, 4.874875, 4.873009, 4.870171, 4.866305, 
    4.862421, 4.857438, 4.851728, 4.845177, 4.838098, 4.830777, 4.823665, 
    4.817146, 4.812004, 4.80843, 4.807797, 4.809296, 4.812929, 4.81851, 
    4.825661, 4.833847, 4.842411, 4.850638, 4.857832, 4.863382, 4.866856, 
    4.868075, 4.867185, 4.864679, 4.861393, 4.858432, 4.857043, 4.85846, 
    4.863751,
  // momentumY(17,3, 0-49)
    4.924704, 4.905055, 4.888456, 4.875116, 4.865107, 4.858351, 4.854629, 
    4.85358, 4.85474, 4.85757, 4.861506, 4.865989, 4.870497, 4.874556, 
    4.877724, 4.879621, 4.88518, 4.884454, 4.882708, 4.879936, 4.876042, 
    4.872316, 4.867249, 4.861258, 4.854124, 4.846151, 4.837596, 4.828926, 
    4.820539, 4.813347, 4.807551, 4.805, 4.804668, 4.806671, 4.810932, 
    4.817171, 4.824917, 4.833555, 4.842372, 4.850632, 4.85764, 4.862832, 
    4.865854, 4.866643, 4.865483, 4.863023, 4.860238, 4.858329, 4.858582, 
    4.862187,
  // momentumY(17,4, 0-49)
    4.925554, 4.906652, 4.890803, 4.878195, 4.868879, 4.862763, 4.859605, 
    4.859044, 4.860619, 4.863809, 4.868073, 4.87288, 4.877728, 4.882148, 
    4.885689, 4.887709, 4.894379, 4.894003, 4.892564, 4.890065, 4.886366, 
    4.88302, 4.878093, 4.872019, 4.8645, 4.855797, 4.846127, 4.835956, 
    4.825689, 4.816328, 4.808094, 4.803315, 4.800786, 4.800761, 4.803308, 
    4.808267, 4.815266, 4.823757, 4.833058, 4.842415, 4.85107, 4.858335, 
    4.863684, 4.866829, 4.867804, 4.867007, 4.865207, 4.863475, 4.863067, 
    4.865251,
  // momentumY(17,5, 0-49)
    4.926895, 4.908814, 4.893754, 4.881882, 4.873228, 4.86768, 4.86499, 
    4.864796, 4.866652, 4.870066, 4.874532, 4.879558, 4.884674, 4.889433, 
    4.893384, 4.89547, 4.903042, 4.903224, 4.902287, 4.900254, 4.896966, 
    4.894212, 4.889642, 4.883701, 4.87602, 4.866802, 4.856206, 4.844675, 
    4.832611, 4.821059, 4.810258, 4.803021, 4.79799, 4.795586, 4.796041, 
    4.799346, 4.805257, 4.813318, 4.822897, 4.833249, 4.843571, 4.853073, 
    4.861067, 4.867047, 4.870778, 4.872372, 4.872322, 4.871489, 4.871013, 
    4.872166,
  // momentumY(17,6, 0-49)
    4.928093, 4.910898, 4.896666, 4.885541, 4.877535, 4.872518, 4.870237, 
    4.870338, 4.872396, 4.875957, 4.880558, 4.885754, 4.891115, 4.89623, 
    4.900664, 4.902766, 4.910966, 4.911911, 4.911652, 4.910261, 4.907574, 
    4.905591, 4.901582, 4.895983, 4.888383, 4.878903, 4.867634, 4.85497, 
    4.841294, 4.827643, 4.814258, 4.804423, 4.796666, 4.791592, 4.789618, 
    4.790914, 4.795382, 4.802684, 4.812258, 4.823384, 4.835237, 4.84695, 
    4.857692, 4.866757, 4.873649, 4.878177, 4.88052, 4.881258, 4.881336, 
    4.881945,
  // momentumY(17,7, 0-49)
    4.928635, 4.912382, 4.89902, 4.888669, 4.88132, 4.87683, 4.874942, 
    4.875315, 4.877554, 4.88124, 4.88596, 4.891318, 4.896939, 4.902454, 
    4.907468, 4.909537, 4.918041, 4.919922, 4.920493, 4.919884, 4.91795, 
    4.916876, 4.913595, 4.908529, 4.901253, 4.891789, 4.880151, 4.866659, 
    4.851659, 4.836112, 4.820251, 4.80779, 4.797184, 4.789228, 4.78455, 
    4.783514, 4.786196, 4.792386, 4.801616, 4.813207, 4.826326, 4.840052, 
    4.853444, 4.865614, 4.875832, 4.883608, 4.8888, 4.891662, 4.892874, 
    4.893465,
  // momentumY(17,8, 0-49)
    4.928143, 4.912886, 4.900441, 4.890904, 4.884245, 4.880311, 4.878841, 
    4.87951, 4.88195, 4.885783, 4.890644, 4.89619, 4.902103, 4.908071, 
    4.913764, 4.915773, 4.92422, 4.927168, 4.928677, 4.928949, 4.927879, 
    4.927794, 4.925365, 4.920992, 4.914267, 4.905104, 4.893435, 4.879482, 
    4.863534, 4.846408, 4.828302, 4.813304, 4.799834, 4.788882, 4.781299, 
    4.777662, 4.778239, 4.782969, 4.791487, 4.803172, 4.817198, 4.83261, 
    4.848373, 4.863461, 4.876935, 4.88804, 4.896313, 4.901678, 4.904503, 
    4.905589,
  // momentumY(17,9, 0-49)
    4.926387, 4.91217, 4.900692, 4.892024, 4.88611, 4.882786, 4.881791, 
    4.882813, 4.88551, 4.889541, 4.894586, 4.900361, 4.906602, 4.913068, 
    4.919524, 4.921489, 4.929521, 4.933596, 4.936105, 4.937315, 4.937177, 
    4.938101, 4.936598, 4.933035, 4.927056, 4.918464, 4.90711, 4.893102, 
    4.876647, 4.85835, 4.838352, 4.821018, 4.804783, 4.790828, 4.780226, 
    4.773788, 4.771987, 4.774931, 4.782368, 4.793742, 4.808257, 4.824928, 
    4.84266, 4.860311, 4.876772, 4.891061, 4.902427, 4.910475, 4.915247, 
    4.917273,
  // momentumY(17,10, 0-49)
    4.923273, 4.910128, 4.899665, 4.891922, 4.886822, 4.884184, 4.883743, 
    4.885196, 4.888224, 4.892519, 4.897807, 4.903848, 4.910443, 4.917434, 
    4.924696, 4.92671, 4.934017, 4.939202, 4.942721, 4.944888, 4.945706, 
    4.947608, 4.947049, 4.944363, 4.939278, 4.931495, 4.920787, 4.907132, 
    4.890639, 4.871647, 4.850207, 4.83084, 4.812048, 4.795187, 4.781552, 
    4.772192, 4.767801, 4.768667, 4.774671, 4.785334, 4.799887, 4.817338, 
    4.836549, 4.856289, 4.875316, 4.892464, 4.906739, 4.917458, 4.924351, 
    4.92766,
  // momentumY(17,11, 0-49)
    4.918819, 4.906762, 4.897353, 4.890594, 4.886381, 4.884509, 4.884711, 
    4.886684, 4.890129, 4.89476, 4.90034, 4.906679, 4.913639, 4.921144, 
    4.929193, 4.931473, 4.937835, 4.944029, 4.948521, 4.951626, 4.953395, 
    4.95619, 4.956545, 4.954758, 4.950663, 4.943872, 4.934094, 4.921172, 
    4.905105, 4.885919, 4.863553, 4.842531, 4.821484, 4.801915, 4.785327, 
    4.773007, 4.765884, 4.764438, 4.768693, 4.778259, 4.792406, 4.810146, 
    4.830305, 4.851591, 4.872667, 4.89222, 4.909069, 4.922284, 4.931321, 
    4.936136,
  // momentumY(17,12, 0-49)
    4.913151, 4.902174, 4.89384, 4.888111, 4.884847, 4.883822, 4.884756, 
    4.887339, 4.891278, 4.896312, 4.90223, 4.908882, 4.91619, 4.924158, 
    4.932895, 4.935816, 4.941145, 4.948177, 4.953555, 4.957557, 4.960253, 
    4.96382, 4.965019, 4.964102, 4.961035, 4.955356, 4.946728, 4.934856, 
    4.919626, 4.900735, 4.877989, 4.855725, 4.832791, 4.810797, 4.791426, 
    4.776199, 4.766277, 4.762349, 4.764593, 4.772719, 4.786045, 4.803592, 
    4.82417, 4.846443, 4.869005, 4.890441, 4.90943, 4.924849, 4.935921, 
    4.942349,
  // momentumY(17,13, 0-49)
    4.906466, 4.896542, 4.889278, 4.884605, 4.882339, 4.882226, 4.883963, 
    4.887234, 4.891738, 4.897228, 4.903514, 4.91048, 4.918095, 4.926425, 
    4.93566, 4.939777, 4.944144, 4.951789, 4.95794, 4.962779, 4.966364, 
    4.970561, 4.972504, 4.972393, 4.970335, 4.96582, 4.958477, 4.947888, 
    4.933827, 4.915659, 4.893061, 4.869974, 4.845552, 4.821473, 4.799566, 
    4.781562, 4.768855, 4.762346, 4.762383, 4.768782, 4.78092, 4.797838, 
    4.818337, 4.841057, 4.864547, 4.887329, 4.907979, 4.925239, 4.938151, 
    4.946199,
  // momentumY(17,14, 0-49)
    4.899024, 4.89009, 4.883871, 4.880249, 4.879004, 4.879846, 4.882438, 
    4.886447, 4.891568, 4.897552, 4.90422, 4.911483, 4.919337, 4.927886, 
    4.937351, 4.943377, 4.947018, 4.955034, 4.961828, 4.967443, 4.971882, 
    4.976558, 4.979132, 4.979733, 4.97862, 4.975255, 4.969245, 4.960069, 
    4.947399, 4.930287, 4.908312, 4.884778, 4.859268, 4.833473, 4.809331, 
    4.788751, 4.773347, 4.764234, 4.761935, 4.766388, 4.777039, 4.792955, 
    4.812939, 4.835619, 4.859524, 4.883137, 4.904978, 4.923697, 4.9382, 
    4.947796,
  // momentumY(17,15, 0-49)
    4.891112, 4.883087, 4.877852, 4.875248, 4.875012, 4.876813, 4.880279, 
    4.885053, 4.890813, 4.897305, 4.904356, 4.911882, 4.919893, 4.928493, 
    4.93788, 4.946609, 4.949912, 4.958069, 4.965397, 4.97174, 4.97701, 
    4.982026, 4.985116, 4.986323, 4.986053, 4.983757, 4.979042, 4.971297, 
    4.960118, 4.944283, 4.923313, 4.899639, 4.873401, 4.84626, 4.820212, 
    4.797309, 4.779364, 4.767699, 4.763014, 4.76538, 4.774317, 4.788934, 
    4.808044, 4.830278, 4.854156, 4.87815, 4.900752, 4.920557, 4.936386, 
    4.947409,
  // momentumY(17,16, 0-49)
    4.883029, 4.875806, 4.871468, 4.869812, 4.870532, 4.873254, 4.877571, 
    4.883094, 4.889482, 4.896476, 4.903892, 4.911646, 4.919736, 4.928235, 
    4.937255, 4.949426, 4.952873, 4.96102, 4.968817, 4.975876, 4.981983, 
    4.987225, 4.990734, 4.992444, 4.992887, 4.991526, 4.987975, 4.981569, 
    4.971848, 4.957378, 4.937684, 4.914083, 4.887414, 4.859268, 4.831649, 
    4.806712, 4.786437, 4.772339, 4.765296, 4.765512, 4.772596, 4.785703, 
    4.803671, 4.825141, 4.84864, 4.872643, 4.89564, 4.916207, 4.933103, 
    4.945402,
  // momentumY(17,17, 0-49)
    4.875055, 4.868514, 4.864955, 4.864135, 4.86571, 4.869261, 4.87435, 
    4.880558, 4.88753, 4.89499, 4.902754, 4.910722, 4.918859, 4.927171, 
    4.935653, 4.951737, 4.955822, 4.963933, 4.972224, 4.980051, 4.987048, 
    4.992446, 4.996313, 4.998434, 4.999444, 4.99883, 4.99623, 4.990953, 
    4.982525, 4.969369, 4.951089, 4.927674, 4.900793, 4.871935, 4.843071, 
    4.816412, 4.794065, 4.777717, 4.768412, 4.766494, 4.771667, 4.783143, 
    4.799794, 4.820279, 4.843141, 4.866875, 4.889984, 4.911039, 4.928771, 
    4.942188,
  // momentumY(17,18, 0-49)
    4.867438, 4.861432, 4.858498, 4.858359, 4.860627, 4.864854, 4.870573, 
    4.87735, 4.884819, 4.892704, 4.900818, 4.909043, 4.917301, 4.925497, 
    4.93346, 4.953443, 4.958536, 4.966762, 4.975693, 4.984436, 4.992451, 
    4.997995, 5.002215, 5.004687, 5.006111, 5.006001, 5.004041, 4.999564, 
    4.992125, 4.980086, 4.963223, 4.940009, 4.913056, 4.88373, 4.853928, 
    4.825867, 4.801744, 4.783382, 4.771981, 4.768018, 4.771304, 4.781112, 
    4.796357, 4.815728, 4.83779, 4.861065, 4.884079, 4.905415, 4.923792, 
    4.938173,
  // momentumY(17,19, 0-49)
    4.860362, 4.854715, 4.852209, 4.85253, 4.855262, 4.859932, 4.866065, 
    4.87323, 4.881079, 4.889356, 4.89789, 4.906549, 4.915184, 4.923564, 
    4.931289, 4.954461, 4.960647, 4.969331, 4.979218, 4.989158, 4.998429, 
    5.004205, 5.008854, 5.011667, 5.013352, 5.01345, 5.011711, 5.007554, 
    5.000636, 4.989366, 4.973771, 4.950686, 4.92374, 4.894152, 4.863704, 
    4.834578, 4.809007, 4.788918, 4.775646, 4.769795, 4.771284, 4.77946, 
    4.793291, 4.811497, 4.83268, 4.855388, 4.878173, 4.899641, 4.918513, 
    4.933718,
  // momentumY(17,20, 0-49)
    4.854655, 4.849918, 4.84861, 4.850455, 4.855026, 4.861779, 4.870096, 
    4.879328, 4.888843, 4.898059, 4.906477, 4.913717, 4.919533, 4.923843, 
    4.926725, 0, 4.976701, 4.980468, 4.985542, 4.99134, 4.997496, 5.000072, 
    5.003079, 5.005518, 5.008004, 5.009818, 5.010391, 5.008807, 5.004483, 
    4.995662, 4.982596, 4.960472, 4.934066, 4.904542, 4.873656, 4.843603, 
    4.816685, 4.794946, 4.779853, 4.772143, 4.771838, 4.778371, 4.790754, 
    4.807751, 4.827991, 4.850053, 4.872515, 4.894001, 4.913239, 4.929135,
  // momentumY(17,21, 0-49)
    4.849359, 4.844958, 4.844018, 4.846222, 4.851108, 4.858102, 4.866564, 
    4.875849, 4.885345, 4.89451, 4.90289, 4.910137, 4.916014, 4.920402, 
    4.923314, 0, 4.978804, 4.983113, 4.98882, 4.995245, 5.001908, 5.003341, 
    5.005481, 5.007151, 5.009163, 5.010862, 5.011708, 5.010763, 5.007414, 
    4.999859, 4.988595, 4.967202, 4.941577, 4.912706, 4.882171, 4.852049, 
    4.824604, 4.801916, 4.785548, 4.776368, 4.774518, 4.77953, 4.790494, 
    4.806223, 4.825388, 4.846598, 4.868461, 4.889622, 4.908823, 4.924966,
  // momentumY(17,22, 0-49)
    4.84491, 4.840719, 4.840024, 4.842488, 4.847629, 4.854852, 4.863504, 
    4.872935, 4.882536, 4.891777, 4.900223, 4.907533, 4.913461, 4.917856, 
    4.920673, 0, 4.980448, 4.985187, 4.991485, 4.998569, 5.005846, 5.006361, 
    5.007894, 5.009054, 5.010793, 5.012468, 5.013533, 5.01302, 5.010294, 
    5.003533, 4.9935, 4.972336, 4.947056, 4.918531, 4.888209, 4.858057, 
    4.830273, 4.806931, 4.789643, 4.779356, 4.776308, 4.780115, 4.789931, 
    4.804622, 4.822892, 4.843383, 4.864727, 4.885594, 4.904738, 4.921063,
  // momentumY(17,23, 0-49)
    4.841343, 4.837268, 4.836722, 4.839362, 4.844692, 4.852111, 4.860959, 
    4.870574, 4.880348, 4.889748, 4.898341, 4.905778, 4.911798, 4.916217, 
    4.918941, 0, 4.982242, 4.987259, 4.993968, 5.001531, 5.009266, 5.00898, 
    5.009981, 5.010692, 5.012161, 5.013753, 5.014909, 5.014637, 5.012286, 
    5.006017, 4.996813, 4.975653, 4.950515, 4.922195, 4.892049, 4.861947, 
    4.834018, 4.810307, 4.792441, 4.781416, 4.77753, 4.780464, 4.789426, 
    4.803322, 4.820889, 4.840794, 4.86169, 4.882262, 4.901279, 4.917653,
  // momentumY(17,24, 0-49)
    4.838642, 4.834622, 4.834155, 4.836901, 4.842365, 4.849943, 4.858972, 
    4.868788, 4.878774, 4.888392, 4.897195, 4.904826, 4.911006, 4.915524, 
    4.918251, 0, 4.984415, 4.98959, 4.996536, 5.004384, 5.012406, 5.011586, 
    5.012234, 5.012639, 5.013902, 5.015387, 5.016535, 5.016338, 5.014139, 
    5.008089, 4.999325, 4.978053, 4.952898, 4.924624, 4.894527, 4.864416, 
    4.836373, 4.812413, 4.794162, 4.782639, 4.778178, 4.7805, 4.788852, 
    4.80217, 4.819218, 4.838678, 4.859221, 4.879544, 4.898427, 4.914783,
  // momentumY(17,25, 0-49)
    4.836769, 4.832759, 4.832325, 4.83513, 4.840688, 4.8484, 4.857604, 
    4.867634, 4.877865, 4.887749, 4.896824, 4.904718, 4.911138, 4.915858, 
    4.918736, 0, 4.986551, 4.991792, 4.998822, 5.006766, 5.014881, 5.013883, 
    5.014416, 5.014708, 5.015873, 5.017272, 5.018345, 5.018085, 5.015834, 
    5.009744, 5.001011, 4.979569, 4.954289, 4.925926, 4.895759, 4.865575, 
    4.83743, 4.813322, 4.794866, 4.783079, 4.778309, 4.780292, 4.788291, 
    4.801262, 4.817979, 4.837139, 4.85742, 4.877531, 4.89625, 4.912501,
  // momentumY(17,26, 0-49)
    4.835672, 4.83165, 4.831218, 4.834058, 4.839693, 4.847535, 4.856926, 
    4.867199, 4.877722, 4.887929, 4.897342, 4.905571, 4.912312, 4.917341, 
    4.920526, 0, 4.988527, 4.993752, 5.000716, 5.008561, 5.016568, 5.015782, 
    5.016457, 5.016857, 5.018059, 5.019417, 5.020375, 5.019933, 5.017445, 
    5.011068, 5.001957, 4.980327, 4.954838, 4.92627, 4.895921, 4.865594, 
    4.837351, 4.813177, 4.794672, 4.782838, 4.778008, 4.779906, 4.787796, 
    4.800632, 4.817194, 4.836185, 4.856286, 4.876206, 4.894732, 4.910787,
  // momentumY(17,27, 0-49)
    4.835305, 4.831254, 4.830816, 4.833688, 4.83941, 4.847407, 4.857031, 
    4.86761, 4.878496, 4.889104, 4.898934, 4.907572, 4.914705, 4.920119, 
    4.923718, 0, 4.990418, 4.995515, 5.002238, 5.00977, 5.01746, 5.017213, 
    5.018252, 5.01895, 5.020303, 5.021653, 5.022446, 5.021699, 5.018786, 
    5.011879, 5.002003, 4.980161, 4.954391, 4.925523, 4.894915, 4.864421, 
    4.836125, 4.812012, 4.793656, 4.782018, 4.777392, 4.779467, 4.787487, 
    4.800394, 4.816962, 4.835893, 4.855869, 4.875599, 4.893869, 4.909608,
  // momentumY(17,28, 0-49)
    4.835628, 4.831538, 4.831094, 4.834014, 4.839862, 4.848079, 4.85802, 
    4.869009, 4.880377, 4.891504, 4.90185, 4.910967, 4.91853, 4.924347, 
    4.928369, 0, 4.992599, 4.997404, 5.003668, 5.010651, 5.017807, 5.018314, 
    5.019859, 5.020988, 5.022568, 5.023917, 5.02448, 5.023301, 5.019778, 
    5.01211, 5.00112, 4.979014, 4.952876, 4.923621, 4.892708, 4.862062, 
    4.833807, 4.809922, 4.791938, 4.780753, 4.776589, 4.779086, 4.787449, 
    4.8006, 4.817302, 4.836254, 4.856133, 4.875648, 4.893589, 4.908889,
  // momentumY(17,29, 0-49)
    4.836607, 4.832465, 4.832018, 4.835017, 4.841056, 4.849597, 4.859998, 
    4.871566, 4.883592, 4.8954, 4.906381, 4.916035, 4.924014, 4.930147, 
    4.934448, 0, 4.994762, 4.999057, 5.004619, 5.010811, 5.01722, 5.01852, 
    5.020604, 5.022212, 5.02405, 5.025388, 5.025658, 5.023925, 5.019612, 
    5.010951, 4.998516, 4.976011, 4.949397, 4.919718, 4.888555, 4.857924, 
    4.829979, 4.806665, 4.789436, 4.779088, 4.77575, 4.778986, 4.787952, 
    4.80154, 4.818505, 4.837532, 4.857296, 4.876508, 4.89396, 4.908601,
  // momentumY(17,30, 0-49)
    4.837832, 4.833149, 4.831962, 4.833973, 4.838768, 4.84586, 4.854743, 
    4.86493, 4.875998, 4.887613, 4.899509, 4.911485, 4.923332, 4.93478, 
    4.945404, 4.975517, 4.979926, 4.9902, 5.001615, 5.01291, 5.023316, 
    5.028723, 5.033325, 5.036073, 5.037669, 5.037555, 5.035443, 5.030748, 
    5.023216, 5.011344, 4.995587, 4.971336, 4.943355, 4.912786, 4.881282, 
    4.850867, 4.823629, 4.801392, 4.785451, 4.776451, 4.77439, 4.778745, 
    4.788615, 4.802867, 4.820241, 4.839418, 4.859073, 4.87792, 4.894762, 
    4.908581,
  // momentumY(17,31, 0-49)
    4.840512, 4.836057, 4.835127, 4.837435, 4.842564, 4.85002, 4.85927, 
    4.869801, 4.881155, 4.892956, 4.904926, 4.916868, 4.928643, 4.940125, 
    4.951134, 4.976396, 4.981072, 4.990958, 5.001443, 5.011515, 5.020609, 
    5.025819, 5.029953, 5.032291, 5.033554, 5.033181, 5.03083, 5.025838, 
    5.017842, 5.005279, 4.988306, 4.964038, 4.936157, 4.905926, 4.875092, 
    4.845701, 4.81979, 4.799075, 4.784719, 4.777233, 4.77651, 4.781954, 
    4.792624, 4.80736, 4.824892, 4.843892, 4.863036, 4.881039, 4.896733, 
    4.90915,
  // momentumY(17,32, 0-49)
    4.84394, 4.839687, 4.838961, 4.84147, 4.8468, 4.854445, 4.863869, 
    4.874544, 4.886004, 4.897867, 4.909857, 4.921802, 4.933619, 4.9453, 
    4.956847, 4.976905, 4.981479, 4.991234, 5.00101, 5.010061, 5.018018, 
    5.023118, 5.026866, 5.028792, 5.02958, 5.028664, 5.025671, 5.019921, 
    5.011018, 4.997434, 4.979104, 4.954812, 4.927166, 4.897542, 4.867736, 
    4.839773, 4.815597, 4.796778, 4.784322, 4.7786, 4.779403, 4.786065, 
    4.797607, 4.812852, 4.830517, 4.849267, 4.867775, 4.88477, 4.899115, 
    4.909908,
  // momentumY(17,33, 0-49)
    4.848188, 4.844136, 4.843581, 4.846228, 4.851653, 4.859349, 4.868777, 
    4.879411, 4.890791, 4.902544, 4.914413, 4.926251, 4.938032, 4.949833, 
    4.961806, 4.976944, 4.981427, 4.991122, 5.000261, 5.008378, 5.015282, 
    5.02028, 5.023657, 5.025142, 5.025333, 5.023657, 5.019734, 5.012911, 
    5.002809, 4.988014, 4.968327, 4.944061, 4.916827, 4.88808, 4.859641, 
    4.83347, 4.811376, 4.794761, 4.784458, 4.780696, 4.783165, 4.791138, 
    4.803601, 4.819355, 4.837107, 4.855516, 4.87325, 4.889057, 4.901842, 
    4.910791,
  // momentumY(17,34, 0-49)
    4.853289, 4.849438, 4.849027, 4.851749, 4.857172, 4.864788, 4.874062, 
    4.88448, 4.895594, 4.907053, 4.91862, 4.930174, 4.941731, 4.953428, 
    4.965522, 4.976438, 4.981064, 4.990592, 4.999053, 5.006239, 5.012118, 
    5.01695, 5.019924, 5.020919, 5.020409, 5.017825, 5.01279, 5.004707, 
    4.993249, 4.9772, 4.956297, 4.932189, 4.905595, 4.878024, 4.85128, 
    4.827223, 4.8075, 4.793324, 4.785354, 4.783679, 4.787896, 4.797219, 
    4.810601, 4.826828, 4.844588, 4.862535, 4.879337, 4.893764, 4.904784, 
    4.911689,
  // momentumY(17,35, 0-49)
    4.859222, 4.855562, 4.855252, 4.857974, 4.863289, 4.870693, 4.879658, 
    4.889689, 4.900362, 4.911344, 4.922421, 4.933497, 4.944608, 4.955915, 
    4.967728, 4.975316, 4.980386, 4.989532, 4.997201, 5.003416, 5.00826, 
    5.012824, 5.015333, 5.015789, 5.014503, 5.010921, 5.004682, 4.995273, 
    4.982435, 4.965222, 4.943371, 4.919636, 4.893962, 4.867884, 4.843148, 
    4.82148, 4.804347, 4.792766, 4.787225, 4.787683, 4.793653, 4.804296, 
    4.81854, 4.835147, 4.852794, 4.870125, 4.885816, 4.898671, 4.907736, 
    4.912441,
  // momentumY(17,36, 0-49)
    4.865902, 4.862398, 4.862123, 4.86475, 4.869839, 4.876892, 4.885399, 
    4.894885, 4.904952, 4.915292, 4.925711, 4.936127, 4.946576, 4.957216, 
    4.968345, 4.973502, 4.979285, 4.987776, 4.994511, 4.999691, 5.003481, 
    5.007654, 5.009626, 5.009497, 5.007393, 5.002791, 4.995346, 4.984653, 
    4.97054, 4.952381, 4.929957, 4.90688, 4.882451, 4.858187, 4.835741, 
    4.816682, 4.802279, 4.793364, 4.790259, 4.792812, 4.800456, 4.812315, 
    4.827287, 4.844121, 4.861478, 4.877997, 4.892375, 4.903469, 4.910425, 
    4.912837,
  // momentumY(17,37, 0-49)
    4.873171, 4.869758, 4.869428, 4.871847, 4.876582, 4.883149, 4.891055, 
    4.899855, 4.909174, 4.918733, 4.928355, 4.93796, 4.947573, 4.957314, 
    4.967422, 4.970922, 4.977585, 4.98515, 4.990809, 4.994896, 4.997612, 
    5.001259, 5.002623, 5.001882, 4.998955, 4.993373, 4.984812, 4.972988, 
    4.957819, 4.939039, 4.916505, 4.894428, 4.871589, 4.849447, 4.829532, 
    4.813232, 4.801623, 4.795353, 4.794603, 4.799121, 4.808279, 4.821166, 
    4.836657, 4.853489, 4.870317, 4.885788, 4.898634, 4.907787, 4.91253, 
    4.912643,
  // momentumY(17,38, 0-49)
    4.880799, 4.877385, 4.876884, 4.878968, 4.88322, 4.889169, 4.896352, 
    4.904349, 4.912816, 4.921493, 4.930215, 4.938902, 4.947552, 4.956231, 
    4.965086, 4.967517, 4.975098, 4.981501, 4.985966, 4.988914, 4.990543, 
    4.993541, 4.994239, 4.992883, 4.989176, 4.982718, 4.973215, 4.960507, 
    4.944603, 4.925617, 4.903484, 4.88278, 4.861875, 4.842131, 4.824929, 
    4.811468, 4.802634, 4.798907, 4.800348, 4.806618, 4.817043, 4.830686, 
    4.846407, 4.862938, 4.878937, 4.893082, 4.904164, 4.911223, 4.913716, 
    4.911637,
  // momentumY(17,39, 0-49)
    4.8885, 4.884964, 4.884163, 4.885783, 4.889422, 4.894643, 4.901007, 
    4.908122, 4.915665, 4.923398, 4.931163, 4.938869, 4.946483, 4.95401, 
    4.961489, 4.963247, 4.971654, 4.976719, 4.979917, 4.981703, 4.982242, 
    4.984488, 4.984486, 4.982543, 4.978146, 4.970976, 4.960778, 4.947517, 
    4.931282, 4.912557, 4.891349, 4.872391, 4.853734, 4.836616, 4.822244, 
    4.811627, 4.805473, 4.804114, 4.807503, 4.815238, 4.826606, 4.840658, 
    4.856246, 4.87211, 4.886935, 4.899451, 4.908543, 4.913409, 4.913702, 
    4.909656,
  // momentumY(17,40, 0-49)
    4.895968, 4.892166, 4.890924, 4.891946, 4.894863, 4.899263, 4.90474, 
    4.910928, 4.917522, 4.924296, 4.931087, 4.937795, 4.944351, 4.950702, 
    4.956784, 4.958094, 4.967124, 4.970757, 4.972659, 4.973285, 4.972751, 
    4.974173, 4.973469, 4.971002, 4.966048, 4.958385, 4.947799, 4.934374, 
    4.918255, 4.900277, 4.880496, 4.863629, 4.847486, 4.833153, 4.821659, 
    4.813825, 4.810189, 4.810955, 4.815989, 4.824837, 4.836764, 4.850812, 
    4.865849, 4.880637, 4.893913, 4.904496, 4.911415, 4.914057, 4.912313, 
    4.906664,
  // momentumY(17,41, 0-49)
    4.902921, 4.898695, 4.89686, 4.897158, 4.899249, 4.902759, 4.907311, 
    4.91256, 4.918214, 4.924046, 4.929891, 4.935626, 4.941149, 4.946351, 
    4.951089, 4.952054, 4.96143, 4.963621, 4.964247, 4.963741, 4.962173, 
    4.962739, 4.96137, 4.958476, 4.95314, 4.945245, 4.934614, 4.921438, 
    4.905893, 4.88913, 4.871221, 4.856738, 4.843309, 4.831854, 4.823215, 
    4.818036, 4.816703, 4.819304, 4.825633, 4.835196, 4.847248, 4.860843, 
    4.874875, 4.888161, 4.899525, 4.907917, 4.912551, 4.913051, 4.909559, 
    4.9028,
  // momentumY(17,42, 0-49)
    4.909159, 4.904336, 4.901761, 4.901208, 4.902383, 4.904947, 4.90855, 
    4.912868, 4.917612, 4.922549, 4.9275, 4.932313, 4.936859, 4.940983, 
    4.944482, 4.945125, 4.954541, 4.955351, 4.954765, 4.953189, 4.95065, 
    4.950379, 4.948419, 4.945224, 4.939711, 4.931865, 4.921547, 4.909028, 
    4.894497, 4.879364, 4.863691, 4.851813, 4.841222, 4.832664, 4.826799, 
    4.8241, 4.824811, 4.828923, 4.836165, 4.846019, 4.857746, 4.870423, 
    4.883003, 4.894386, 4.903529, 4.90956, 4.911921, 4.910494, 4.905684, 
    4.898421,
  // momentumY(17,43, 0-49)
    4.914628, 4.909033, 4.905563, 4.904037, 4.904203, 4.905764, 4.908397, 
    4.91179, 4.915656, 4.919752, 4.923867, 4.927831, 4.931473, 4.934608, 
    4.936998, 4.937302, 4.946457, 4.946009, 4.944318, 4.94176, 4.938349, 
    4.937307, 4.934862, 4.93152, 4.926051, 4.91854, 4.908878, 4.897394, 
    4.884263, 4.871099, 4.857931, 4.848797, 4.84109, 4.835384, 4.832156, 
    4.83172, 4.834194, 4.839475, 4.847241, 4.856964, 4.867921, 4.879242, 
    4.889966, 4.899126, 4.905847, 4.909483, 4.909735, 4.906756, 4.901185, 
    4.894104,
  // momentumY(17,44, 0-49)
    4.919461, 4.912925, 4.908408, 4.905779, 4.904836, 4.90532, 4.90694, 
    4.909394, 4.912395, 4.915678, 4.919009, 4.92218, 4.924991, 4.92723, 
    4.928645, 4.928577, 4.937214, 4.935669, 4.933005, 4.929586, 4.925431, 
    4.923725, 4.920937, 4.917611, 4.91241, 4.905505, 4.896807, 4.88668, 
    4.875265, 4.864319, 4.85382, 4.847488, 4.84264, 4.839678, 4.838911, 
    4.8405, 4.844442, 4.850554, 4.858476, 4.867672, 4.877462, 4.887057, 
    4.895621, 4.902356, 4.906611, 4.907991, 4.906475, 4.902468, 4.896797, 
    4.890616,
  // momentumY(17,45, 0-49)
    4.924008, 4.916375, 4.910664, 4.906796, 4.904622, 4.903929, 4.904456, 
    4.905918, 4.908018, 4.910478, 4.913033, 4.91544, 4.91747, 4.918889, 
    4.919441, 4.918964, 4.926886, 4.924419, 4.920935, 4.916797, 4.912052, 
    4.909824, 4.906849, 4.903707, 4.898986, 4.892923, 4.885447, 4.876929, 
    4.86746, 4.858889, 4.851131, 4.847575, 4.845493, 4.84512, 4.846608, 
    4.849974, 4.855102, 4.861737, 4.869482, 4.877822, 4.886137, 4.893749, 
    4.899987, 4.904269, 4.906194, 4.90565, 4.902875, 4.898486, 4.893424, 
    4.888831,
  // momentumY(17,46, 0-49)
    4.928825, 4.919962, 4.912918, 4.90767, 4.904126, 4.902122, 4.90143, 
    4.901784, 4.902892, 4.904456, 4.906185, 4.907807, 4.909061, 4.909698, 
    4.909465, 4.908536, 4.915604, 4.912388, 4.908238, 4.903537, 4.898368, 
    4.895784, 4.892784, 4.88998, 4.885921, 4.880892, 4.874827, 4.868092, 
    4.860718, 4.854588, 4.849548, 4.848677, 4.849215, 4.851243, 4.854764, 
    4.859663, 4.865725, 4.87262, 4.879941, 4.887194, 4.89385, 4.899375, 
    4.903301, 4.905291, 4.905223, 4.903256, 4.899861, 4.895799, 4.892039, 
    4.889628,
  // momentumY(17,47, 0-49)
    4.934628, 4.924436, 4.915936, 4.909171, 4.904103, 4.900622, 4.898542, 
    4.897622, 4.897577, 4.898103, 4.89889, 4.899638, 4.900064, 4.899903, 
    4.898912, 4.897471, 4.903601, 4.899779, 4.895105, 4.889996, 4.884573, 
    4.881795, 4.878922, 4.876583, 4.873326, 4.869465, 4.864933, 4.860072, 
    4.85486, 4.851156, 4.848743, 4.850405, 4.853375, 4.857594, 4.862926, 
    4.869143, 4.875928, 4.882905, 4.889649, 4.895721, 4.900694, 4.904212, 
    4.906034, 4.906089, 4.904534, 4.901772, 4.898455, 4.895413, 4.893567, 
    4.893793,
  // momentumY(17,48, 0-49)
    4.942206, 4.930628, 4.920584, 4.912177, 4.905432, 4.900293, 4.896624, 
    4.894217, 4.892807, 4.892093, 4.891754, 4.891472, 4.890954, 4.889923, 
    4.888144, 4.886106, 4.891249, 4.886915, 4.881835, 4.876449, 4.870919, 
    4.868098, 4.865475, 4.863686, 4.861314, 4.858688, 4.855734, 4.852766, 
    4.84971, 4.848352, 4.848417, 4.852421, 4.857611, 4.863803, 4.870745, 
    4.878098, 4.885471, 4.89244, 4.898585, 4.903532, 4.906981, 4.908762, 
    4.908873, 4.907512, 4.905091, 4.902219, 4.899659, 4.898243, 4.898774, 
    4.901918,
  // momentumY(17,49, 0-49)
    4.959617, 4.946238, 4.934052, 4.923233, 4.913883, 4.906022, 4.89959, 
    4.894449, 4.890389, 4.887144, 4.884412, 4.881876, 4.879222, 4.876143, 
    4.872361, 4.869101, 4.880398, 4.874001, 4.866947, 4.860031, 4.853502, 
    4.852767, 4.852791, 4.85458, 4.855067, 4.854731, 4.853221, 4.850918, 
    4.847435, 4.846223, 4.846673, 4.853611, 4.861576, 4.870242, 4.879228, 
    4.888075, 4.896299, 4.903437, 4.909089, 4.912979, 4.914989, 4.915207, 
    4.913942, 4.911713, 4.909215, 4.907247, 4.906631, 4.908108, 4.91226, 
    4.919442,
  // momentumY(18,0, 0-49)
    4.884809, 4.871144, 4.860725, 4.853534, 4.849423, 4.848121, 4.849251, 
    4.852354, 4.856926, 4.862458, 4.868456, 4.874484, 4.880164, 4.885192, 
    4.88933, 4.892411, 4.895638, 4.896484, 4.896322, 4.895182, 4.893073, 
    4.890365, 4.886718, 4.882278, 4.87701, 4.871042, 4.864499, 4.857598, 
    4.850573, 4.843819, 4.837571, 4.832456, 4.82845, 4.825788, 4.824625, 
    4.825011, 4.826875, 4.830015, 4.834108, 4.838731, 4.843399, 4.84762, 
    4.850959, 4.853108, 4.853957, 4.853652, 4.852622, 4.851551, 4.851324, 
    4.852911,
  // momentumY(18,1, 0-49)
    4.884934, 4.871832, 4.862022, 4.855465, 4.85199, 4.851309, 4.853025, 
    4.856676, 4.861752, 4.867746, 4.874176, 4.880609, 4.886672, 4.892051, 
    4.896487, 4.899747, 4.904272, 4.905182, 4.905079, 4.903979, 4.901849, 
    4.899334, 4.895684, 4.891092, 4.885404, 4.878729, 4.871161, 4.862932, 
    4.854278, 4.845744, 4.837555, 4.830768, 4.825129, 4.820971, 4.818543, 
    4.817976, 4.819256, 4.822213, 4.826527, 4.831753, 4.837351, 4.842746, 
    4.847396, 4.850862, 4.852898, 4.853511, 4.853005, 4.851987, 4.851309, 
    4.851967,
  // momentumY(18,2, 0-49)
    4.886409, 4.873914, 4.864717, 4.858756, 4.855839, 4.85566, 4.857812, 
    4.861832, 4.867219, 4.87348, 4.880151, 4.886819, 4.893123, 4.898752, 
    4.903427, 4.906798, 4.912543, 4.913613, 4.913682, 4.912762, 4.910775, 
    4.908639, 4.905188, 4.900646, 4.894743, 4.887562, 4.879149, 4.869736, 
    4.859549, 4.849249, 4.839058, 4.830468, 4.823002, 4.817106, 4.813138, 
    4.811329, 4.811743, 4.814265, 4.818604, 4.82431, 4.830813, 4.837478, 
    4.84367, 4.848833, 4.852573, 4.854734, 4.855453, 4.855189, 4.854686, 
    4.854899,
  // momentumY(18,3, 0-49)
    4.888647, 4.876785, 4.868192, 4.862783, 4.86035, 4.860566, 4.863028, 
    4.867271, 4.872816, 4.879192, 4.885966, 4.892745, 4.899195, 4.905011, 
    4.909902, 4.913323, 4.920159, 4.921499, 4.921853, 4.921245, 4.919561, 
    4.917976, 4.914915, 4.910623, 4.904731, 4.897276, 4.888249, 4.877862, 
    4.866318, 4.854356, 4.842188, 4.831735, 4.822308, 4.814471, 4.808708, 
    4.805367, 4.804612, 4.806405, 4.810504, 4.816482, 4.823758, 4.831663, 
    4.839493, 4.846585, 4.852404, 4.856616, 4.859165, 4.860306, 4.860612, 
    4.860924,
  // momentumY(18,4, 0-49)
    4.89114, 4.879928, 4.871926, 4.867028, 4.865009, 4.865537, 4.868205, 
    4.872565, 4.878159, 4.884547, 4.891326, 4.898142, 4.904681, 4.910653, 
    4.915773, 4.919184, 4.926921, 4.92865, 4.929398, 4.929215, 4.927966, 
    4.927078, 4.924573, 4.920717, 4.91506, 4.907583, 4.898214, 4.887125, 
    4.874485, 4.861058, 4.847029, 4.834742, 4.823296, 4.813377, 4.805604, 
    4.800458, 4.798227, 4.798971, 4.802519, 4.808488, 4.816317, 4.825317, 
    4.834739, 4.843832, 4.851933, 4.858536, 4.863369, 4.866457, 4.868152, 
    4.869117,
  // momentumY(18,5, 0-49)
    4.893487, 4.882936, 4.875515, 4.871094, 4.869439, 4.870214, 4.873019, 
    4.877421, 4.882993, 4.889328, 4.89606, 4.90287, 4.909472, 4.915598, 
    4.920979, 4.924315, 4.932712, 4.934937, 4.936172, 4.936502, 4.935794, 
    4.935705, 4.933889, 4.930626, 4.925414, 4.918171, 4.908759, 4.897293, 
    4.883885, 4.869284, 4.853611, 4.839611, 4.826176, 4.814109, 4.80417, 
    4.796988, 4.792989, 4.792358, 4.795018, 4.800653, 4.808738, 4.818592, 
    4.829433, 4.840447, 4.85086, 4.860002, 4.867395, 4.872821, 4.876379, 
    4.878513,
  // momentumY(18,6, 0-49)
    4.895404, 4.88553, 4.878681, 4.874718, 4.873394, 4.874374, 4.877271, 
    4.881673, 4.887185, 4.893434, 4.900091, 4.906876, 4.913533, 4.919827, 
    4.925513, 4.928716, 4.937472, 4.940289, 4.942079, 4.942984, 4.942886, 
    4.94365, 4.942612, 4.940061, 4.935476, 4.928711, 4.919563, 4.908076, 
    4.894294, 4.878877, 4.861876, 4.846375, 4.831077, 4.816886, 4.8047, 
    4.795306, 4.789286, 4.78697, 4.788401, 4.79335, 4.801349, 4.811738, 
    4.823725, 4.836451, 4.849043, 4.860695, 4.870737, 4.878716, 4.884475, 
    4.888203,
  // momentumY(18,7, 0-49)
    4.896717, 4.887537, 4.881267, 4.877753, 4.876744, 4.877908, 4.880875, 
    4.885259, 4.890693, 4.896843, 4.903419, 4.910171, 4.916884, 4.92336, 
    4.929397, 4.932419, 4.941206, 4.944678, 4.947065, 4.948576, 4.949125, 
    4.950751, 4.950533, 4.948766, 4.944954, 4.938883, 4.930294, 4.919146, 
    4.905412, 4.889598, 4.871658, 4.854958, 4.838015, 4.821816, 4.807391, 
    4.795682, 4.787444, 4.783171, 4.783046, 4.786955, 4.794499, 4.80506, 
    4.81785, 4.831971, 4.846484, 4.860461, 4.873067, 4.88364, 4.891777, 
    4.897409,
  // momentumY(18,8, 0-49)
    4.897334, 4.888876, 4.8832, 4.880144, 4.879449, 4.880795, 4.88383, 
    4.888193, 4.893551, 4.899602, 4.906095, 4.912813, 4.919581, 4.926244, 
    4.932665, 4.935491, 4.943973, 4.948122, 4.951126, 4.953247, 4.954448, 
    4.956897, 4.957495, 4.956541, 4.953597, 4.948393, 4.940624, 4.930164, 
    4.916898, 4.901135, 4.882703, 4.865164, 4.846878, 4.828883, 4.812316, 
    4.798274, 4.78769, 4.78124, 4.779273, 4.781801, 4.788523, 4.798871, 
    4.812071, 4.82721, 4.843288, 4.859285, 4.874232, 4.887288, 4.897826, 
    4.905539,
  // momentumY(18,9, 0-49)
    4.897227, 4.889523, 4.884467, 4.881888, 4.881528, 4.883073, 4.886189, 
    4.890546, 4.895837, 4.901796, 4.908204, 4.914883, 4.921696, 4.928542, 
    4.935356, 4.938022, 4.945889, 4.950691, 4.9543, 4.957017, 4.958854, 
    4.962049, 4.963417, 4.963258, 4.96123, 4.957014, 4.950277, 4.940805, 
    4.928404, 4.913132, 4.894676, 4.876698, 4.85743, 4.837928, 4.819408, 
    4.803104, 4.790129, 4.78135, 4.777303, 4.778151, 4.783701, 4.793451, 
    4.806657, 4.822395, 4.839628, 4.857264, 4.874227, 4.889527, 4.902359, 
    4.912195,
  // momentumY(18,10, 0-49)
    4.896404, 4.88949, 4.885093, 4.883026, 4.883033, 4.884808, 4.888037, 
    4.892411, 4.897654, 4.903532, 4.909855, 4.916485, 4.923323, 4.930325, 
    4.937502, 4.940127, 4.947123, 4.952506, 4.956683, 4.959964, 4.962405, 
    4.966238, 4.968298, 4.968881, 4.967768, 4.964606, 4.959049, 4.950807, 
    4.939605, 4.925227, 4.90721, 4.889191, 4.869336, 4.848673, 4.828465, 
    4.810056, 4.79473, 4.783552, 4.777253, 4.776168, 4.780232, 4.789024, 
    4.80184, 4.817754, 4.835709, 4.854557, 4.873146, 4.890373, 4.905285, 
    4.917168,
  // momentumY(18,11, 0-49)
    4.894901, 4.888815, 4.885118, 4.88361, 4.884029, 4.886082, 4.889462, 
    4.893889, 4.899112, 4.904922, 4.911164, 4.917727, 4.924558, 4.931664, 
    4.939128, 4.941932, 4.947885, 4.95373, 4.958413, 4.962218, 4.965225, 
    4.969569, 4.972219, 4.97346, 4.973217, 4.971121, 4.966827, 4.95998, 
    4.950234, 4.937087, 4.91993, 4.90224, 4.882188, 4.860743, 4.839166, 
    4.818886, 4.801331, 4.787762, 4.779115, 4.775909, 4.778225, 4.785737, 
    4.797791, 4.813478, 4.831725, 4.851353, 4.87115, 4.889936, 4.906639, 
    4.920398,
  // momentumY(18,12, 0-49)
    4.892765, 4.88754, 4.884587, 4.88369, 4.884581, 4.886966, 4.890554, 
    4.89508, 4.900316, 4.906077, 4.912237, 4.918715, 4.925493, 4.932621, 
    4.940238, 4.94356, 4.948406, 4.954556, 4.959667, 4.963951, 4.967489, 
    4.972205, 4.97533, 4.977124, 4.977676, 4.976608, 4.973598, 4.968228, 
    4.960105, 4.94844, 4.9325, 4.915447, 4.895557, 4.873702, 4.851109, 
    4.829243, 4.809653, 4.793781, 4.782765, 4.777319, 4.777685, 4.783647, 
    4.794613, 4.809704, 4.827843, 4.847833, 4.868425, 4.888381, 4.906549, 
    4.921947,
  // momentumY(18,13, 0-49)
    4.890054, 4.885715, 4.88355, 4.883318, 4.884742, 4.887525, 4.891382, 
    4.89606, 4.901348, 4.907085, 4.913165, 4.919536, 4.926205, 4.93325, 
    4.940831, 4.945117, 4.948902, 4.955187, 4.960639, 4.96536, 4.969398, 
    4.97435, 4.977834, 4.980072, 4.981319, 4.981205, 4.979434, 4.975549, 
    4.969117, 4.959093, 4.944644, 4.928452, 4.909022, 4.887101, 4.86384, 
    4.840705, 4.81933, 4.801309, 4.787976, 4.780247, 4.778527, 4.782729, 
    4.792338, 4.806513, 4.824186, 4.844155, 4.865149, 4.885897, 4.905189, 
    4.921952,
  // momentumY(18,14, 0-49)
    4.886841, 4.883399, 4.882051, 4.882535, 4.884551, 4.887797, 4.891985, 
    4.896872, 4.902257, 4.907996, 4.914003, 4.920245, 4.926744, 4.933584, 
    4.940909, 4.94667, 4.949551, 4.95581, 4.961526, 4.966652, 4.971175, 
    4.976239, 4.979972, 4.982547, 4.984378, 4.98511, 4.984487, 4.982019, 
    4.977257, 4.968933, 4.956161, 4.94096, 4.922206, 4.900504, 4.876897, 
    4.852814, 4.829932, 4.809971, 4.794442, 4.784451, 4.780582, 4.782882, 
    4.790926, 4.803923, 4.820827, 4.840441, 4.861489, 4.882676, 4.90276, 
    4.920603,
  // momentumY(18,15, 0-49)
    4.883207, 4.880651, 4.880136, 4.881371, 4.884029, 4.887794, 4.892372, 
    4.897519, 4.903045, 4.908817, 4.914763, 4.920861, 4.927134, 4.93365, 
    4.940502, 4.948238, 4.950455, 4.956568, 4.962499, 4.96802, 4.973034, 
    4.978105, 4.982003, 4.984821, 4.987122, 4.988574, 4.988962, 4.987782, 
    4.984583, 4.977922, 4.966918, 4.952744, 4.934793, 4.913519, 4.889838, 
    4.865107, 4.84101, 4.819353, 4.801796, 4.789631, 4.783615, 4.783937, 
    4.790273, 4.801894, 4.817789, 4.836773, 4.857575, 4.878895, 4.899468, 
    4.918118,
  // momentumY(18,16, 0-49)
    4.879242, 4.87754, 4.87785, 4.879844, 4.883172, 4.887492, 4.892501, 
    4.897952, 4.903658, 4.909498, 4.915406, 4.921362, 4.92738, 4.933488, 
    4.939705, 4.949776, 4.951613, 4.95754, 4.963687, 4.969635, 4.975175, 
    4.98018, 4.984186, 4.987179, 4.989842, 4.991875, 4.993103, 4.993021, 
    4.991203, 4.986084, 4.976843, 4.963641, 4.946527, 4.925811, 4.902266, 
    4.877148, 4.852115, 4.829021, 4.809649, 4.795449, 4.787349, 4.785682, 
    4.790234, 4.800347, 4.815056, 4.8332, 4.853517, 4.874714, 4.895517, 
    4.914725,
  // momentumY(18,17, 0-49)
    4.875041, 4.874127, 4.875218, 4.87795, 4.881939, 4.886819, 4.892274, 
    4.898053, 4.903974, 4.909922, 4.915837, 4.921696, 4.927484, 4.933181, 
    4.938707, 4.951196, 4.952917, 4.958723, 4.965165, 4.971624, 4.977774, 
    4.982686, 4.986784, 4.989913, 4.992849, 4.995311, 4.997171, 4.997947, 
    4.997252, 4.993465, 4.9859, 4.973534, 4.95721, 4.937099, 4.913828, 
    4.888538, 4.862826, 4.838557, 4.817604, 4.801552, 4.791484, 4.787878, 
    4.790633, 4.799174, 4.812584, 4.829738, 4.849395, 4.870271, 4.891096, 
    4.910655,
  // momentumY(18,18, 0-49)
    4.870688, 4.87046, 4.872247, 4.875643, 4.880235, 4.885635, 4.891515, 
    4.897624, 4.90379, 4.909906, 4.91592, 4.921796, 4.927487, 4.932893, 
    4.937829, 4.952391, 4.954152, 4.960028, 4.966936, 4.974069, 4.980973, 
    4.985815, 4.99005, 4.993322, 4.99646, 4.999198, 5.001451, 5.002779, 
    5.002877, 5.000129, 4.994055, 4.982319, 4.966665, 4.947137, 4.924218, 
    4.898921, 4.872756, 4.847573, 4.825289, 4.807601, 4.795727, 4.790283, 
    4.791286, 4.798248, 4.810311, 4.826389, 4.84527, 4.865687, 4.886379, 
    4.906126,
  // momentumY(18,19, 0-49)
    4.86625, 4.86655, 4.868883, 4.872808, 4.877879, 4.883698, 4.889936, 
    4.896357, 4.902807, 4.909202, 4.915492, 4.921624, 4.927492, 4.932897, 
    4.937518, 4.953274, 4.955041, 4.961284, 4.968928, 4.976991, 4.984876, 
    4.989754, 4.994244, 4.997727, 5.001033, 5.003887, 5.006248, 5.007756, 
    5.008227, 5.006122, 5.001248, 4.98988, 4.974717, 4.955695, 4.933158, 
    4.907983, 4.881572, 4.855722, 4.832371, 4.813286, 4.799805, 4.792671, 
    4.792016, 4.797443, 4.808165, 4.823141, 4.841189, 4.861065, 4.881521, 
    4.901341,
  // momentumY(18,20, 0-49)
    4.862615, 4.864183, 4.867981, 4.873559, 4.880429, 4.888097, 4.896105, 
    4.904039, 4.91155, 4.918352, 4.924236, 4.929071, 4.932817, 4.935514, 
    4.937287, 0, 4.967083, 4.970193, 4.974487, 4.979447, 4.9848, 4.986744, 
    4.989418, 4.992031, 4.995424, 4.999174, 5.003032, 5.006403, 5.008925, 
    5.008933, 5.006418, 4.996209, 4.982046, 4.963815, 4.941799, 4.916811, 
    4.8902, 4.86374, 4.83939, 4.818989, 4.803974, 4.79521, 4.792936, 
    4.796848, 4.806228, 4.820079, 4.837255, 4.856534, 4.87668, 4.896485,
  // momentumY(18,21, 0-49)
    4.858526, 4.860593, 4.864909, 4.870983, 4.878288, 4.886311, 4.89458, 
    4.902694, 4.910328, 4.917231, 4.923228, 4.928211, 4.932137, 4.935033, 
    4.936998, 0, 4.96749, 4.971151, 4.976059, 4.981626, 4.987492, 4.988534, 
    4.990527, 4.992525, 4.995533, 4.999171, 5.003212, 5.007048, 5.010316, 
    5.011328, 5.010325, 5.000771, 4.987464, 4.970185, 4.949078, 4.924807, 
    4.898589, 4.872103, 4.847268, 4.82596, 4.809701, 4.799472, 4.795639, 
    4.798006, 4.805933, 4.818489, 4.834568, 4.852976, 4.872499, 4.891943,
  // momentumY(18,22, 0-49)
    4.854605, 4.857058, 4.861805, 4.868328, 4.876069, 4.884493, 4.893115, 
    4.901526, 4.909408, 4.916522, 4.922707, 4.927864, 4.931949, 4.93498, 
    4.937038, 0, 4.968196, 4.972306, 4.977769, 4.98394, 4.990365, 4.990649, 
    4.992125, 4.993677, 4.996429, 5.000011, 5.004191, 5.008338, 5.01208, 
    5.013722, 5.013745, 5.004387, 4.991473, 4.974729, 4.954206, 4.930459, 
    4.904589, 4.878174, 4.853073, 4.831153, 4.813982, 4.802622, 4.797538, 
    4.798625, 4.805327, 4.816769, 4.831888, 4.849522, 4.86848, 4.887581,
  // momentumY(18,23, 0-49)
    4.850917, 4.853661, 4.858761, 4.865675, 4.873829, 4.882668, 4.891686, 
    4.900468, 4.908682, 4.916094, 4.922538, 4.927917, 4.932185, 4.935344, 
    4.93747, 0, 4.969583, 4.973991, 4.979832, 4.98642, 4.993236, 4.992826, 
    4.993824, 4.99496, 4.99745, 5.000928, 5.005152, 5.009469, 5.013495, 
    5.015525, 5.016229, 5.006853, 4.994095, 4.977653, 4.95752, 4.934175, 
    4.908624, 4.882356, 4.857164, 4.834885, 4.817104, 4.804931, 4.798903, 
    4.798989, 4.804698, 4.81521, 4.8295, 4.846437, 4.864852, 4.883585,
  // momentumY(18,24, 0-49)
    4.847519, 4.850479, 4.85586, 4.863112, 4.871647, 4.880895, 4.890332, 
    4.899526, 4.908134, 4.915905, 4.92267, 4.928324, 4.932813, 4.936135, 
    4.938357, 0, 4.971826, 4.976392, 4.982431, 4.989242, 4.996271, 4.995375, 
    4.996037, 4.996878, 4.999168, 5.002536, 5.006739, 5.011106, 5.015255, 
    5.017463, 5.018531, 5.009044, 4.996279, 4.979924, 4.959941, 4.936765, 
    4.911347, 4.885115, 4.859817, 4.837259, 4.819028, 4.806264, 4.799543, 
    4.798884, 4.803843, 4.813639, 4.827281, 4.843661, 4.86163, 4.880041,
  // momentumY(18,25, 0-49)
    4.84447, 4.847589, 4.853196, 4.860741, 4.869628, 4.879272, 4.889136, 
    4.898769, 4.907809, 4.915988, 4.923122, 4.929097, 4.933853, 4.937385, 
    4.939763, 0, 4.974479, 4.979081, 4.985147, 4.991983, 4.999034, 4.997939, 
    4.99846, 4.999179, 5.001375, 5.00467, 5.008821, 5.013151, 5.017279, 
    5.019472, 5.020578, 5.010951, 4.998077, 4.981641, 4.961603, 4.938382, 
    4.91291, 4.88659, 4.861147, 4.838369, 4.819839, 4.806698, 4.799538, 
    4.7984, 4.802862, 4.81217, 4.825348, 4.841312, 4.858924, 4.877048,
  // momentumY(18,26, 0-49)
    4.841846, 4.845082, 4.850876, 4.858679, 4.867893, 4.877924, 4.888223, 
    4.898314, 4.907815, 4.916437, 4.923976, 4.930305, 4.935359, 4.939139, 
    4.941726, 0, 4.977385, 4.981901, 4.98783, 4.994493, 5.001371, 5.000391, 
    5.000994, 5.001788, 5.004019, 5.007303, 5.01139, 5.015614, 5.019589, 
    5.021584, 5.022406, 5.012643, 4.999584, 4.982924, 4.962636, 4.939158, 
    4.913439, 4.886895, 4.861254, 4.838302, 4.819606, 4.806296, 4.798949, 
    4.797599, 4.801824, 4.810872, 4.823782, 4.839473, 4.856821, 4.874699,
  // momentumY(18,27, 0-49)
    4.839744, 4.843068, 4.84902, 4.857059, 4.866587, 4.877005, 4.887747, 
    4.898317, 4.908307, 4.917399, 4.925366, 4.932062, 4.937419, 4.941448, 
    4.944248, 0, 4.980576, 4.984866, 4.990472, 4.996755, 5.003257, 5.002659, 
    5.003529, 5.004568, 5.006943, 5.01026, 5.014267, 5.018305, 5.021995, 
    5.023608, 5.023826, 5.013915, 5.000586, 4.983556, 4.962839, 4.938921, 
    4.912803, 4.885948, 4.860112, 4.837081, 4.818402, 4.805168, 4.797915, 
    4.796639, 4.800896, 4.809918, 4.822744, 4.838297, 4.855458, 4.873108,
  // momentumY(18,28, 0-49)
    4.838279, 4.841671, 4.847761, 4.856022, 4.86586, 4.876674, 4.887884, 
    4.898968, 4.909482, 4.919071, 4.927473, 4.934519, 4.940135, 4.94435, 
    4.94729, 0, 4.984393, 4.988278, 4.993347, 4.999027, 5.004954, 5.004905, 
    5.006158, 5.007552, 5.010141, 5.013506, 5.017393, 5.021155, 5.024417, 
    5.025462, 5.024777, 5.014656, 5.000932, 4.983361, 4.962024, 4.937493, 
    4.910855, 4.883649, 4.857671, 4.834711, 4.816276, 4.803395, 4.796536, 
    4.795633, 4.800196, 4.80943, 4.82236, 4.837905, 4.854949, 4.872379,
  // momentumY(18,29, 0-49)
    4.837578, 4.841016, 4.847223, 4.855696, 4.865859, 4.8771, 4.888828, 
    4.900484, 4.911574, 4.921689, 4.930514, 4.937848, 4.943614, 4.94786, 
    4.950751, 0, 4.988549, 4.991818, 4.996123, 5.000973, 5.006124, 5.006631, 
    5.00827, 5.010037, 5.012847, 5.016247, 5.019962, 5.023355, 5.02604, 
    5.026312, 5.024417, 5.013925, 4.999619, 4.981328, 4.959243, 4.93405, 
    4.906947, 4.879553, 4.853701, 4.831154, 4.813352, 4.801226, 4.795144, 
    4.794957, 4.800112, 4.80978, 4.822963, 4.83858, 4.855508, 4.872646,
  // momentumY(18,30, 0-49)
    4.837201, 4.839952, 4.84534, 4.852841, 4.861905, 4.872, 4.882656, 
    4.893489, 4.904216, 4.914642, 4.924639, 4.934104, 4.942914, 4.950874, 
    4.957664, 4.980512, 4.978384, 4.985451, 4.993881, 5.002621, 5.011064, 
    5.015289, 5.019503, 5.022801, 5.026014, 5.028763, 5.03095, 5.032186, 
    5.032328, 5.02988, 5.02498, 5.012665, 4.996644, 4.97683, 4.95351, 
    4.927465, 4.899968, 4.872666, 4.847361, 4.825732, 4.809091, 4.798231, 
    4.793395, 4.794331, 4.800419, 4.81079, 4.824425, 4.840233, 4.8571, 
    4.873925,
  // momentumY(18,31, 0-49)
    4.838711, 4.841673, 4.847275, 4.855004, 4.864307, 4.874646, 4.885531, 
    4.896559, 4.907419, 4.917896, 4.927857, 4.937228, 4.945951, 4.953948, 
    4.961065, 4.980995, 4.980417, 4.987096, 4.994756, 5.002519, 5.00993, 
    5.014159, 5.018117, 5.021186, 5.024208, 5.026828, 5.028913, 5.029993, 
    5.029801, 5.02675, 5.020671, 5.008065, 4.991631, 4.971384, 4.94774, 
    4.9216, 4.89433, 4.86762, 4.843251, 4.822825, 4.807539, 4.798059, 
    4.794508, 4.796546, 4.803485, 4.814416, 4.828295, 4.844025, 4.860487, 
    4.876597,
  // momentumY(18,32, 0-49)
    4.841342, 4.844412, 4.850084, 4.857855, 4.867183, 4.877531, 4.888418, 
    4.899436, 4.910273, 4.920713, 4.930632, 4.93998, 4.948754, 4.956964, 
    4.964594, 4.980965, 4.981505, 4.988069, 4.995195, 5.002202, 5.00878, 
    5.013144, 5.016983, 5.019907, 5.02272, 5.025066, 5.026776, 5.02734, 
    5.026409, 5.022374, 5.014822, 5.001704, 4.984722, 4.964009, 4.940114, 
    4.914057, 4.88728, 4.861488, 4.838411, 4.819547, 4.80595, 4.798151, 
    4.796151, 4.799515, 4.807491, 4.819123, 4.833344, 4.849035, 4.865076, 
    4.880392,
  // momentumY(18,33, 0-49)
    4.845201, 4.848296, 4.853919, 4.861576, 4.870737, 4.880888, 4.891561, 
    4.902365, 4.912999, 4.923262, 4.933043, 4.942318, 4.951126, 4.959552, 
    4.967697, 4.980441, 4.981912, 4.988523, 4.995258, 5.001646, 5.007523, 
    5.012081, 5.015876, 5.018697, 5.021259, 5.023195, 5.024305, 5.02406, 
    5.022061, 5.016749, 5.007536, 4.993733, 4.976113, 4.954939, 4.930896, 
    4.905118, 4.879101, 4.85454, 4.833084, 4.816096, 4.804484, 4.798627, 
    4.798405, 4.803288, 4.812459, 4.824915, 4.839553, 4.855231, 4.870821, 
    4.885258,
  // momentumY(18,34, 0-49)
    4.850313, 4.853356, 4.858818, 4.866215, 4.875041, 4.884804, 4.895066, 
    4.905462, 4.915716, 4.925641, 4.935148, 4.944232, 4.952967, 4.961494, 
    4.970001, 4.979457, 4.981847, 4.98854, 4.994935, 5.000776, 5.006025, 
    5.010772, 5.014541, 5.01726, 5.019513, 5.020917, 5.02124, 5.019953, 
    5.016633, 5.00984, 4.998881, 4.98429, 4.966008, 4.944437, 4.920403, 
    4.895131, 4.870153, 4.847122, 4.82758, 4.812739, 4.803346, 4.799632, 
    4.801355, 4.8079, 4.818378, 4.831736, 4.846831, 4.862496, 4.877587, 
    4.891049,
  // momentumY(18,35, 0-49)
    4.85662, 4.859527, 4.864711, 4.871711, 4.880044, 4.889249, 4.898926, 
    4.908741, 4.918445, 4.927876, 4.936965, 4.94572, 4.954232, 4.962675, 
    4.971297, 4.978046, 4.981433, 4.988136, 4.99417, 4.999484, 5.004143, 
    5.009024, 5.012743, 5.015333, 5.017207, 5.017971, 5.017355, 5.014852, 
    5.01003, 5.001642, 4.988949, 4.973538, 4.954648, 4.932821, 4.909005, 
    4.884502, 4.860847, 4.839624, 4.822244, 4.809759, 4.80275, 4.801305, 
    4.805072, 4.813345, 4.825176, 4.839457, 4.855005, 4.870616, 4.885136, 
    4.89752,
  // momentumY(18,36, 0-49)
    4.863973, 4.866647, 4.871443, 4.877914, 4.885613, 4.894113, 4.903052, 
    4.912133, 4.921141, 4.929941, 4.938475, 4.946762, 4.954895, 4.963057, 
    4.971507, 4.97621, 4.980695, 4.987263, 4.992869, 4.997642, 5.001723, 
    5.006649, 5.010259, 5.012672, 5.014094, 5.014126, 5.01246, 5.008624, 
    5.0022, 4.992191, 4.977875, 4.961699, 4.942339, 4.920467, 4.897135, 
    4.87369, 4.85164, 4.83247, 4.817447, 4.807454, 4.802914, 4.80378, 
    4.809597, 4.819584, 4.832732, 4.847884, 4.863813, 4.879286, 4.893135, 
    4.904335,
  // momentumY(18,37, 0-49)
    4.872146, 4.874485, 4.878777, 4.884603, 4.891544, 4.899216, 4.907293, 
    4.91552, 4.923715, 4.931767, 4.939631, 4.947328, 4.954942, 4.962633, 
    4.970646, 4.973928, 4.979574, 4.985822, 4.990914, 4.995116, 4.99861, 
    5.003463, 5.006887, 5.00906, 5.009962, 5.009189, 5.006405, 5.001185, 
    4.993144, 4.981586, 4.965855, 4.949062, 4.929453, 4.907815, 4.885276, 
    4.863191, 4.843011, 4.8261, 4.813562, 4.806119, 4.804044, 4.807168, 
    4.814948, 4.826537, 4.840876, 4.856761, 4.872931, 4.888124, 4.901169, 
    4.911073,
  // momentumY(18,38, 0-49)
    4.880842, 4.882741, 4.886423, 4.891498, 4.897586, 4.904336, 4.911465, 
    4.918751, 4.926048, 4.933264, 4.940367, 4.947376, 4.954354, 4.961426, 
    4.968778, 4.971156, 4.977955, 4.983696, 4.988179, 4.991767, 4.994656, 
    4.999306, 5.002451, 5.004314, 5.004631, 5.003013, 4.999096, 4.992517, 
    4.982934, 4.969998, 4.953146, 4.935975, 4.916419, 4.895351, 4.873941, 
    4.853517, 4.83544, 4.820933, 4.810941, 4.806021, 4.806313, 4.811546, 
    4.821102, 4.834083, 4.849388, 4.86578, 4.881971, 4.896688, 4.908768, 
    4.917272,
  // momentumY(18,39, 0-49)
    4.889717, 4.891066, 4.894044, 4.898291, 4.903454, 4.909225, 4.915352, 
    4.921652, 4.927999, 4.934326, 4.940608, 4.946858, 4.953117, 4.959458, 
    4.965996, 4.96784, 4.975702, 4.980766, 4.984552, 4.987484, 4.989732, 
    4.99404, 4.996809, 4.998293, 4.997983, 4.995514, 4.990504, 4.982667, 
    4.971714, 4.957668, 4.940073, 4.922842, 4.903699, 4.883575, 4.863635, 
    4.84515, 4.829363, 4.817347, 4.809879, 4.807374, 4.809848, 4.816947, 
    4.827996, 4.842059, 4.858009, 4.874594, 4.890515, 4.904504, 4.915439, 
    4.922453,
  // momentumY(18,40, 0-49)
    4.8984, 4.899097, 4.90129, 4.904646, 4.908849, 4.913617, 4.91873, 
    4.924032, 4.929419, 4.934838, 4.940274, 4.945725, 4.951211, 4.956755, 
    4.96239, 4.963936, 4.972683, 4.976931, 4.979949, 4.982178, 4.983747, 
    4.987577, 4.989875, 4.990921, 4.989964, 4.98668, 4.98068, 4.971765, 
    4.959704, 4.944898, 4.927004, 4.910091, 4.891764, 4.872965, 4.854824, 
    4.838517, 4.825151, 4.815638, 4.810602, 4.81032, 4.814709, 4.823346, 
    4.835516, 4.850266, 4.866456, 4.882841, 4.898137, 4.911113, 4.920713, 
    4.926178,
  // momentumY(18,41, 0-49)
    4.906529, 4.906476, 4.907814, 4.910242, 4.91347, 4.917244, 4.921369, 
    4.925701, 4.930154, 4.934687, 4.939281, 4.94393, 4.948625, 4.953344, 
    4.958044, 4.959407, 4.968792, 4.97213, 4.974324, 4.975806, 4.976653, 
    4.979882, 4.981626, 4.98219, 4.980597, 4.976579, 4.969752, 4.960011, 
    4.947186, 4.932035, 4.914319, 4.898144, 4.881041, 4.863939, 4.847887, 
    4.833943, 4.823065, 4.816005, 4.813236, 4.814918, 4.820882, 4.830656, 
    4.843504, 4.858468, 4.874428, 4.890163, 4.904439, 4.916101, 4.924196, 
    4.928107,
  // momentumY(18,42, 0-49)
    4.913782, 4.912883, 4.913308, 4.914782, 4.917043, 4.919858, 4.923043, 
    4.926467, 4.93005, 4.933751, 4.937549, 4.941423, 4.945343, 4.949245, 
    4.953024, 4.954234, 4.963964, 4.96634, 4.967675, 4.96837, 4.968452, 
    4.970979, 4.972106, 4.972164, 4.969982, 4.965353, 4.957918, 4.947659, 
    4.934467, 4.919428, 4.902383, 4.887368, 4.871888, 4.856811, 4.843086, 
    4.831631, 4.823244, 4.818518, 4.817794, 4.821123, 4.82827, 4.83873, 
    4.851759, 4.866421, 4.881636, 4.896245, 4.9091, 4.919161, 4.925624, 
    4.928048,
  // momentumY(18,43, 0-49)
    4.919908, 4.918075, 4.917529, 4.918031, 4.919343, 4.921244, 4.923561, 
    4.926164, 4.928969, 4.931925, 4.934999, 4.938159, 4.941349, 4.944471, 
    4.947376, 4.948405, 4.958177, 4.959578, 4.960035, 4.959912, 4.959199, 
    4.960948, 4.961421, 4.960978, 4.958283, 4.953208, 4.945422, 4.934996, 
    4.921866, 4.907401, 4.8915, 4.878047, 4.864542, 4.851766, 4.840542, 
    4.831635, 4.82568, 4.823121, 4.824172, 4.828796, 4.8367, 4.847362, 
    4.860054, 4.873881, 4.887831, 4.900847, 4.911908, 4.920138, 4.924921, 
    4.926015,
  // momentumY(18,44, 0-49)
    4.924776, 4.921913, 4.92034, 4.91985, 4.920226, 4.921264, 4.92279, 
    4.924667, 4.926798, 4.929115, 4.931567, 4.934095, 4.936621, 4.939024, 
    4.941122, 4.941914, 4.951438, 4.951888, 4.951467, 4.95051, 4.94899, 
    4.94992, 4.94973, 4.948813, 4.945714, 4.940386, 4.932531, 4.9223, 
    4.909667, 4.896218, 4.881884, 4.870344, 4.859107, 4.848838, 4.840219, 
    4.833856, 4.830224, 4.829626, 4.832157, 4.837701, 4.845929, 4.856311, 
    4.868156, 4.880635, 4.89284, 4.903851, 4.912822, 4.91908, 4.922236, 
    4.922259,
  // momentumY(18,45, 0-49)
    4.928407, 4.924418, 4.921751, 4.920234, 4.919677, 4.919885, 4.920683, 
    4.921923, 4.923484, 4.925271, 4.927204, 4.929194, 4.931141, 4.932897, 
    4.934264, 4.934757, 4.943786, 4.943328, 4.942047, 4.94026, 4.937941, 
    4.93805, 4.937223, 4.935887, 4.932515, 4.927137, 4.9195, 4.909817, 
    4.898086, 4.886047, 4.873634, 4.864293, 4.855537, 4.847908, 4.841933, 
    4.838057, 4.836599, 4.837729, 4.841436, 4.847537, 4.855672, 4.865327, 
    4.875862, 4.886545, 4.896604, 4.9053, 4.912002, 4.916276, 4.917975, 
    4.917284,
  // momentumY(18,46, 0-49)
    4.931002, 4.925789, 4.921949, 4.919353, 4.917837, 4.917222, 4.917328, 
    4.917989, 4.919061, 4.920411, 4.921917, 4.92346, 4.924904, 4.926087, 
    4.926797, 4.926932, 4.935273, 4.933967, 4.931861, 4.929269, 4.926188, 
    4.925509, 4.924102, 4.922422, 4.918921, 4.9137, 4.906552, 4.897737, 
    4.887263, 4.876956, 4.866735, 4.859797, 4.853657, 4.848723, 4.845367, 
    4.843875, 4.844419, 4.84704, 4.851633, 4.857956, 4.865634, 4.87418, 
    4.883031, 4.891579, 4.899223, 4.905437, 4.90984, 4.912262, 4.912797, 
    4.911825,
  // momentumY(18,47, 0-49)
    4.932955, 4.926421, 4.921322, 4.91757, 4.91504, 4.913567, 4.912973, 
    4.913074, 4.91369, 4.914652, 4.915792, 4.916949, 4.917954, 4.91862, 
    4.918736, 4.91845, 4.925973, 4.923887, 4.921003, 4.917657, 4.913873, 
    4.912481, 4.910572, 4.908642, 4.905159, 4.900286, 4.893863, 4.88618, 
    4.877249, 4.868914, 4.861065, 4.856644, 4.853178, 4.850926, 4.850114, 
    4.850874, 4.853234, 4.85712, 4.862342, 4.86861, 4.875546, 4.88271, 
    4.88963, 4.895852, 4.900975, 4.904717, 4.906961, 4.907805, 4.907571, 
    4.906791,
  // momentumY(18,48, 0-49)
    4.934845, 4.9269, 4.920446, 4.915445, 4.911812, 4.909406, 4.908049, 
    4.907547, 4.907685, 4.908252, 4.909031, 4.909818, 4.910404, 4.910583, 
    4.91014, 4.909373, 4.916004, 4.9132, 4.909599, 4.905562, 4.90116, 
    4.899149, 4.896842, 4.894763, 4.891435, 4.887076, 4.881566, 4.875215, 
    4.868028, 4.861816, 4.856431, 4.854557, 4.85374, 4.854105, 4.855721, 
    4.858578, 4.862577, 4.867533, 4.873183, 4.879201, 4.885219, 4.890858, 
    4.895762, 4.899647, 4.902333, 4.903794, 4.904185, 4.903849, 4.903304, 
    4.90318,
  // momentumY(18,49, 0-49)
    4.943079, 4.933022, 4.92444, 4.917368, 4.911783, 4.907586, 4.904629, 
    4.902708, 4.901586, 4.901, 4.900681, 4.900353, 4.899747, 4.898587, 
    4.896599, 4.894702, 4.907625, 4.902482, 4.896469, 4.890329, 4.884231, 
    4.883526, 4.882961, 4.883486, 4.882074, 4.87913, 4.874318, 4.868094, 
    4.860242, 4.854196, 4.849467, 4.851037, 4.85378, 4.857646, 4.86253, 
    4.868235, 4.874485, 4.880953, 4.887276, 4.893087, 4.898046, 4.901875, 
    4.904406, 4.905601, 4.905601, 4.904716, 4.90344, 4.902396, 4.902278, 
    4.903772,
  // momentumY(19,0, 0-49)
    4.863467, 4.857262, 4.854007, 4.853439, 4.855211, 4.858918, 4.86413, 
    4.870421, 4.877393, 4.884692, 4.892019, 4.899126, 4.905809, 4.911901, 
    4.917256, 4.921696, 4.926414, 4.929109, 4.930936, 4.931877, 4.931879, 
    4.93122, 4.92947, 4.92665, 4.922586, 4.917221, 4.910484, 4.902398, 
    4.893026, 4.882643, 4.871445, 4.860118, 4.848811, 4.838039, 4.828342, 
    4.820229, 4.814119, 4.8103, 4.808887, 4.80981, 4.812818, 4.817494, 
    4.823306, 4.829645, 4.835906, 4.841548, 4.846171, 4.849586, 4.85186, 
    4.853332,
  // momentumY(19,1, 0-49)
    4.865608, 4.859947, 4.857208, 4.857111, 4.8593, 4.863361, 4.868865, 
    4.875392, 4.882556, 4.890017, 4.897492, 4.904748, 4.911586, 4.917842, 
    4.923354, 4.927824, 4.933651, 4.936447, 4.938407, 4.939521, 4.939701, 
    4.939492, 4.938069, 4.935489, 4.931462, 4.925898, 4.918675, 4.909807, 
    4.899339, 4.887649, 4.874897, 4.862156, 4.849326, 4.837008, 4.825834, 
    4.816401, 4.809213, 4.804626, 4.802801, 4.803697, 4.807059, 4.812455, 
    4.8193, 4.826921, 4.834619, 4.841738, 4.847753, 4.85234, 4.855436, 
    4.857277,
  // momentumY(19,2, 0-49)
    4.868079, 4.86294, 4.86067, 4.86098, 4.863502, 4.867823, 4.873523, 
    4.880189, 4.887453, 4.894991, 4.90254, 4.909874, 4.91681, 4.923179, 
    4.928813, 4.933246, 4.940066, 4.942986, 4.945104, 4.946426, 4.946843, 
    4.947165, 4.946175, 4.943969, 4.940157, 4.934615, 4.927167, 4.917808, 
    4.90655, 4.893838, 4.879786, 4.865834, 4.851622, 4.837819, 4.825143, 
    4.814283, 4.805833, 4.800229, 4.7977, 4.798252, 4.801656, 4.807476, 
    4.815114, 4.823852, 4.832918, 4.841565, 4.849153, 4.855217, 4.859553, 
    4.862253,
  // momentumY(19,3, 0-49)
    4.870552, 4.86591, 4.864064, 4.864718, 4.867503, 4.872014, 4.877833, 
    4.884569, 4.891868, 4.899426, 4.906993, 4.914361, 4.921353, 4.927806, 
    4.93355, 4.937875, 4.945512, 4.948591, 4.950888, 4.952444, 4.953139, 
    4.954044, 4.953572, 4.95185, 4.948418, 4.943113, 4.935712, 4.926178, 
    4.914483, 4.901093, 4.886057, 4.871165, 4.855776, 4.840611, 4.826462, 
    4.814105, 4.804229, 4.797366, 4.793829, 4.793693, 4.796775, 4.802673, 
    4.810785, 4.820376, 4.830633, 4.840738, 4.84995, 4.857678, 4.863564, 
    4.867543,
  // momentumY(19,4, 0-49)
    4.872817, 4.868643, 4.867184, 4.868135, 4.871129, 4.875768, 4.881651, 
    4.888405, 4.895691, 4.903227, 4.910775, 4.918141, 4.92516, 4.931677, 
    4.937528, 4.941673, 4.949905, 4.953179, 4.955673, 4.957477, 4.958472, 
    4.959987, 4.960082, 4.958926, 4.956011, 4.951143, 4.944056, 4.934675, 
    4.922916, 4.909231, 4.893579, 4.878071, 4.861773, 4.845433, 4.829899, 
    4.816028, 4.804605, 4.796266, 4.79143, 4.790257, 4.792642, 4.798227, 
    4.806442, 4.816557, 4.827739, 4.839124, 4.849892, 4.859341, 4.866971, 
    4.872547,
  // momentumY(19,5, 0-49)
    4.874774, 4.871048, 4.869942, 4.871148, 4.874307, 4.879029, 4.884934, 
    4.891664, 4.898901, 4.906378, 4.913873, 4.921207, 4.928225, 4.93479, 
    4.940752, 4.944649, 4.953211, 4.956712, 4.959419, 4.961472, 4.962777, 
    4.964893, 4.965576, 4.96503, 4.962738, 4.958478, 4.951951, 4.943034, 
    4.931594, 4.918012, 4.902144, 4.886379, 4.869491, 4.852226, 4.835463, 
    4.820125, 4.807089, 4.797104, 4.790708, 4.788169, 4.789482, 4.79436, 
    4.802285, 4.812552, 4.824332, 4.836738, 4.848891, 4.860003, 4.869445, 
    4.876825,
  // momentumY(19,6, 0-49)
    4.876401, 4.873109, 4.872334, 4.873767, 4.877055, 4.881827, 4.887718, 
    4.894387, 4.901539, 4.90892, 4.916327, 4.923593, 4.930583, 4.937176, 
    4.943255, 4.946844, 4.955447, 4.959205, 4.962132, 4.964428, 4.966038, 
    4.968722, 4.969982, 4.970057, 4.968456, 4.964935, 4.959171, 4.951004, 
    4.94024, 4.92715, 4.911473, 4.895832, 4.878706, 4.860817, 4.843043, 
    4.826352, 4.811706, 4.799966, 4.7918, 4.78761, 4.787505, 4.791297, 
    4.798542, 4.808578, 4.820599, 4.833713, 4.847009, 4.85963, 4.870845, 
    4.880115,
  // momentumY(19,7, 0-49)
    4.877742, 4.87488, 4.87442, 4.876059, 4.879453, 4.884243, 4.890086, 
    4.896661, 4.903688, 4.910936, 4.918213, 4.925372, 4.932297, 4.938896, 
    4.945095, 4.948344, 4.956688, 4.960714, 4.963864, 4.966398, 4.968299, 
    4.971492, 4.973291, 4.973963, 4.973082, 4.970386, 4.965547, 4.958364, 
    4.94859, 4.936349, 4.921254, 4.906102, 4.889108, 4.870925, 4.852411, 
    4.83455, 4.818367, 4.804838, 4.79476, 4.78869, 4.78687, 4.789238, 
    4.795435, 4.80487, 4.816771, 4.830261, 4.844414, 4.858326, 4.871181, 
    4.882321,
  // momentumY(19,8, 0-49)
    4.878867, 4.876438, 4.876289, 4.878121, 4.881602, 4.886387, 4.892151, 
    4.898596, 4.90546, 4.912529, 4.919632, 4.926641, 4.93346, 4.940037, 
    4.946343, 4.94926, 4.957064, 4.961346, 4.964719, 4.967476, 4.969651, 
    4.973279, 4.975556, 4.976775, 4.976603, 4.974774, 4.970967, 4.964946, 
    4.956418, 4.94533, 4.931167, 4.916834, 4.900319, 4.88219, 4.863243, 
    4.844447, 4.826875, 4.811594, 4.799544, 4.791435, 4.787673, 4.788329, 
    4.793161, 4.801657, 4.813101, 4.826638, 4.841345, 4.856289, 4.87059, 
    4.883487,
  // momentumY(19,9, 0-49)
    4.879853, 4.877869, 4.878036, 4.880059, 4.883614, 4.888375, 4.894034, 
    4.900314, 4.906975, 4.913821, 4.920701, 4.927508, 4.934181, 4.940696, 
    4.94708, 4.94973, 4.956745, 4.961252, 4.964836, 4.967809, 4.970237, 
    4.974212, 4.976891, 4.978584, 4.979081, 4.978118, 4.975397, 4.970651, 
    4.963554, 4.953855, 4.940918, 4.927673, 4.911951, 4.894206, 4.875144, 
    4.855691, 4.836935, 4.820017, 4.80601, 4.795788, 4.789926, 4.788655, 
    4.791863, 4.799135, 4.809819, 4.823099, 4.838062, 4.853761, 4.86927, 
    4.883741,
  // momentumY(19,10, 0-49)
    4.880766, 4.879248, 4.879743, 4.881961, 4.885587, 4.890312, 4.895844, 
    4.901929, 4.90835, 4.91493, 4.921543, 4.928103, 4.934577, 4.940979, 
    4.947385, 4.949909, 4.955944, 4.960614, 4.964392, 4.967567, 4.970238, 
    4.974462, 4.977457, 4.979537, 4.980639, 4.980505, 4.978874, 4.975456, 
    4.969903, 4.961752, 4.950266, 4.938305, 4.923625, 4.906556, 4.887687, 
    4.867873, 4.848182, 4.829807, 4.813938, 4.801608, 4.79357, 4.79023, 
    4.79162, 4.797441, 4.807114, 4.819869, 4.834813, 4.850992, 4.867447, 
    4.883266,
  // momentumY(19,11, 0-49)
    4.881644, 4.880621, 4.881466, 4.883892, 4.887596, 4.892278, 4.897672, 
    4.903541, 4.909692, 4.91597, 4.922273, 4.92854, 4.934764, 4.94099, 
    4.94733, 4.949949, 4.954883, 4.959633, 4.963575, 4.966947, 4.969853, 
    4.974226, 4.977445, 4.979825, 4.981448, 4.982079, 4.9815, 4.979406, 
    4.975439, 4.968922, 4.95904, 4.948476, 4.935015, 4.918853, 4.900454, 
    4.880566, 4.860214, 4.840611, 4.823038, 4.80868, 4.798471, 4.792996, 
    4.792449, 4.796651, 4.805115, 4.817122, 4.8318, 4.8482, 4.865337, 4.882246,
  // momentumY(19,12, 0-49)
    4.882496, 4.881999, 4.883224, 4.885882, 4.889676, 4.894325, 4.899577, 
    4.90522, 4.911082, 4.917034, 4.922996, 4.928931, 4.934853, 4.940827, 
    4.946981, 4.949989, 4.95378, 4.958515, 4.962585, 4.966149, 4.969291, 
    4.973717, 4.977075, 4.979658, 4.981715, 4.983027, 4.983429, 4.982606, 
    4.9802, 4.975337, 4.967144, 4.958006, 4.945863, 4.930773, 4.913065, 
    4.893366, 4.872625, 4.852049, 4.832983, 4.816743, 4.804437, 4.796834, 
    4.794295, 4.796777, 4.803885, 4.814964, 4.829169, 4.845552, 4.863111, 
    4.880845,
  // momentumY(19,13, 0-49)
    4.883292, 4.883357, 4.884997, 4.887918, 4.891829, 4.896464, 4.901587, 
    4.907006, 4.912575, 4.918189, 4.923789, 4.929358, 4.934927, 4.940565, 
    4.94639, 4.950139, 4.952823, 4.957446, 4.961614, 4.96537, 4.968758, 
    4.973145, 4.976562, 4.979265, 4.981663, 4.983564, 4.98485, 4.985204, 
    4.984283, 4.981029, 4.974552, 4.966794, 4.955986, 4.942058, 4.9252, 
    4.905908, 4.885034, 4.863748, 4.84343, 4.825501, 4.811233, 4.801569, 
    4.797047, 4.797762, 4.803423, 4.813437, 4.826993, 4.84315, 4.86089, 
    4.879182,
  // momentumY(19,14, 0-49)
    4.883975, 4.884635, 4.886726, 4.889947, 4.894012, 4.898662, 4.903681, 
    4.908897, 4.914186, 4.919464, 4.924696, 4.929881, 4.935049, 4.940267, 
    4.945613, 4.950459, 4.952142, 4.956577, 4.960824, 4.964785, 4.968439, 
    4.972709, 4.976121, 4.978877, 4.981533, 4.983922, 4.985978, 4.987384, 
    4.98782, 4.986081, 4.981294, 4.974806, 4.965281, 4.952532, 4.936615, 
    4.917893, 4.897106, 4.875359, 4.85404, 4.83465, 4.818594, 4.806993, 
    4.800546, 4.799497, 4.803661, 4.812512, 4.825278, 4.841026, 4.858731, 
    4.877334,
  // momentumY(19,15, 0-49)
    4.884464, 4.885746, 4.888322, 4.891884, 4.896142, 4.900849, 4.905801, 
    4.910846, 4.915881, 4.920848, 4.925724, 4.930517, 4.93526, 4.939989, 
    4.94473, 4.95096, 4.951797, 4.956015, 4.960347, 4.964542, 4.968503, 
    4.972597, 4.97596, 4.978716, 4.981555, 4.984333, 4.987031, 4.989339, 
    4.990971, 4.990606, 4.987436, 4.98206, 4.973706, 4.962089, 4.94714, 
    4.929091, 4.908561, 4.886575, 4.864501, 4.843886, 4.82625, 4.812865, 
    4.804594, 4.801823, 4.804478, 4.812106, 4.823973, 4.83916, 4.856639, 
    4.875334,
  // momentumY(19,16, 0-49)
    4.884663, 4.88658, 4.889668, 4.893605, 4.898099, 4.902907, 4.907837, 
    4.912756, 4.917584, 4.922279, 4.926834, 4.931263, 4.935582, 4.939795, 
    4.943863, 4.951606, 4.951766, 4.955799, 4.960267, 4.964756, 4.969089, 
    4.972967, 4.976264, 4.978997, 4.981962, 4.985034, 4.988237, 4.991272, 
    4.993902, 4.994734, 4.993072, 4.988607, 4.981264, 4.970675, 4.956662, 
    4.93933, 4.919178, 4.897139, 4.874533, 4.85293, 4.833932, 4.818943, 
    4.808976, 4.804556, 4.805722, 4.812094, 4.822984, 4.837489, 4.854583, 
    4.873177,
  // momentumY(19,17, 0-49)
    4.884471, 4.887014, 4.890623, 4.894957, 4.899719, 4.904669, 4.909626, 
    4.914478, 4.919161, 4.923654, 4.92796, 4.932091, 4.936043, 4.939777, 
    4.943196, 4.952326, 4.951941, 4.9559, 4.960605, 4.965496, 4.970294, 
    4.973958, 4.977208, 4.979924, 4.982979, 4.986258, 4.989816, 4.993383, 
    4.996779, 4.998592, 4.998283, 4.994504, 4.987976, 4.978271, 4.96511, 
    4.948489, 4.928789, 4.90684, 4.883897, 4.861527, 4.841388, 4.824988, 
    4.813472, 4.8075, 4.807219, 4.81233, 4.822189, 4.835921, 4.852504, 
    4.870842,
  // momentumY(19,18, 0-49)
    4.883793, 4.886919, 4.891025, 4.895751, 4.900793, 4.905913, 4.910947, 
    4.915798, 4.920425, 4.924825, 4.929009, 4.932978, 4.936702, 4.940094, 
    4.94299, 4.953041, 4.952164, 4.956231, 4.961337, 4.966779, 4.972184, 
    4.975669, 4.978938, 4.981686, 4.984823, 4.988232, 4.991991, 4.995869, 
    4.999767, 5.002297, 5.003136, 4.999793, 4.993859, 4.984858, 4.972429, 
    4.956472, 4.937254, 4.915499, 4.892387, 4.869453, 4.848384, 4.830771, 
    4.817868, 4.810457, 4.808792, 4.812659, 4.821465, 4.834362, 4.850341, 
    4.868311,
  // momentumY(19,19, 0-49)
    4.882538, 4.886151, 4.890681, 4.895749, 4.901048, 4.906345, 4.911496, 
    4.916429, 4.921131, 4.92561, 4.929882, 4.933926, 4.937669, 4.94096, 
    4.943571, 4.95371, 4.952253, 4.956655, 4.962374, 4.968572, 4.974777, 
    4.978183, 4.981593, 4.984472, 4.987724, 4.991202, 4.994999, 4.998935, 
    5.003021, 5.00595, 5.007671, 5.004481, 4.998894, 4.990393, 4.978553, 
    4.963183, 4.944447, 4.922963, 4.899824, 4.876513, 4.854719, 4.836087, 
    4.821965, 4.813243, 4.810278, 4.812939, 4.820692, 4.832723, 4.848042, 
    4.865566,
  // momentumY(19,20, 0-49)
    4.881588, 4.886601, 4.892593, 4.899169, 4.905969, 4.912692, 4.919097, 
    4.924998, 4.930258, 4.934787, 4.938541, 4.941516, 4.943758, 4.94535, 
    4.946416, 0, 4.960864, 4.963375, 4.966852, 4.970822, 4.975077, 4.975944, 
    4.977604, 4.979422, 4.982367, 4.986216, 4.99093, 4.996161, 5.00179, 
    5.006393, 5.010077, 5.007852, 5.003162, 4.995485, 4.98438, 4.969624, 
    4.951338, 4.930086, 4.906902, 4.883231, 4.860764, 4.841182, 4.825912, 
    4.815937, 4.811708, 4.813176, 4.819865, 4.831002, 4.845614, 4.862631,
  // momentumY(19,21, 0-49)
    4.87942, 4.884988, 4.891505, 4.898539, 4.905715, 4.912723, 4.919326, 
    4.92536, 4.930717, 4.935334, 4.939191, 4.942301, 4.944708, 4.946493, 
    4.947779, 0, 4.960035, 4.963074, 4.967126, 4.971672, 4.976431, 4.976584, 
    4.977723, 4.979072, 4.98174, 4.985524, 4.990396, 4.995993, 5.002195, 
    5.007564, 5.012428, 5.010612, 5.006535, 4.999634, 4.989399, 4.975526, 
    4.958041, 4.937399, 4.914538, 4.890834, 4.867946, 4.84758, 4.831234, 
    4.819987, 4.814397, 4.814506, 4.819916, 4.829904, 4.843533, 4.859751,
  // momentumY(19,22, 0-49)
    4.876799, 4.882879, 4.889917, 4.897455, 4.905089, 4.912499, 4.919439, 
    4.925747, 4.931327, 4.936132, 4.940154, 4.943415, 4.945968, 4.947898, 
    4.949335, 0, 4.959913, 4.963387, 4.967949, 4.973043, 4.978314, 4.977839, 
    4.978555, 4.979537, 4.982003, 4.985746, 4.990732, 4.996574, 5.003149, 
    5.009007, 5.014683, 5.012933, 5.009101, 5.002608, 4.992905, 4.97964, 
    4.962763, 4.942643, 4.920128, 4.896511, 4.873403, 4.852501, 4.835343, 
    4.823078, 4.816355, 4.815298, 4.819583, 4.828539, 4.841269, 4.856745,
  // momentumY(19,23, 0-49)
    4.873835, 4.880381, 4.887924, 4.895979, 4.904121, 4.912008, 4.91938, 
    4.926068, 4.931972, 4.937049, 4.941298, 4.944747, 4.947457, 4.949518, 
    4.951072, 0, 4.960715, 4.964478, 4.969381, 4.974841, 4.980453, 4.979389, 
    4.979692, 4.980315, 4.982558, 4.986212, 4.991232, 4.997212, 5.004019, 
    5.010185, 5.016409, 5.014583, 5.010819, 5.004539, 4.995176, 4.982343, 
    4.96594, 4.946269, 4.924097, 4.900642, 4.877457, 4.856218, 4.838474, 
    4.825424, 4.817783, 4.815747, 4.819055, 4.827091, 4.838994, 4.853765,
  // momentumY(19,24, 0-49)
    4.870672, 4.877634, 4.885653, 4.894224, 4.902894, 4.911297, 4.91916, 
    4.926295, 4.932595, 4.93801, 4.94254, 4.946218, 4.949106, 4.951304, 
    4.952971, 0, 4.962595, 4.966502, 4.971569, 4.977206, 4.982986, 4.981498, 
    4.981503, 4.981868, 4.98394, 4.987504, 4.992511, 4.998539, 5.005456, 
    5.011777, 5.018311, 5.016373, 5.012581, 5.006359, 4.997128, 4.984486, 
    4.968306, 4.948847, 4.926829, 4.903417, 4.880123, 4.858602, 4.840403, 
    4.826757, 4.818415, 4.815626, 4.818173, 4.82548, 4.836718, 4.850913,
  // momentumY(19,25, 0-49)
    4.867481, 4.874813, 4.883271, 4.892335, 4.901527, 4.91046, 4.918839, 
    4.926459, 4.933195, 4.938988, 4.943835, 4.947769, 4.950856, 4.953206, 
    4.954986, 0, 4.965112, 4.969028, 4.974089, 4.979712, 4.985476, 4.983797, 
    4.983668, 4.983923, 4.985918, 4.989429, 4.994407, 5.000427, 5.007351, 
    5.013689, 5.020282, 5.018254, 5.014394, 5.008122, 4.998861, 4.986204, 
    4.970013, 4.950536, 4.92847, 4.904962, 4.881504, 4.859735, 4.841204, 
    4.827145, 4.818328, 4.815025, 4.817045, 4.823834, 4.834585, 4.848341,
  // momentumY(19,26, 0-49)
    4.864459, 4.87211, 4.880964, 4.890482, 4.900172, 4.909622, 4.918519, 
    4.926631, 4.933817, 4.940006, 4.945184, 4.949382, 4.952669, 4.955164, 
    4.957052, 0, 4.968115, 4.971904, 4.97679, 4.98221, 4.987775, 4.986162, 
    4.986086, 4.986403, 4.988436, 4.991954, 4.996908, 5.002874, 5.009715, 
    5.015938, 5.022344, 5.020271, 5.016323, 5.009913, 5.00047, 4.98759, 
    4.971152, 4.951414, 4.929086, 4.905328, 4.881636, 4.859649, 4.840906, 
    4.826628, 4.817581, 4.814027, 4.815778, 4.822286, 4.832751, 4.846226,
  // momentumY(19,27, 0-49)
    4.861812, 4.869731, 4.878926, 4.888848, 4.898993, 4.908931, 4.918322, 
    4.926916, 4.934547, 4.941125, 4.946622, 4.951062, 4.954522, 4.957128, 
    4.959073, 0, 4.97163, 4.975142, 4.979673, 4.984694, 4.989872, 4.988544, 
    4.988675, 4.989195, 4.991359, 4.994929, 4.999852, 5.005712, 5.012372, 
    5.018343, 5.024315, 5.022226, 5.018149, 5.011499, 5.001717, 4.988418, 
    4.971513, 4.951303, 4.928545, 4.904437, 4.880499, 4.858378, 4.839594, 
    4.825338, 4.816338, 4.812825, 4.814583, 4.821054, 4.831435, 4.844779,
  // momentumY(19,28, 0-49)
    4.859741, 4.867873, 4.877347, 4.887616, 4.898163, 4.908547, 4.918406, 
    4.927459, 4.935514, 4.942453, 4.948228, 4.952856, 4.956412, 4.959038, 
    4.960937, 0, 4.975993, 4.979054, 4.983034, 4.987453, 4.992063, 4.991148, 
    4.991572, 4.99238, 4.994724, 4.998356, 5.003215, 5.008902, 5.015275, 
    5.020853, 5.026161, 5.024028, 5.019733, 5.012695, 5.002378, 4.988438, 
    4.970845, 4.949972, 4.926649, 4.90214, 4.87801, 4.8559, 4.837305, 
    4.823361, 4.814726, 4.811572, 4.813638, 4.820332, 4.830835, 4.844201,
  // momentumY(19,29, 0-49)
    4.858432, 4.866712, 4.876399, 4.88695, 4.897851, 4.908648, 4.918948, 
    4.92844, 4.936892, 4.944144, 4.950123, 4.95483, 4.958349, 4.960835, 
    4.962511, 0, 4.980938, 4.983357, 4.986584, 4.990198, 4.994048, 4.993536, 
    4.994227, 4.995311, 4.997817, 5.001482, 5.006229, 5.011665, 5.017635, 
    5.022667, 5.027061, 5.024763, 5.020088, 5.012481, 5.00145, 4.986721, 
    4.968343, 4.946784, 4.922968, 4.898229, 4.874156, 4.852381, 4.834337, 
    4.821075, 4.813166, 4.810695, 4.81334, 4.820467, 4.831241, 4.8447,
  // momentumY(19,30, 0-49)
    4.857325, 4.864811, 4.87362, 4.883223, 4.89315, 4.903017, 4.912543, 
    4.921545, 4.929926, 4.937651, 4.944711, 4.951098, 4.956753, 4.961548, 
    4.965257, 4.981699, 4.974598, 4.979191, 4.985151, 4.991585, 4.998013, 
    5.000706, 5.003804, 5.006528, 5.009774, 5.013294, 5.017124, 5.021049, 
    5.02509, 5.027961, 5.029866, 5.026049, 5.019855, 5.010766, 4.998342, 
    4.982376, 4.962988, 4.940724, 4.916574, 4.891904, 4.868294, 4.847318, 
    4.830311, 4.818207, 4.811459, 4.810057, 4.813608, 4.821434, 4.832671, 
    4.846352,
  // momentumY(19,31, 0-49)
    4.858174, 4.865802, 4.874738, 4.884463, 4.894507, 4.904485, 4.9141, 
    4.923157, 4.931543, 4.939215, 4.946176, 4.952444, 4.958014, 4.962843, 
    4.966795, 4.981744, 4.976817, 4.98103, 4.986337, 4.99197, 4.997562, 
    5.000377, 5.003357, 5.005968, 5.009114, 5.01259, 5.016417, 5.020319, 
    5.02421, 5.026711, 5.027736, 5.023791, 5.017277, 5.007711, 4.994723, 
    4.978187, 4.958328, 4.935792, 4.911653, 4.88733, 4.8644, 4.844378, 
    4.828509, 4.817608, 4.812016, 4.811631, 4.815988, 4.824363, 4.835867, 
    4.849523,
  // momentumY(19,32, 0-49)
    4.860078, 4.867659, 4.876506, 4.886116, 4.896039, 4.905897, 4.915404, 
    4.924363, 4.932662, 4.940258, 4.947163, 4.953413, 4.959052, 4.964091, 
    4.968487, 4.981169, 4.978074, 4.982155, 4.987026, 4.992065, 4.997014, 
    5.000091, 5.003103, 5.005722, 5.008819, 5.012202, 5.015869, 5.019507, 
    5.02294, 5.024753, 5.024618, 5.020299, 5.013247, 5.003031, 4.989363, 
    4.972216, 4.95193, 4.929254, 4.905345, 4.881649, 4.859718, 4.840992, 
    4.826592, 4.817206, 4.813052, 4.813928, 4.819293, 4.828377, 4.840262, 
    4.853956,
  // momentumY(19,33, 0-49)
    4.863094, 4.870475, 4.879053, 4.888352, 4.897948, 4.907487, 4.916703, 
    4.925407, 4.9335, 4.940943, 4.947758, 4.953999, 4.959738, 4.965044, 
    4.969951, 4.980079, 4.97859, 4.982728, 4.987326, 4.991925, 4.996374, 
    4.999796, 5.002942, 5.005651, 5.008716, 5.011941, 5.015303, 5.018456, 
    5.021159, 5.022017, 5.020511, 5.015593, 5.007808, 4.996795, 4.982359, 
    4.964593, 4.943953, 4.921297, 4.897847, 4.875063, 4.854445, 4.837331, 
    4.824705, 4.817112, 4.814642, 4.816987, 4.823531, 4.833456, 4.845809, 
    4.859584,
  // momentumY(19,34, 0-49)
    4.867206, 4.874252, 4.882409, 4.891233, 4.900333, 4.909385, 4.918148, 
    4.926455, 4.934219, 4.941414, 4.948065, 4.954243, 4.960041, 4.96557, 
    4.970939, 4.978593, 4.978584, 4.98288, 4.987299, 4.991557, 4.995606, 
    4.999401, 5.002732, 5.005574, 5.008594, 5.011591, 5.014505, 5.016977, 
    5.018713, 5.018397, 5.015368, 5.009659, 5.000988, 4.989071, 4.973829, 
    4.955482, 4.934607, 4.912163, 4.889425, 4.867839, 4.848833, 4.833615, 
    4.823024, 4.817452, 4.816856, 4.820828, 4.828676, 4.839528, 4.852401, 
    4.86627,
  // momentumY(19,35, 0-49)
    4.872328, 4.878919, 4.886526, 4.89474, 4.903203, 4.911632, 4.919809, 
    4.927599, 4.934926, 4.941772, 4.948174, 4.954204, 4.959976, 4.965626, 
    4.971318, 4.976828, 4.978239, 4.982703, 4.986978, 4.990948, 4.99466, 
    4.998809, 5.002337, 5.005319, 5.008259, 5.010948, 5.01328, 5.014896, 
    5.015461, 5.013795, 5.009148, 5.002493, 4.992821, 4.979948, 4.963921, 
    4.945088, 4.92415, 4.90215, 4.880391, 4.860284, 4.843158, 4.83008, 
    4.821725, 4.818338, 4.819746, 4.825438, 4.834654, 4.84647, 4.859871, 
    4.873812,
  // momentumY(19,36, 0-49)
    4.878319, 4.884347, 4.891294, 4.898786, 4.906506, 4.914204, 4.921698, 
    4.928871, 4.935667, 4.942079, 4.948146, 4.953941, 4.95958, 4.965217, 
    4.97104, 4.974863, 4.977667, 4.982239, 4.986354, 4.99006, 4.993469, 
    4.997919, 5.001616, 5.004714, 5.007523, 5.009817, 5.011443, 5.012049, 
    5.011275, 5.008129, 5.00182, 4.994109, 4.98338, 4.969563, 4.952835, 
    4.933675, 4.912894, 4.891598, 4.871095, 4.852732, 4.837718, 4.826962, 
    4.820982, 4.819872, 4.823338, 4.830776, 4.841359, 4.854115, 4.868001, 
    4.881951,
  // momentumY(19,37, 0-49)
    4.884991, 4.890361, 4.896557, 4.903244, 4.910141, 4.917033, 4.923767, 
    4.930253, 4.936448, 4.942355, 4.948011, 4.953487, 4.958893, 4.964376, 
    4.97013, 4.972736, 4.976905, 4.981477, 4.985387, 4.988821, 4.991942, 
    4.996607, 5.000417, 5.003583, 5.006192, 5.008002, 5.008813, 5.008285, 
    5.006043, 5.001339, 4.993384, 4.98456, 4.972786, 4.958107, 4.940834, 
    4.921567, 4.901206, 4.880898, 4.861922, 4.845537, 4.832814, 4.824502, 
    4.820959, 4.822139, 4.827637, 4.836768, 4.848647, 4.862257, 4.876529, 
    4.890384,
  // momentumY(19,38, 0-49)
    4.892121, 4.896754, 4.902132, 4.907953, 4.913973, 4.920011, 4.92594, 
    4.931687, 4.937231, 4.942576, 4.947761, 4.952847, 4.957928, 4.963131, 
    4.968633, 4.970451, 4.975925, 4.980362, 4.984005, 4.987148, 4.989974, 
    4.994747, 4.99859, 5.001753, 5.004083, 5.005324, 5.005226, 5.003472, 
    4.999688, 4.993407, 4.983876, 4.973956, 4.96122, 4.945838, 4.928244, 
    4.909145, 4.889503, 4.870472, 4.853275, 4.839058, 4.828744, 4.82292, 
    4.821793, 4.825191, 4.832617, 4.843311, 4.856339, 4.870652, 4.885157, 
    4.898771,
  // momentumY(19,39, 0-49)
    4.899467, 4.903297, 4.907806, 4.912726, 4.917843, 4.923001, 4.928099, 
    4.933086, 4.937946, 4.942693, 4.947358, 4.951997, 4.95668, 4.961504, 
    4.966603, 4.967971, 4.974646, 4.978811, 4.982118, 4.984936, 4.987445, 
    4.992202, 4.995981, 4.999056, 5.00102, 5.001617, 5.000542, 4.997513, 
    4.99217, 4.984358, 4.973391, 4.962465, 4.948932, 4.93308, 4.915452, 
    4.896836, 4.878227, 4.860754, 4.845551, 4.833638, 4.825777, 4.822405, 
    4.823591, 4.829056, 4.838219, 4.850267, 4.864228, 4.879025, 4.893557, 
    4.906746,
  // momentumY(19,40, 0-49)
    4.906766, 4.909746, 4.913357, 4.917359, 4.921566, 4.925843, 4.930111, 
    4.934331, 4.938495, 4.942622, 4.94674, 4.950891, 4.95512, 4.959492, 
    4.964085, 4.965239, 4.97296, 4.976724, 4.979627, 4.98208, 4.984232, 
    4.988842, 4.992447, 4.995337, 4.996855, 4.996744, 4.994654, 4.990354, 
    4.983506, 4.974283, 4.962084, 4.950325, 4.936236, 4.920212, 4.902885, 
    4.885092, 4.867829, 4.852161, 4.839121, 4.829577, 4.824143, 4.823107, 
    4.82642, 4.833713, 4.844347, 4.857467, 4.872072, 4.887079, 4.901387, 
    4.913939,
  // momentumY(19,41, 0-49)
    4.913755, 4.915848, 4.918544, 4.921631, 4.924941, 4.928359, 4.931815, 
    4.935283, 4.938761, 4.942267, 4.945827, 4.949466, 4.953209, 4.957081, 
    4.961106, 4.962186, 4.970744, 4.974006, 4.976444, 4.97848, 4.980226, 
    4.984553, 4.987868, 4.990473, 4.991469, 4.990608, 4.987513, 4.982002, 
    4.973772, 4.963334, 4.950175, 4.93783, 4.923496, 4.90765, 4.890987, 
    4.874359, 4.858728, 4.845076, 4.8343, 4.827125, 4.824011, 4.825119, 
    4.830297, 4.839108, 4.850871, 4.864708, 4.879611, 4.894502, 4.908296, 
    4.919983,
  // momentumY(19,42, 0-49)
    4.92017, 4.921348, 4.923127, 4.925314, 4.927758, 4.930353, 4.933038, 
    4.935792, 4.938614, 4.94152, 4.944527, 4.94765, 4.950894, 4.954247, 
    4.957675, 4.958741, 4.967895, 4.970575, 4.972492, 4.974058, 4.975332, 
    4.979243, 4.982157, 4.984379, 4.984793, 4.983174, 4.979122, 4.97252, 
    4.963109, 4.951718, 4.937935, 4.92532, 4.911098, 4.895811, 4.880182, 
    4.865045, 4.851295, 4.839802, 4.83133, 4.826448, 4.825478, 4.828466, 
    4.835182, 4.845138, 4.857627, 4.871772, 4.886574, 4.900981, 4.913953, 
    4.924549,
  // momentumY(19,43, 0-49)
    4.925763, 4.926003, 4.926868, 4.928182, 4.929801, 4.931626, 4.933599, 
    4.935696, 4.937914, 4.94026, 4.942748, 4.945375, 4.948125, 4.950956, 
    4.953793, 4.954841, 4.96433, 4.966375, 4.967723, 4.968758, 4.969495, 
    4.972867, 4.975272, 4.977025, 4.97682, 4.974465, 4.969556, 4.962043, 
    4.951717, 4.939699, 4.925668, 4.913147, 4.899427, 4.885087, 4.87084, 
    4.857475, 4.845798, 4.836551, 4.830351, 4.827622, 4.828561, 4.833115, 
    4.840987, 4.851663, 4.86443, 4.878427, 4.892694, 4.906231, 4.91807, 
    4.927366,
  // momentumY(19,44, 0-49)
    4.930317, 4.929597, 4.929554, 4.930022, 4.930867, 4.931989, 4.933323, 
    4.934839, 4.936524, 4.938376, 4.940395, 4.942565, 4.944849, 4.94718, 
    4.949445, 4.950438, 4.960001, 4.961379, 4.962115, 4.96256, 4.962694, 
    4.965418, 4.967226, 4.968439, 4.967605, 4.964572, 4.95895, 4.950758, 
    4.93984, 4.927562, 4.913687, 4.901648, 4.888824, 4.875793, 4.863242, 
    4.85188, 4.842403, 4.835417, 4.831395, 4.830625, 4.833188, 4.838951, 
    4.847569, 4.85851, 4.87108, 4.884458, 4.897746, 4.910027, 4.920442, 
    4.928277,
  // momentumY(19,45, 0-49)
    4.933671, 4.931966, 4.931014, 4.930665, 4.930786, 4.931273, 4.932052, 
    4.933077, 4.934319, 4.935762, 4.937385, 4.939156, 4.941019, 4.942884, 
    4.944615, 4.945492, 4.954885, 4.955587, 4.955676, 4.955476, 4.954947, 
    4.956939, 4.958081, 4.958708, 4.957262, 4.953647, 4.947495, 4.938894, 
    4.92774, 4.915594, 4.902283, 4.89111, 4.879552, 4.868159, 4.857555, 
    4.848358, 4.841139, 4.836369, 4.834379, 4.835332, 4.839209, 4.845804, 
    4.854742, 4.86549, 4.877389, 4.889682, 4.901563, 4.912237, 4.920988, 
    4.927265,
  // momentumY(19,46, 0-49)
    4.935753, 4.933025, 4.931156, 4.930007, 4.929449, 4.929368, 4.929675, 
    4.930304, 4.931202, 4.932328, 4.933641, 4.935088, 4.936592, 4.938042, 
    4.939281, 4.939974, 4.948993, 4.949016, 4.948432, 4.947545, 4.946309, 
    4.947513, 4.947949, 4.947968, 4.945961, 4.941886, 4.935413, 4.926697, 
    4.915676, 4.904049, 4.89169, 4.881741, 4.871771, 4.862283, 4.853815, 
    4.846878, 4.841915, 4.83926, 4.839114, 4.841527, 4.846392, 4.853445, 
    4.862292, 4.872415, 4.883203, 4.893989, 4.904093, 4.912873, 4.919795, 
    4.924508,
  // momentumY(19,47, 0-49)
    4.936611, 4.932811, 4.929999, 4.92805, 4.926839, 4.926242, 4.92615, 
    4.92647, 4.927119, 4.928027, 4.929121, 4.930323, 4.931534, 4.932622, 
    4.93342, 4.933862, 4.942347, 4.941703, 4.94043, 4.938825, 4.936858, 
    4.937251, 4.936972, 4.936396, 4.933905, 4.929514, 4.922946, 4.914406, 
    4.903878, 4.893131, 4.882066, 4.873648, 4.86553, 4.858142, 4.851929, 
    4.847281, 4.844512, 4.843832, 4.84532, 4.848924, 4.854459, 4.861622, 
    4.870004, 4.879118, 4.888425, 4.897368, 4.905418, 4.912122, 4.917159, 
    4.920394,
  // momentumY(19,48, 0-49)
    4.936437, 4.931505, 4.927708, 4.924939, 4.923077, 4.921989, 4.921544, 
    4.921619, 4.922096, 4.922868, 4.923826, 4.924857, 4.925838, 4.926618, 
    4.92702, 4.927145, 4.934983, 4.93369, 4.931725, 4.929393, 4.926692, 
    4.926288, 4.925319, 4.924188, 4.921313, 4.916768, 4.910326, 4.90224, 
    4.892526, 4.88297, 4.87348, 4.866836, 4.860761, 4.855598, 4.851686, 
    4.849298, 4.848623, 4.849751, 4.852652, 4.857186, 4.863106, 4.870075, 
    4.877688, 4.885501, 4.89306, 4.89994, 4.905788, 4.910366, 4.913583, 
    4.915535,
  // momentumY(19,49, 0-49)
    4.939479, 4.932686, 4.927199, 4.922946, 4.919828, 4.917706, 4.916431, 
    4.915837, 4.915757, 4.916022, 4.916465, 4.916909, 4.91717, 4.917032, 
    4.916247, 4.915366, 4.929752, 4.926197, 4.921779, 4.917198, 4.912539, 
    4.913105, 4.913378, 4.914213, 4.912521, 4.90855, 4.901885, 4.89297, 
    4.881677, 4.871408, 4.861761, 4.857852, 4.85482, 4.852896, 4.852281, 
    4.853092, 4.855345, 4.858965, 4.86378, 4.869527, 4.875886, 4.882484, 
    4.888945, 4.894903, 4.900057, 4.904189, 4.907223, 4.909227, 4.910436, 
    4.91124,
  // momentumY(20,0, 0-49)
    4.860252, 4.86001, 4.861908, 4.865577, 4.870636, 4.876714, 4.883478, 
    4.890644, 4.897981, 4.905314, 4.912512, 4.919477, 4.926129, 4.932405, 
    4.938227, 4.943402, 4.949084, 4.953224, 4.956752, 4.959602, 4.961658, 
    4.963098, 4.963417, 4.962541, 4.960215, 4.956271, 4.950531, 4.9429, 
    4.933327, 4.921966, 4.908915, 4.894793, 4.879703, 4.864185, 4.848875, 
    4.834458, 4.821619, 4.810974, 4.803027, 4.798102, 4.796328, 4.797613, 
    4.801653, 4.80796, 4.815895, 4.82473, 4.833702, 4.842091, 4.849298, 
    4.854918,
  // momentumY(20,1, 0-49)
    4.862436, 4.862621, 4.86489, 4.86887, 4.874181, 4.880456, 4.887374, 
    4.894657, 4.902087, 4.909499, 4.91677, 4.923805, 4.93053, 4.936876, 
    4.94276, 4.947818, 4.954359, 4.958505, 4.962062, 4.965001, 4.967188, 
    4.969077, 4.969801, 4.969337, 4.967341, 4.963618, 4.957946, 4.950209, 
    4.94033, 4.92852, 4.914805, 4.900119, 4.884272, 4.867824, 4.851451, 
    4.835898, 4.821912, 4.810189, 4.8013, 4.795636, 4.793375, 4.794456, 
    4.798588, 4.805271, 4.813842, 4.823527, 4.833501, 4.842969, 4.851245, 
    4.857827,
  // momentumY(20,2, 0-49)
    4.864428, 4.86499, 4.867573, 4.871808, 4.877315, 4.883739, 4.890766, 
    4.898131, 4.905627, 4.913094, 4.920412, 4.927494, 4.934264, 4.94065, 
    4.946568, 4.951439, 4.958696, 4.962821, 4.966372, 4.969354, 4.971641, 
    4.973957, 4.97509, 4.97507, 4.97349, 4.970134, 4.964743, 4.957186, 
    4.947346, 4.935463, 4.921481, 4.90663, 4.890397, 4.873343, 4.856158, 
    4.839617, 4.824526, 4.811648, 4.801634, 4.794953, 4.791851, 4.792322, 
    4.79611, 4.802735, 4.811536, 4.821715, 4.832422, 4.842813, 4.852137, 
    4.85981,
  // momentumY(20,3, 0-49)
    4.866155, 4.86705, 4.869899, 4.874338, 4.879996, 4.886528, 4.893631, 
    4.90105, 4.908585, 4.916081, 4.923425, 4.930527, 4.937315, 4.943715, 
    4.949641, 4.954255, 4.962042, 4.966132, 4.969641, 4.972626, 4.974976, 
    4.977679, 4.979204, 4.979639, 4.978534, 4.975669, 4.970754, 4.963642, 
    4.954173, 4.94259, 4.928738, 4.914125, 4.897903, 4.880599, 4.862891, 
    4.845562, 4.829454, 4.815392, 4.804106, 4.796156, 4.791875, 4.791333, 
    4.794338, 4.800455, 4.809047, 4.819333, 4.830458, 4.841559, 4.851843, 
    4.860661,
  // momentumY(20,4, 0-49)
    4.867635, 4.868824, 4.871896, 4.876496, 4.882263, 4.888866, 4.896011, 
    4.903454, 4.910999, 4.918499, 4.925837, 4.932927, 4.939702, 4.946087, 
    4.952006, 4.956291, 4.964385, 4.968431, 4.971873, 4.974825, 4.977198, 
    4.980241, 4.982126, 4.982999, 4.982406, 4.980123, 4.975844, 4.969408, 
    4.960617, 4.949678, 4.936331, 4.922343, 4.906526, 4.889344, 4.871434, 
    4.85356, 4.836578, 4.82136, 4.808711, 4.799289, 4.793529, 4.791602, 
    4.793405, 4.798576, 4.80653, 4.816529, 4.827738, 4.8393, 4.850401, 
    4.860345,
  // momentumY(20,5, 0-49)
    4.868941, 4.870391, 4.873652, 4.878376, 4.884216, 4.890854, 4.898007, 
    4.905436, 4.912956, 4.920418, 4.927711, 4.934752, 4.941473, 4.947814, 
    4.953711, 4.957606, 4.965757, 4.969759, 4.973117, 4.976005, 4.978372, 
    4.981693, 4.983891, 4.98517, 4.985097, 4.983453, 4.979932, 4.97436, 
    4.966503, 4.956503, 4.944001, 4.930983, 4.915935, 4.899241, 4.881466, 
    4.863327, 4.845665, 4.82938, 4.815343, 4.80431, 4.796834, 4.793207, 
    4.793438, 4.797264, 4.804183, 4.813521, 4.824488, 4.836249, 4.84799, 
    4.858978,
  // momentumY(20,6, 0-49)
    4.870184, 4.871867, 4.875287, 4.880104, 4.885983, 4.892617, 4.899735, 
    4.907109, 4.914557, 4.921935, 4.929136, 4.936078, 4.942703, 4.948964, 
    4.95482, 4.958287, 4.966236, 4.970192, 4.97346, 4.976264, 4.978598, 
    4.982133, 4.984593, 4.986225, 4.986656, 4.985677, 4.982993, 4.978419, 
    4.971696, 4.962874, 4.95149, 4.939726, 4.925767, 4.9099, 4.892593, 
    4.874488, 4.856383, 4.83918, 4.823804, 4.8111, 4.801749, 4.796178, 
    4.794536, 4.796683, 4.802223, 4.810569, 4.820991, 4.832695, 4.844877, 
    4.856782,
  // momentumY(20,7, 0-49)
    4.871486, 4.873385, 4.876938, 4.881816, 4.887699, 4.894289, 4.901329, 
    4.908598, 4.915922, 4.923161, 4.930209, 4.936997, 4.943477, 4.949618, 
    4.955414, 4.958443, 4.965936, 4.969844, 4.97302, 4.975732, 4.978019, 
    4.981705, 4.984363, 4.986288, 4.987187, 4.986865, 4.985055, 4.981565, 
    4.976113, 4.968638, 4.958585, 4.948279, 4.935663, 4.92091, 4.904378, 
    4.886606, 4.868324, 4.850407, 4.833809, 4.819458, 4.808159, 4.800493, 
    4.796761, 4.796972, 4.800858, 4.807934, 4.81755, 4.828959, 4.841378, 
    4.854039,
  // momentumY(20,8, 0-49)
    4.872965, 4.875064, 4.878729, 4.883643, 4.889493, 4.895999, 4.902913, 
    4.910024, 4.917163, 4.924199, 4.931038, 4.937615, 4.943896, 4.949877, 
    4.955583, 4.958203, 4.965009, 4.968857, 4.971947, 4.974571, 4.976808, 
    4.980578, 4.983373, 4.98552, 4.986834, 4.987137, 4.986202, 4.983829, 
    4.979728, 4.973704, 4.965117, 4.956395, 4.945295, 4.931881, 4.916384, 
    4.899226, 4.88104, 4.862648, 4.845007, 4.829113, 4.815887, 4.806065, 
    4.800118, 4.798223, 4.800258, 4.805854, 4.81445, 4.825356, 4.837813, 
    4.851048,
  // momentumY(20,9, 0-49)
    4.874715, 4.877008, 4.88077, 4.885693, 4.891478, 4.897859, 4.904594, 
    4.911492, 4.918387, 4.925161, 4.931726, 4.938032, 4.944063, 4.949836, 
    4.955409, 4.957707, 4.963628, 4.967393, 4.970406, 4.972955, 4.975152, 
    4.978941, 4.981811, 4.984108, 4.985774, 4.98665, 4.986557, 4.985291, 
    4.982565, 4.978032, 4.970989, 4.96389, 4.954402, 4.942473, 4.928211, 
    4.911908, 4.894079, 4.87547, 4.857014, 4.839749, 4.824699, 4.812755, 
    4.804565, 4.800483, 4.800548, 4.804519, 4.811933, 4.82216, 4.834473, 
    4.848091,
  // momentumY(20,10, 0-49)
    4.876799, 4.879285, 4.883133, 4.888045, 4.893735, 4.899947, 4.906461, 
    4.913087, 4.919682, 4.926131, 4.932365, 4.938345, 4.944074, 4.949587, 
    4.954967, 4.957089, 4.961978, 4.965627, 4.968569, 4.971067, 4.973243, 
    4.97699, 4.979874, 4.98225, 4.984199, 4.985584, 4.986276, 4.986076, 
    4.984701, 4.981645, 4.976162, 4.970654, 4.962789, 4.952418, 4.939521, 
    4.924259, 4.907021, 4.88845, 4.869433, 4.851023, 4.834328, 4.82038, 
    4.810005, 4.803736, 4.801787, 4.804056, 4.810177, 4.819589, 4.831591, 
    4.845403,
  // momentumY(20,11, 0-49)
    4.879239, 4.881923, 4.885851, 4.890735, 4.896304, 4.902315, 4.908561, 
    4.91487, 4.921111, 4.927186, 4.933039, 4.938643, 4.944018, 4.949213, 
    4.954324, 4.956469, 4.960239, 4.963728, 4.966609, 4.969083, 4.971266, 
    4.974913, 4.977757, 4.980145, 4.982306, 4.984129, 4.985535, 4.986328, 
    4.986242, 4.98461, 4.980663, 4.976647, 4.97035, 4.961532, 4.950062, 
    4.935967, 4.919504, 4.901208, 4.881889, 4.862591, 4.844482, 4.828718, 
    4.816289, 4.807916, 4.80398, 4.804524, 4.80929, 4.81778, 4.829328, 
    4.843155,
  // momentumY(20,12, 0-49)
    4.88201, 4.884904, 4.888915, 4.893763, 4.899191, 4.904974, 4.910917, 
    4.916871, 4.922716, 4.928374, 4.933802, 4.938989, 4.943964, 4.948782, 
    4.953533, 4.95595, 4.958569, 4.961857, 4.964685, 4.967168, 4.969397, 
    4.972889, 4.975645, 4.977991, 4.980297, 4.982482, 4.984518, 4.986214, 
    4.987322, 4.987028, 4.984559, 4.981891, 4.977048, 4.969718, 4.959666, 
    4.946801, 4.93125, 4.913426, 4.894051, 4.874133, 4.854875, 4.837531, 
    4.823242, 4.812902, 4.807063, 4.805912, 4.809299, 4.816798, 4.827771, 
    4.841449,
  // momentumY(20,13, 0-49)
    4.885045, 4.888165, 4.892267, 4.897079, 4.902358, 4.907895, 4.913514, 
    4.919086, 4.924509, 4.929721, 4.934696, 4.939434, 4.943967, 4.948348, 
    4.952642, 4.955595, 4.957088, 4.960145, 4.962937, 4.965468, 4.967791, 
    4.971079, 4.973709, 4.975964, 4.978357, 4.980833, 4.98341, 4.985902, 
    4.98809, 4.989025, 4.987952, 4.986454, 4.982911, 4.976952, 4.968254, 
    4.956622, 4.942061, 4.92486, 4.905646, 4.885368, 4.865235, 4.846574, 
    4.830656, 4.818532, 4.810918, 4.808143, 4.810166, 4.816629, 4.826932, 
    4.840311,
  // momentumY(20,14, 0-49)
    4.888229, 4.8916, 4.895807, 4.900593, 4.905726, 4.911015, 4.916304, 
    4.921482, 4.92647, 4.931225, 4.935732, 4.940003, 4.944067, 4.947958, 
    4.951711, 4.955437, 4.955875, 4.958696, 4.961479, 4.964108, 4.966577, 
    4.969624, 4.9721, 4.974234, 4.976667, 4.979364, 4.98239, 4.985562, 
    4.988698, 4.990733, 4.990968, 4.99044, 4.988013, 4.983267, 4.975816, 
    4.965367, 4.951819, 4.935346, 4.916467, 4.896061, 4.875321, 4.855616, 
    4.838318, 4.824619, 4.815388, 4.811089, 4.811786, 4.817195, 4.826753, 
    4.839705,
  // momentumY(20,15, 0-49)
    4.891417, 4.895063, 4.899403, 4.904181, 4.909182, 4.914233, 4.919199, 
    4.923991, 4.928551, 4.932856, 4.936903, 4.940707, 4.944289, 4.947664, 
    4.950818, 4.955467, 4.954948, 4.957564, 4.96039, 4.963179, 4.965862, 
    4.968639, 4.970955, 4.972952, 4.975391, 4.978249, 4.981628, 4.985358, 
    4.989294, 4.99229, 4.993727, 4.993963, 4.99245, 4.988739, 4.982389, 
    4.973036, 4.96048, 4.944787, 4.926372, 4.906035, 4.884928, 4.864438, 
    4.846014, 4.830963, 4.820285, 4.814578, 4.81401, 4.818363, 4.827119, 
    4.839538,
  // momentumY(20,16, 0-49)
    4.894438, 4.898385, 4.902883, 4.90768, 4.912577, 4.917415, 4.922084, 
    4.926518, 4.93068, 4.934565, 4.938181, 4.941544, 4.944665, 4.94753, 
    4.950081, 4.955651, 4.954271, 4.956758, 4.959707, 4.962741, 4.965721, 
    4.968219, 4.970386, 4.972255, 4.974681, 4.977648, 4.981289, 4.985443, 
    4.990022, 4.993821, 4.99635, 4.997137, 4.996331, 4.993463, 4.98805, 
    4.97967, 4.968042, 4.953138, 4.935272, 4.915156, 4.893888, 4.87285, 
    4.853538, 4.837351, 4.825407, 4.818417, 4.816652, 4.819967, 4.827884, 
    4.839682,
  // momentumY(20,17, 0-49)
    4.897111, 4.901378, 4.906057, 4.910903, 4.915725, 4.920388, 4.924805, 
    4.92893, 4.93275, 4.936276, 4.939528, 4.942516, 4.945239, 4.947652, 
    4.949658, 4.955938, 4.95375, 4.956237, 4.959424, 4.962814, 4.966193, 
    4.968428, 4.970485, 4.972262, 4.974679, 4.977714, 4.981524, 4.985966, 
    4.991012, 4.995444, 4.99893, 5.000061, 4.999754, 4.997528, 4.992876, 
    4.985324, 4.974533, 4.960389, 4.943113, 4.92333, 4.90207, 4.880688, 
    4.860705, 4.843585, 4.830546, 4.822402, 4.819518, 4.82182, 4.828876, 
    4.839989,
  // momentumY(20,18, 0-49)
    4.899259, 4.903844, 4.908713, 4.913628, 4.918412, 4.922945, 4.927167, 
    4.931057, 4.934627, 4.9379, 4.940901, 4.943637, 4.946083, 4.948168, 
    4.94976, 4.956294, 4.953275, 4.955921, 4.959491, 4.963376, 4.967283, 
    4.969299, 4.971318, 4.973071, 4.97551, 4.97859, 4.98248, 4.987064, 
    4.992386, 4.997256, 5.001545, 5.002809, 5.002788, 5.001004, 4.996927, 
    4.990052, 4.979986, 4.966546, 4.949867, 4.930487, 4.909364, 4.887812, 
    4.867347, 4.849483, 4.83551, 4.826337, 4.822413, 4.823737, 4.829926, 
    4.840314,
  // momentumY(20,19, 0-49)
    4.900722, 4.905582, 4.910621, 4.915603, 4.920366, 4.924819, 4.928921, 
    4.932685, 4.936142, 4.939328, 4.942264, 4.944942, 4.947306, 4.949254, 
    4.950626, 4.956723, 4.952731, 4.955709, 4.959822, 4.964365, 4.968961, 
    4.970843, 4.972939, 4.974776, 4.977301, 4.980426, 4.984317, 4.988889, 
    4.994273, 4.99935, 5.004237, 5.005415, 5.005468, 5.00392, 5.000231, 
    4.993872, 4.984408, 4.971598, 4.9555, 4.936566, 4.915679, 4.894096, 
    4.873318, 4.854876, 4.840123, 4.83004, 4.825162, 4.825555, 4.830888, 
    4.840529,
  // momentumY(20,20, 0-49)
    4.90239, 4.908547, 4.914843, 4.921025, 4.926898, 4.932327, 4.937214, 
    4.9415, 4.945158, 4.948183, 4.950596, 4.952441, 4.953793, 4.954744, 
    4.955407, 0, 4.958249, 4.960236, 4.962961, 4.965996, 4.969181, 4.968955, 
    4.969491, 4.97025, 4.972277, 4.975456, 4.979868, 4.985317, 4.991841, 
    4.998215, 5.004694, 5.006587, 5.007314, 5.006402, 5.00332, 4.997553, 
    4.988664, 4.976397, 4.960779, 4.942212, 4.921516, 4.899904, 4.878851, 
    4.859899, 4.844436, 4.83351, 4.827723, 4.827208, 4.831687, 4.840559,
  // momentumY(20,21, 0-49)
    4.902546, 4.909152, 4.915813, 4.922264, 4.928308, 4.93382, 4.938725, 
    4.942987, 4.946609, 4.949608, 4.952027, 4.953918, 4.955361, 4.956449, 
    4.957307, 0, 4.95625, 4.958742, 4.96202, 4.965616, 4.96931, 4.968532, 
    4.968688, 4.969118, 4.970976, 4.974154, 4.978734, 4.984498, 4.991485, 
    4.998459, 5.005868, 5.007966, 5.009057, 5.008655, 5.006201, 5.001147, 
    4.99302, 4.981514, 4.966591, 4.948582, 4.928237, 4.906707, 4.885434, 
    4.865964, 4.849724, 4.837832, 4.830966, 4.829334, 4.832719, 4.840568,
  // momentumY(20,22, 0-49)
    4.902033, 4.909122, 4.916215, 4.92303, 4.929366, 4.935092, 4.940144, 
    4.944501, 4.948182, 4.951223, 4.953678, 4.955619, 4.957127, 4.958311, 
    4.959311, 0, 4.955119, 4.958027, 4.96179, 4.965904, 4.970087, 4.968813, 
    4.968649, 4.968804, 4.970531, 4.973706, 4.978404, 4.984384, 4.991682, 
    4.999045, 5.007104, 5.009167, 5.010358, 5.010189, 5.00809, 5.003501, 
    4.995925, 4.985018, 4.970692, 4.953214, 4.933263, 4.911923, 4.89059, 
    4.870792, 4.853981, 4.841319, 4.833551, 4.830953, 4.833365, 4.84028,
  // momentumY(20,23, 0-49)
    4.900946, 4.908532, 4.916096, 4.92334, 4.930048, 4.936085, 4.941385, 
    4.945931, 4.949752, 4.952897, 4.955433, 4.95744, 4.959013, 4.96027, 
    4.961375, 0, 4.954969, 4.958154, 4.962238, 4.966699, 4.971208, 4.969459, 
    4.96897, 4.968847, 4.970413, 4.973536, 4.978281, 4.984387, 4.991886, 
    4.999502, 5.008006, 5.009949, 5.011131, 5.011066, 5.009185, 5.00492, 
    4.99776, 4.987338, 4.973525, 4.956533, 4.936977, 4.915878, 4.894584, 
    4.874597, 4.857371, 4.844103, 4.835588, 4.832156, 4.833704, 4.839765,
  // momentumY(20,24, 0-49)
    4.899428, 4.907504, 4.915555, 4.92326, 4.930388, 4.936795, 4.942407, 
    4.947209, 4.951232, 4.95453, 4.957183, 4.959279, 4.96092, 4.962241, 
    4.963425, 0, 4.95597, 4.959291, 4.963529, 4.968157, 4.972827, 4.970741, 
    4.970021, 4.969701, 4.971145, 4.974215, 4.978966, 4.985128, 4.992729, 
    5.000482, 5.009243, 5.011076, 5.012208, 5.012159, 5.010361, 5.006243, 
    4.999289, 4.98912, 4.975582, 4.958858, 4.939522, 4.918553, 4.897259, 
    4.877122, 4.859592, 4.845881, 4.836812, 4.832757, 4.833642, 4.839036,
  // momentumY(20,25, 0-49)
    4.897653, 4.906196, 4.91472, 4.922887, 4.93045, 4.937253, 4.943209, 
    4.948304, 4.952564, 4.956049, 4.958841, 4.961037, 4.962751, 4.964127, 
    4.965363, 0, 4.957728, 4.961046, 4.96527, 4.969884, 4.974544, 4.972311, 
    4.971497, 4.971106, 4.972506, 4.975554, 4.980302, 4.986476, 4.994102, 
    5.001885, 5.010712, 5.012488, 5.013579, 5.013506, 5.011698, 5.007585, 
    5.000655, 4.990522, 4.977032, 4.960351, 4.941041, 4.920062, 4.898702, 
    4.878432, 4.860693, 4.846697, 4.837277, 4.832819, 4.833266, 4.838201,
  // momentumY(20,26, 0-49)
    4.895818, 4.904783, 4.913742, 4.922344, 4.930325, 4.937515, 4.943821, 
    4.949216, 4.953726, 4.957407, 4.960343, 4.962636, 4.964409, 4.965817, 
    4.967063, 0, 4.960133, 4.963308, 4.967357, 4.971776, 4.976251, 4.974082, 
    4.973327, 4.973009, 4.974462, 4.977538, 4.982289, 4.98844, 4.996022, 
    5.003737, 5.012439, 5.014235, 5.015309, 5.015183, 5.013282, 5.009041, 
    5.001948, 4.99163, 4.97794, 4.961062, 4.941566, 4.920424, 4.898925, 
    4.878536, 4.860688, 4.846581, 4.837034, 4.832421, 4.832682, 4.8374,
  // momentumY(20,27, 0-49)
    4.894114, 4.903435, 4.912771, 4.921757, 4.930116, 4.937665, 4.944301, 
    4.949985, 4.954732, 4.958596, 4.961658, 4.964022, 4.965817, 4.967206, 
    4.968397, 0, 4.96324, 4.966122, 4.969824, 4.973864, 4.97798, 4.976048, 
    4.975473, 4.975338, 4.976915, 4.98005, 4.984796, 4.990885, 4.998345, 
    5.00589, 5.014274, 5.016143, 5.01721, 5.016988, 5.014902, 5.010391, 
    5.002958, 4.992247, 4.978143, 4.960862, 4.941015, 4.919603, 4.897938, 
    4.87749, 4.859674, 4.845661, 4.836235, 4.831735, 4.832074, 4.836821,
  // momentumY(20,28, 0-49)
    4.892716, 4.902316, 4.911954, 4.921258, 4.92994, 4.937809, 4.94474, 
    4.950686, 4.955645, 4.959659, 4.962801, 4.965176, 4.966919, 4.9682, 
    4.969231, 0, 4.967395, 4.969824, 4.972999, 4.976473, 4.980055, 4.978459, 
    4.97812, 4.978223, 4.979947, 4.983134, 4.987837, 4.993802, 5.001053, 
    5.008318, 5.016205, 5.018162, 5.019183, 5.018777, 5.016371, 5.011417, 
    5.00344, 4.992121, 4.977393, 4.95953, 4.939205, 4.917471, 4.895676, 
    4.875288, 4.8577, 4.844033, 4.835011, 4.830916, 4.831614, 4.836638,
  // momentumY(20,29, 0-49)
    4.891768, 4.901561, 4.91142, 4.920973, 4.929929, 4.938075, 4.945275, 
    4.951451, 4.956579, 4.960682, 4.963824, 4.966108, 4.967679, 4.968717, 
    4.969442, 0, 4.972353, 4.974166, 4.976633, 4.979355, 4.982222, 4.980926, 
    4.980772, 4.981068, 4.982892, 4.986081, 4.990681, 4.996451, 5.003397, 
    5.010265, 5.017463, 5.019434, 5.020311, 5.019595, 5.016734, 5.011202, 
    5.002559, 4.990538, 4.975133, 4.956691, 4.935954, 4.914032, 4.892297, 
    4.872213, 4.855128, 4.842093, 4.833755, 4.830319, 4.831594, 4.837072,
  // momentumY(20,30, 0-49)
    4.890552, 4.899473, 4.908428, 4.917069, 4.925149, 4.932522, 4.939125, 
    4.94497, 4.950115, 4.954631, 4.958583, 4.961999, 4.964857, 4.967066, 
    4.968472, 4.979602, 4.96907, 4.971892, 4.976008, 4.980648, 4.98542, 
    4.986781, 4.988743, 4.990612, 4.993301, 4.996634, 5.000715, 5.005429, 
    5.010921, 5.01609, 5.021275, 5.022079, 5.021772, 5.019878, 5.015864, 
    5.009229, 4.99956, 4.986626, 4.970476, 4.951515, 4.930534, 4.90868, 
    4.887331, 4.867914, 4.851709, 4.839678, 4.832371, 4.829907, 4.832027, 
    4.838179,
  // momentumY(20,31, 0-49)
    4.890921, 4.899925, 4.908952, 4.91766, 4.925797, 4.93321, 4.939828, 
    4.945653, 4.950732, 4.95514, 4.958956, 4.962236, 4.965003, 4.967213, 
    4.968752, 4.979363, 4.971177, 4.97361, 4.977141, 4.98109, 4.985148, 
    4.986675, 4.988585, 4.990395, 4.993023, 4.996342, 5.00046, 5.005226, 
    5.010689, 5.015679, 5.020274, 5.021196, 5.02085, 5.01876, 5.014407, 
    5.007318, 4.997122, 4.983652, 4.967027, 4.947731, 4.926632, 4.904924, 
    4.883998, 4.865252, 4.849897, 4.83881, 4.832448, 4.830843, 4.833675, 
    4.840341,
  // momentumY(20,32, 0-49)
    4.891858, 4.900726, 4.909607, 4.918174, 4.926184, 4.933486, 4.940012, 
    4.945757, 4.950766, 4.955113, 4.958885, 4.962158, 4.964985, 4.967364, 
    4.969228, 4.978518, 4.972463, 4.974708, 4.977826, 4.98125, 4.984755, 
    4.986572, 4.988569, 4.990442, 4.993085, 4.996394, 5.000472, 5.005139, 
    5.010365, 5.014951, 5.01875, 5.019603, 5.019039, 5.016583, 5.011744, 
    5.004078, 4.993276, 4.979236, 4.962163, 4.942626, 4.921564, 4.900208, 
    4.879947, 4.86213, 4.847888, 4.837993, 4.832799, 4.832254, 4.835965, 
    4.843286,
  // momentumY(20,33, 0-49)
    4.893402, 4.901961, 4.910522, 4.918782, 4.926514, 4.933579, 4.93991, 
    4.945505, 4.950407, 4.954688, 4.958445, 4.961763, 4.964719, 4.96735, 
    4.96964, 4.977197, 4.973083, 4.975312, 4.978167, 4.981205, 4.984287, 
    4.986477, 4.98866, 4.990693, 4.993394, 4.996678, 5.000629, 5.005051, 
    5.009844, 5.013827, 5.016671, 5.017282, 5.016326, 5.013347, 5.00788, 
    4.999536, 4.988063, 4.973445, 4.955978, 4.936319, 4.915467, 4.894683, 
    4.87533, 4.858694, 4.845803, 4.83732, 4.833489, 4.834168, 4.838899, 
    4.846986,
  // momentumY(20,34, 0-49)
    4.89555, 4.903658, 4.911766, 4.919588, 4.926923, 4.933646, 4.939695, 
    4.945072, 4.949821, 4.954011, 4.957741, 4.961105, 4.964197, 4.967091, 
    4.969819, 4.975549, 4.97322, 4.975553, 4.978248, 4.981001, 4.983756, 
    4.986354, 4.988786, 4.991036, 4.993814, 4.997042, 5.000778, 5.004812, 
    5.008993, 5.012204, 5.01397, 5.014173, 5.01267, 5.009023, 5.002813, 
    4.993709, 4.981535, 4.966369, 4.9486, 4.928967, 4.908524, 4.88854, 
    4.870338, 4.855117, 4.843793, 4.836905, 4.834589, 4.836618, 4.842463, 
    4.851387,
  // momentumY(20,35, 0-49)
    4.898267, 4.905814, 4.913355, 4.920641, 4.92749, 4.933788, 4.939488, 
    4.944591, 4.949139, 4.953203, 4.956876, 4.960257, 4.963455, 4.966567, 
    4.969674, 4.973719, 4.973058, 4.975548, 4.978137, 4.98067, 4.983167, 
    4.986171, 4.988875, 4.991373, 4.994223, 4.997348, 5.000774, 5.004288, 
    5.007689, 5.009979, 5.010575, 5.010211, 5.008013, 5.003575, 4.996533, 
    4.986623, 4.973759, 4.958113, 4.940172, 4.920749, 4.900939, 4.881996, 
    4.865181, 4.851587, 4.842009, 4.83686, 4.836168, 4.83962, 4.846628, 
    4.856417,
  // momentumY(20,36, 0-49)
    4.901495, 4.908389, 4.915284, 4.921958, 4.92825, 4.934066, 4.939364, 
    4.944149, 4.948456, 4.952359, 4.955939, 4.959299, 4.962548, 4.965801, 
    4.969179, 4.971826, 4.972733, 4.975375, 4.977877, 4.980225, 4.982509, 
    4.985884, 4.988856, 4.991599, 4.994495, 4.99746, 5.00048, 5.003342, 
    5.005812, 5.007051, 5.006406, 5.005326, 5.002304, 4.996975, 4.989042, 
    4.97832, 4.964816, 4.948807, 4.930867, 4.911874, 4.892938, 4.87528, 
    4.860076, 4.848299, 4.84061, 4.837299, 4.838289, 4.843188, 4.85136, 
    4.861993,
  // momentumY(20,37, 0-49)
    4.905167, 4.911334, 4.917521, 4.923526, 4.929215, 4.934506, 4.939363, 
    4.943795, 4.947833, 4.95154, 4.954994, 4.958288, 4.961529, 4.964836, 
    4.968349, 4.969948, 4.972336, 4.975077, 4.977478, 4.979656, 4.981754, 
    4.985441, 4.988646, 4.991607, 4.994504, 4.99724, 4.999755, 5.001844, 
    5.003247, 5.003323, 5.001387, 4.999458, 4.995503, 4.989217, 4.980371, 
    4.968874, 4.954834, 4.938624, 4.9209, 4.902584, 4.884777, 4.868644, 
    4.855253, 4.845448, 4.839749, 4.838326, 4.841006, 4.847328, 4.856611, 
    4.868018,
  // momentumY(20,38, 0-49)
    4.909193, 4.914583, 4.920015, 4.925317, 4.930371, 4.935106, 4.939497, 
    4.943548, 4.947289, 4.950776, 4.954073, 4.957259, 4.960435, 4.96371, 
    4.967225, 4.968122, 4.971893, 4.974655, 4.976923, 4.97893, 4.980852, 
    4.984771, 4.988155, 4.991285, 4.994119, 4.996551, 4.998464, 4.999669, 
    4.999884, 4.99871, 4.995449, 4.992558, 4.987595, 4.98032, 4.970589, 
    4.958406, 4.943982, 4.927779, 4.910518, 4.893145, 4.876726, 4.862342, 
    4.85094, 4.84322, 4.839568, 4.840035, 4.844362, 4.852028, 4.862319, 
    4.874377,
  // momentumY(20,39, 0-49)
    4.913477, 4.918053, 4.922704, 4.927279, 4.931678, 4.93584, 4.939745, 
    4.943396, 4.946823, 4.950062, 4.953173, 4.956218, 4.959277, 4.962446, 
    4.965847, 4.966341, 4.971383, 4.974071, 4.976166, 4.977993, 4.979737, 
    4.983795, 4.987283, 4.990516, 4.993211, 4.995252, 4.99647, 4.996691, 
    4.995628, 4.99314, 4.988544, 4.984612, 4.978605, 4.970356, 4.959818, 
    4.94709, 4.932482, 4.916533, 4.900011, 4.883851, 4.869068, 4.856631, 
    4.847351, 4.841784, 4.840184, 4.842492, 4.848373, 4.857256, 4.868401, 
    4.880943,
  // momentumY(20,40, 0-49)
    4.917906, 4.921646, 4.925501, 4.929339, 4.933074, 4.936653, 4.940061, 
    4.9433, 4.946392, 4.949367, 4.952266, 4.955137, 4.958039, 4.961041, 
    4.964238, 4.964564, 4.970736, 4.97326, 4.975143, 4.976772, 4.978323, 
    4.982419, 4.985922, 4.989172, 4.991644, 4.993212, 4.993649, 4.99281, 
    4.990404, 4.98657, 4.980658, 4.975645, 4.968606, 4.959457, 4.948241, 
    4.93516, 4.920611, 4.905192, 4.889691, 4.87501, 4.86208, 4.851747, 
    4.844676, 4.84128, 4.841683, 4.845729, 4.853019, 4.862945, 4.874746, 
    4.887564,
  // momentumY(20,41, 0-49)
    4.922345, 4.925241, 4.928298, 4.9314, 4.934471, 4.937466, 4.940372, 
    4.943191, 4.945935, 4.948627, 4.951293, 4.953965, 4.956676, 4.95947, 
    4.9624, 4.962718, 4.969854, 4.972135, 4.973769, 4.975179, 4.976512, 
    4.980538, 4.983962, 4.987133, 4.989291, 4.9903, 4.98989, 4.987938, 
    4.984165, 4.978992, 4.971818, 4.965739, 4.957735, 4.94781, 4.936104, 
    4.92291, 4.908694, 4.894094, 4.879889, 4.866925, 4.856025, 4.847902, 
    4.84307, 4.841802, 4.844105, 4.849738, 4.858246, 4.868992, 4.881212, 
    4.894058,
  // momentumY(20,42, 0-49)
    4.926642, 4.928699, 4.930964, 4.93334, 4.935758, 4.938178, 4.940584, 
    4.942979, 4.945368, 4.947763, 4.950179, 4.95263, 4.955127, 4.957681, 
    4.960309, 4.96071, 4.96862, 4.970598, 4.971952, 4.973114, 4.974197, 
    4.978046, 4.981288, 4.98428, 4.986035, 4.986415, 4.985108, 4.982025, 
    4.976905, 4.970449, 4.962109, 4.955034, 4.946192, 4.935675, 4.923714, 
    4.910677, 4.897085, 4.88359, 4.870934, 4.859879, 4.851132, 4.845262, 
    4.842635, 4.843394, 4.847439, 4.854456, 4.863945, 4.875252, 4.887619, 
    4.900222,
  // momentumY(20,43, 0-49)
    4.930626, 4.931849, 4.933344, 4.935014, 4.936798, 4.938658, 4.940579, 
    4.942554, 4.944587, 4.94668, 4.948834, 4.951047, 4.953313, 4.955612, 
    4.957922, 4.958442, 4.966921, 4.968552, 4.9696, 4.970482, 4.971275, 
    4.974844, 4.977806, 4.980515, 4.981785, 4.981482, 4.979256, 4.975064, 
    4.968668, 4.961029, 4.951668, 4.943729, 4.934234, 4.923361, 4.911418, 
    4.898832, 4.886153, 4.874021, 4.86312, 4.854114, 4.847578, 4.843935, 
    4.843416, 4.846041, 4.851618, 4.85977, 4.869962, 4.881538, 4.893755, 
    4.905829,
  // momentumY(20,44, 0-49)
    4.93411, 4.934515, 4.935261, 4.936253, 4.937433, 4.938762, 4.940217, 
    4.941791, 4.943477, 4.94527, 4.94716, 4.949131, 4.951157, 4.953195, 
    4.955183, 4.955816, 4.964656, 4.965913, 4.966628, 4.967195, 4.967651, 
    4.970848, 4.973435, 4.975765, 4.976482, 4.975461, 4.972332, 4.967094, 
    4.959548, 4.950883, 4.940692, 4.93208, 4.922171, 4.911213, 4.89958, 
    4.887739, 4.876243, 4.865695, 4.856701, 4.849814, 4.845474, 4.843967, 
    4.845396, 4.84967, 4.856519, 4.865516, 4.876104, 4.887634, 4.899394, 
    4.910653,
  // momentumY(20,45, 0-49)
    4.936903, 4.936502, 4.936521, 4.936871, 4.937485, 4.938321, 4.939349, 
    4.940551, 4.941915, 4.943424, 4.945058, 4.946791, 4.948578, 4.950358, 
    4.952039, 4.952745, 4.961742, 4.962612, 4.962971, 4.963184, 4.963254, 
    4.965993, 4.968124, 4.96999, 4.970107, 4.968362, 4.964381, 4.958209, 
    4.949688, 4.940206, 4.929422, 4.920379, 4.910328, 4.899585, 4.888559, 
    4.877738, 4.867655, 4.858856, 4.851855, 4.847086, 4.844861, 4.845332, 
    4.848487, 4.854145, 4.861969, 4.87149, 4.882148, 4.893308, 4.904304, 
    4.914479,
  // momentumY(20,46, 0-49)
    4.938819, 4.937624, 4.936943, 4.936685, 4.936779, 4.93717, 4.937817, 
    4.938693, 4.939772, 4.94103, 4.942434, 4.943947, 4.945509, 4.947042, 
    4.948433, 4.949158, 4.958127, 4.958603, 4.958583, 4.958401, 4.958039, 
    4.960252, 4.961856, 4.963193, 4.962687, 4.960245, 4.955501, 4.948549, 
    4.939279, 4.929226, 4.918125, 4.908927, 4.899035, 4.888804, 4.878668, 
    4.869109, 4.860616, 4.853668, 4.848677, 4.845958, 4.845698, 4.847935, 
    4.852553, 4.859291, 4.86776, 4.877473, 4.887864, 4.898334, 4.908283, 
    4.91715,
  // momentumY(20,47, 0-49)
    4.93972, 4.937729, 4.936366, 4.935534, 4.935153, 4.935151, 4.935477, 
    4.936083, 4.936932, 4.937986, 4.939202, 4.940526, 4.941891, 4.9432, 
    4.944324, 4.945001, 4.953781, 4.953864, 4.95344, 4.952825, 4.951988, 
    4.953621, 4.954652, 4.955418, 4.954295, 4.951216, 4.945836, 4.938297, 
    4.928536, 4.918194, 4.907071, 4.898016, 4.888585, 4.879151, 4.870152, 
    4.862043, 4.85526, 4.850199, 4.847168, 4.84637, 4.847877, 4.851622, 
    4.857403, 4.864896, 4.873673, 4.883236, 4.893039, 4.902533, 4.911198, 
    4.918588,
  // momentumY(20,48, 0-49)
    4.939519, 4.93672, 4.934682, 4.933303, 4.932487, 4.932148, 4.932213, 
    4.932616, 4.933301, 4.934213, 4.935294, 4.936477, 4.937681, 4.938794, 
    4.939677, 4.940239, 4.948703, 4.94839, 4.94754, 4.946457, 4.945107, 
    4.946132, 4.946567, 4.946746, 4.945043, 4.94142, 4.935561, 4.927656, 
    4.917686, 4.907351, 4.896503, 4.88789, 4.879201, 4.870818, 4.863158, 
    4.856635, 4.85162, 4.848419, 4.847244, 4.848188, 4.851223, 4.856192, 
    4.862821, 4.870739, 4.879495, 4.888591, 4.89752, 4.905799, 4.913006, 
    4.918834,
  // momentumY(20,49, 0-49)
    4.940613, 4.936409, 4.933164, 4.930776, 4.929138, 4.928135, 4.927667, 
    4.927631, 4.927937, 4.928491, 4.9292, 4.92996, 4.930647, 4.931097, 
    4.931102, 4.930818, 4.946164, 4.943949, 4.940964, 4.937904, 4.934816, 
    4.936986, 4.938692, 4.94071, 4.939893, 4.93633, 4.929495, 4.919771, 
    4.907046, 4.894641, 4.882136, 4.8747, 4.867539, 4.861034, 4.855579, 
    4.851521, 4.849131, 4.84859, 4.849968, 4.853214, 4.858169, 4.864559, 
    4.872037, 4.88018, 4.888537, 4.896647, 4.90409, 4.910515, 4.915682, 
    4.919499,
  // momentumY(21,0, 0-49)
    4.867756, 4.87136, 4.876185, 4.881904, 4.888227, 4.894917, 4.901782, 
    4.908686, 4.915534, 4.922264, 4.928842, 4.935246, 4.941461, 4.947464, 
    4.953222, 4.958513, 4.964422, 4.96916, 4.973463, 4.977247, 4.98037, 
    4.982961, 4.984521, 4.984962, 4.984047, 4.981614, 4.977492, 4.971577, 
    4.963781, 4.95417, 4.942726, 4.929893, 4.915575, 4.900093, 4.883879, 
    4.867457, 4.851445, 4.836494, 4.823259, 4.812335, 4.804196, 4.799148, 
    4.797297, 4.798529, 4.802532, 4.808812, 4.816741, 4.82561, 4.834689, 
    4.843285,
  // momentumY(21,1, 0-49)
    4.869227, 4.873135, 4.878213, 4.88414, 4.890633, 4.897455, 4.904428, 
    4.911416, 4.918332, 4.925114, 4.931731, 4.938162, 4.944387, 4.950385, 
    4.956112, 4.961147, 4.967659, 4.972268, 4.976444, 4.980152, 4.983257, 
    4.986171, 4.988067, 4.988924, 4.988447, 4.98646, 4.982759, 4.977232, 
    4.969764, 4.960455, 4.949201, 4.93672, 4.922586, 4.907089, 4.890637, 
    4.87375, 4.857055, 4.841236, 4.827, 4.815002, 4.805791, 4.799745, 
    4.797029, 4.797587, 4.801143, 4.807224, 4.815208, 4.824379, 4.833981, 
    4.843285,
  // momentumY(21,2, 0-49)
    4.87042, 4.874584, 4.879874, 4.885972, 4.892601, 4.899534, 4.906593, 
    4.913648, 4.920613, 4.927431, 4.934066, 4.940497, 4.946706, 4.952666, 
    4.958333, 4.963048, 4.970029, 4.974471, 4.978471, 4.982044, 4.985077, 
    4.988253, 4.990441, 4.991687, 4.991656, 4.99017, 4.987002, 4.982033, 
    4.97512, 4.966384, 4.955632, 4.943846, 4.930265, 4.915128, 4.898799, 
    4.881767, 4.864641, 4.848114, 4.832927, 4.819794, 4.809337, 4.802019, 
    4.798089, 4.79757, 4.800246, 4.805697, 4.813336, 4.822461, 4.832316, 
    4.842153,
  // momentumY(21,3, 0-49)
    4.871417, 4.875794, 4.881257, 4.88749, 4.894225, 4.90124, 4.90836, 
    4.91546, 4.922452, 4.92928, 4.935906, 4.942309, 4.948469, 4.954359, 
    4.959938, 4.964278, 4.971559, 4.975809, 4.979591, 4.982981, 4.985889, 
    4.989264, 4.991691, 4.993279, 4.993685, 4.992729, 4.990175, 4.985899, 
    4.979735, 4.971802, 4.96182, 4.951028, 4.938334, 4.923909, 4.908056, 
    4.891205, 4.873922, 4.856891, 4.840857, 4.826586, 4.81477, 4.805964, 
    4.800524, 4.798568, 4.799973, 4.804396, 4.811304, 4.820037, 4.829866, 
    4.840038,
  // momentumY(21,4, 0-49)
    4.872332, 4.876885, 4.882481, 4.888814, 4.895623, 4.902688, 4.909839, 
    4.916954, 4.923941, 4.930746, 4.937329, 4.943668, 4.949744, 4.955535, 
    4.961005, 4.964917, 4.972301, 4.976346, 4.979885, 4.983051, 4.985792, 
    4.989301, 4.991906, 4.993781, 4.994592, 4.994171, 4.992283, 4.9888, 
    4.983535, 4.976586, 4.967588, 4.958031, 4.946498, 4.933095, 4.91804, 
    4.90169, 4.884544, 4.867239, 4.850518, 4.835167, 4.821952, 4.811521, 
    4.804342, 4.800659, 4.800459, 4.8035, 4.809333, 4.817359, 4.826887, 
    4.837183,
  // momentumY(21,5, 0-49)
    4.873298, 4.87799, 4.883683, 4.890078, 4.896924, 4.904002, 4.91115, 
    4.91824, 4.925184, 4.931925, 4.938425, 4.94466, 4.950615, 4.956275, 
    4.961616, 4.965065, 4.972339, 4.976171, 4.979454, 4.982371, 4.984913, 
    4.988491, 4.99121, 4.993308, 4.994482, 4.994578, 4.993377, 4.990749, 
    4.986489, 4.980652, 4.972798, 4.964639, 4.954481, 4.942347, 4.928371, 
    4.912815, 4.896089, 4.878769, 4.861557, 4.845256, 4.830675, 4.818562, 
    4.809506, 4.803884, 4.801821, 4.803196, 4.807662, 4.8147, 4.823673, 
    4.833878,
  // momentumY(21,6, 0-49)
    4.874443, 4.879241, 4.884993, 4.891414, 4.898254, 4.905306, 4.912405, 
    4.919427, 4.926284, 4.932917, 4.939289, 4.945377, 4.951174, 4.956671, 
    4.961865, 4.964837, 4.971784, 4.975398, 4.97842, 4.981078, 4.983403, 
    4.986985, 4.989758, 4.992006, 4.993488, 4.994068, 4.99355, 4.991801, 
    4.988611, 4.983963, 4.977353, 4.970687, 4.962039, 4.951355, 4.938675, 
    4.924161, 4.908125, 4.891047, 4.87358, 4.856506, 4.840674, 4.826908, 
    4.815924, 4.808243, 4.804142, 4.803638, 4.806506, 4.812325, 4.820523, 
    4.830435,
  // momentumY(21,7, 0-49)
    4.87588, 4.880752, 4.88653, 4.892937, 4.899731, 4.90671, 4.913714, 
    4.920619, 4.927339, 4.933815, 4.940012, 4.945911, 4.951509, 4.956812, 
    4.961838, 4.964347, 4.970757, 4.97415, 4.976916, 4.979318, 4.981421, 
    4.98495, 4.987716, 4.990044, 4.991772, 4.992788, 4.992926, 4.992055, 
    4.989957, 4.986527, 4.981206, 4.976059, 4.968983, 4.959855, 4.948626, 
    4.93535, 4.92023, 4.903647, 4.886172, 4.868548, 4.851635, 4.836328, 
    4.823456, 4.813686, 4.807459, 4.804945, 4.806056, 4.810474, 4.81771, 
    4.82715,
  // momentumY(21,8, 0-49)
    4.8777, 4.882618, 4.888388, 4.894741, 4.901444, 4.908303, 4.915162, 
    4.9219, 4.928433, 4.934703, 4.940678, 4.946343, 4.951704, 4.95678, 
    4.961609, 4.963711, 4.969393, 4.972557, 4.975082, 4.977241, 4.979133, 
    4.982553, 4.985257, 4.987593, 4.989506, 4.990901, 4.99165, 4.991627, 
    4.990613, 4.988391, 4.984363, 4.980696, 4.975188, 4.967651, 4.957954, 
    4.946052, 4.932031, 4.916164, 4.898924, 4.880996, 4.863228, 4.846558, 
    4.831919, 4.82012, 4.811763, 4.807185, 4.806442, 4.80934, 4.81547, 
    4.824277,
  // momentumY(21,9, 0-49)
    4.879959, 4.884899, 4.890628, 4.89689, 4.903462, 4.910154, 4.916817, 
    4.923337, 4.929632, 4.935648, 4.941355, 4.946746, 4.951833, 4.956645, 
    4.961241, 4.963027, 4.967825, 4.970748, 4.97305, 4.974993, 4.976692, 
    4.979956, 4.982547, 4.98483, 4.986863, 4.988575, 4.989882, 4.990657, 
    4.99069, 4.989635, 4.986869, 4.984592, 4.98059, 4.974617, 4.966471, 
    4.956012, 4.943221, 4.928251, 4.911475, 4.893493, 4.87512, 4.857318, 
    4.8411, 4.827405, 4.816993, 4.810369, 4.807745, 4.80905, 4.813972, 
    4.822018,
  // momentumY(21,10, 0-49)
    4.882683, 4.887622, 4.893283, 4.899419, 4.905817, 4.912298, 4.918719, 
    4.924973, 4.930984, 4.936702, 4.942099, 4.947176, 4.951952, 4.956465, 
    4.960778, 4.962388, 4.966177, 4.968843, 4.970945, 4.972705, 4.974249, 
    4.977313, 4.979748, 4.98192, 4.984013, 4.985978, 4.98778, 4.989291, 
    4.99031, 4.990362, 4.988803, 4.987789, 4.985182, 4.980694, 4.97406, 
    4.965057, 4.953567, 4.939633, 4.923513, 4.905717, 4.887003, 4.868331, 
    4.85077, 4.835371, 4.823044, 4.814457, 4.809978, 4.809673, 4.813326, 
    4.820508,
  // momentumY(21,11, 0-49)
    4.885859, 4.890782, 4.896351, 4.902331, 4.90852, 4.914749, 4.920887, 
    4.926834, 4.932517, 4.937896, 4.942946, 4.947676, 4.952104, 4.956275, 
    4.960248, 4.961854, 4.964558, 4.966954, 4.968882, 4.970501, 4.971934, 
    4.974759, 4.977002, 4.979015, 4.981116, 4.983275, 4.985504, 4.987677, 
    4.989609, 4.990688, 4.990268, 4.990361, 4.989007, 4.985883, 4.980674, 
    4.973091, 4.962924, 4.950112, 4.934801, 4.917403, 4.898602, 4.879333, 
    4.860695, 4.843828, 4.829777, 4.819361, 4.813109, 4.811215, 4.813574, 
    4.819819,
  // momentumY(21,12, 0-49)
    4.88944, 4.894337, 4.899799, 4.905598, 4.911548, 4.917494, 4.923313, 
    4.928915, 4.934238, 4.939242, 4.943916, 4.948267, 4.952316, 4.956103, 
    4.959673, 4.961469, 4.963051, 4.965169, 4.966954, 4.968485, 4.96986, 
    4.972414, 4.974438, 4.976257, 4.978319, 4.980617, 4.983204, 4.985958, 
    4.988717, 4.990734, 4.99138, 4.99241, 4.992143, 4.990234, 4.986331, 
    4.980086, 4.971216, 4.959564, 4.945173, 4.928348, 4.909691, 4.890091, 
    4.870652, 4.852578, 4.837027, 4.824958, 4.81705, 4.813632, 4.814701, 
    4.819964,
  // momentumY(21,13, 0-49)
    4.893345, 4.898217, 4.90356, 4.909164, 4.914856, 4.920492, 4.925966, 
    4.931196, 4.936131, 4.94074, 4.945012, 4.948959, 4.952602, 4.955966, 
    4.959073, 4.961245, 4.961709, 4.963559, 4.96524, 4.96674, 4.96812, 
    4.970376, 4.972166, 4.973768, 4.975757, 4.978142, 4.981021, 4.984272, 
    4.987758, 4.990619, 4.99226, 4.994047, 4.99469, 4.993832, 4.991089, 
    4.98607, 4.978432, 4.967936, 4.954527, 4.93841, 4.920095, 4.900408, 
    4.880437, 4.861424, 4.844614, 4.831095, 4.821679, 4.816827, 4.816639, 
    4.820898,
  // momentumY(21,14, 0-49)
    4.897468, 4.902321, 4.907547, 4.912951, 4.918373, 4.923688, 4.928799, 
    4.93364, 4.93817, 4.942365, 4.946223, 4.949754, 4.95297, 4.95588, 
    4.958479, 4.961169, 4.960548, 4.962161, 4.963795, 4.965333, 4.966787, 
    4.968728, 4.97028, 4.971656, 4.973548, 4.975982, 4.979085, 4.982744, 
    4.986854, 4.990458, 4.993018, 4.995389, 4.996763, 4.99678, 4.995036, 
    4.991111, 4.98461, 4.975227, 4.962822, 4.947505, 4.929689, 4.910128, 
    4.889874, 4.870183, 4.852361, 4.837605, 4.826849, 4.820671, 4.819281, 
    4.822535,
  // momentumY(21,15, 0-49)
    4.901683, 4.906533, 4.911652, 4.916859, 4.922011, 4.927, 4.931743, 
    4.936191, 4.94031, 4.944088, 4.94753, 4.950641, 4.953424, 4.955871, 
    4.957943, 4.96121, 4.959546, 4.960984, 4.962644, 4.9643, 4.965909, 
    4.967529, 4.968853, 4.970014, 4.971802, 4.974249, 4.977513, 4.981489, 
    4.986113, 4.990354, 4.993762, 4.996544, 4.998473, 4.999189, 4.998278, 
    4.995298, 4.989818, 4.981478, 4.970063, 4.955593, 4.938392, 4.919131, 
    4.898813, 4.878683, 4.860091, 4.844313, 4.832389, 4.825014, 4.822492, 
    4.824755,
  // momentumY(21,16, 0-49)
    4.905852, 4.910719, 4.915746, 4.92077, 4.925663, 4.930331, 4.934713, 
    4.938773, 4.942492, 4.945868, 4.948905, 4.951612, 4.953979, 4.955981, 
    4.95755, 4.961321, 4.958642, 4.960001, 4.961782, 4.963653, 4.965511, 
    4.966817, 4.967943, 4.968918, 4.970611, 4.973051, 4.976418, 4.980618, 
    4.985636, 4.9904, 4.994579, 4.99761, 4.999923, 5.001165, 5.00092, 
    4.99873, 4.994142, 4.986749, 4.976277, 4.962667, 4.946156, 4.927331, 
    4.907132, 4.886779, 4.86764, 4.851046, 4.838132, 4.82969, 4.826118, 
    4.82742,
  // momentumY(21,17, 0-49)
    4.909837, 4.914738, 4.919692, 4.924548, 4.929195, 4.93356, 4.9376, 
    4.941293, 4.944641, 4.947648, 4.950324, 4.95267, 4.954671, 4.956281, 
    4.957415, 4.961463, 4.957752, 4.959157, 4.961174, 4.963372, 4.965584, 
    4.966605, 4.967587, 4.968428, 4.970053, 4.97248, 4.975895, 4.980227, 
    4.985517, 4.99068, 4.995541, 4.998661, 5.001194, 5.002797, 5.003052, 
    5.001498, 4.997662, 4.991107, 4.98151, 4.968741, 4.95296, 4.934667, 
    4.914736, 4.894343, 4.874856, 4.857644, 4.843911, 4.834536, 4.83, 4.830382,
  // momentumY(21,18, 0-49)
    4.913497, 4.918441, 4.923331, 4.928032, 4.932451, 4.936535, 4.940263, 
    4.943635, 4.946665, 4.949371, 4.951762, 4.953833, 4.955557, 4.956873, 
    4.957686, 4.961622, 4.956789, 4.958377, 4.96076, 4.963412, 4.9661, 
    4.966885, 4.967799, 4.968584, 4.970194, 4.972615, 4.97604, 4.980412, 
    4.985839, 4.991264, 4.996696, 4.999753, 5.002348, 5.004149, 5.004743, 
    5.003669, 5.000443, 4.994608, 4.985798, 4.973829, 4.958785, 4.94109, 
    4.921543, 4.901266, 4.881607, 4.863956, 4.849568, 4.839391, 4.833985, 
    4.833497,
  // momentumY(21,19, 0-49)
    4.9167, 4.921665, 4.926477, 4.931019, 4.93522, 4.939054, 4.942522, 
    4.945646, 4.948455, 4.950972, 4.953205, 4.955136, 4.956722, 4.957885, 
    4.958528, 4.961836, 4.95568, 4.957586, 4.960464, 4.963702, 4.967002, 
    4.967633, 4.968585, 4.96942, 4.971097, 4.973547, 4.976954, 4.981276, 
    4.986701, 4.992226, 4.998084, 5.00092, 5.003414, 5.00525, 5.006023, 
    5.005275, 5.00252, 4.997281, 4.989166, 4.977938, 4.963619, 4.94656, 
    4.927482, 4.90745, 4.887774, 4.869849, 4.854956, 4.84411, 4.837931, 
    4.836633,
  // momentumY(21,20, 0-49)
    4.920373, 4.926408, 4.932198, 4.937615, 4.942574, 4.947017, 4.95092, 
    4.954266, 4.957061, 4.959322, 4.961086, 4.962402, 4.963344, 4.963996, 
    4.96446, 0, 4.958336, 4.959911, 4.962055, 4.964373, 4.966731, 4.965669, 
    4.965298, 4.965133, 4.966242, 4.968559, 4.972223, 4.977122, 4.983384, 
    4.989923, 4.997092, 5.000469, 5.003476, 5.005798, 5.007044, 5.006776, 
    5.004527, 4.999839, 4.992319, 4.981717, 4.96802, 4.951524, 4.932887, 
    4.913119, 4.893489, 4.875374, 4.860076, 4.848648, 4.841766, 4.839701,
  // momentumY(21,21, 0-49)
    4.922716, 4.928973, 4.934875, 4.9403, 4.945176, 4.949471, 4.95318, 
    4.956317, 4.958914, 4.96101, 4.962654, 4.963908, 4.964848, 4.965567, 
    4.966182, 0, 4.955145, 4.957202, 4.959885, 4.962759, 4.965636, 4.964164, 
    4.963536, 4.963161, 4.964198, 4.966575, 4.970424, 4.975614, 4.982278, 
    4.989311, 4.997245, 5.000715, 5.003937, 5.006592, 5.008276, 5.008539, 
    5.006902, 5.002893, 4.996096, 4.986228, 4.97323, 4.957343, 4.939162, 
    4.919639, 4.900001, 4.881614, 4.865797, 4.85364, 4.845881, 4.842846,
  // momentumY(21,22, 0-49)
    4.924577, 4.931123, 4.937216, 4.942735, 4.947618, 4.951845, 4.955435, 
    4.958422, 4.960857, 4.962803, 4.964324, 4.965492, 4.966395, 4.967139, 
    4.967857, 0, 4.952854, 4.955309, 4.958461, 4.96184, 4.965202, 4.963355, 
    4.962503, 4.961944, 4.962914, 4.96533, 4.96931, 4.974701, 4.981636, 
    4.988995, 4.997468, 5.000855, 5.004099, 5.006884, 5.008801, 5.009401, 
    5.008202, 5.004722, 4.998529, 4.989316, 4.976982, 4.961714, 4.944051, 
    4.92488, 4.905382, 4.886895, 4.870741, 4.858034, 4.849556, 4.845685,
  // momentumY(21,23, 0-49)
    4.925975, 4.932854, 4.939191, 4.944864, 4.949818, 4.954044, 4.957575, 
    4.960462, 4.962778, 4.964598, 4.966004, 4.967083, 4.967932, 4.968668, 
    4.969452, 0, 4.951511, 4.954235, 4.957705, 4.961428, 4.965119, 4.962908, 
    4.961822, 4.961064, 4.961936, 4.964339, 4.968385, 4.973899, 4.98101, 
    4.988581, 4.997424, 5.000678, 5.003872, 5.006702, 5.008762, 5.009603, 
    5.008744, 5.0057, 5.000029, 4.9914, 4.97968, 4.96501, 4.947873, 4.929098, 
    4.909818, 4.891339, 4.874972, 4.861847, 4.852779, 4.848183,
  // momentumY(21,24, 0-49)
    4.926955, 4.934186, 4.940796, 4.946662, 4.951729, 4.956, 4.959518, 
    4.962349, 4.964579, 4.966302, 4.96761, 4.968601, 4.969385, 4.970094, 
    4.970906, 0, 4.951337, 4.954191, 4.957818, 4.961719, 4.965586, 4.963124, 
    4.961879, 4.96099, 4.961792, 4.964177, 4.968248, 4.973822, 4.981027, 
    4.988714, 4.997774, 5.000921, 5.004061, 5.006891, 5.009009, 5.009973, 
    5.009304, 5.006517, 5.001168, 4.992916, 4.981607, 4.967354, 4.950599, 
    4.932136, 4.913054, 4.894632, 4.878164, 4.864782, 4.855316, 4.850201,
  // momentumY(21,25, 0-49)
    4.927581, 4.93516, 4.94205, 4.948121, 4.953326, 4.957671, 4.961206, 
    4.964014, 4.96619, 4.967835, 4.969058, 4.969966, 4.970678, 4.971337, 
    4.972132, 0, 4.951993, 4.954841, 4.958466, 4.962369, 4.966248, 4.963695, 
    4.962402, 4.961487, 4.962284, 4.964675, 4.968763, 4.974359, 4.981592, 
    4.989312, 4.998431, 5.001542, 5.004662, 5.007491, 5.009628, 5.010636, 
    5.010038, 5.007354, 5.002141, 4.994059, 4.982945, 4.968903, 4.952358, 
    4.934081, 4.915137, 4.896785, 4.880301, 4.866809, 4.857136, 4.851721,
  // momentumY(21,26, 0-49)
    4.927925, 4.935825, 4.942978, 4.949254, 4.954605, 4.959037, 4.962613, 
    4.965418, 4.967557, 4.969142, 4.970285, 4.971105, 4.971728, 4.972306, 
    4.973034, 0, 4.953425, 4.95613, 4.959591, 4.963326, 4.96705, 4.964577, 
    4.963362, 4.962536, 4.963402, 4.965837, 4.969944, 4.975535, 4.982742, 
    4.990416, 4.999442, 5.002605, 5.005761, 5.008602, 5.010732, 5.011711, 
    5.011069, 5.008329, 5.003057, 4.994917, 4.983764, 4.969701, 4.953165, 
    4.934923, 4.91604, 4.89776, 4.881342, 4.867894, 4.858222, 4.852753,
  // momentumY(21,27, 0-49)
    4.92806, 4.936237, 4.943624, 4.950087, 4.955577, 4.960105, 4.963733, 
    4.96655, 4.968665, 4.970191, 4.971249, 4.971961, 4.972464, 4.972912, 
    4.973501, 0, 4.955719, 4.958138, 4.961273, 4.964661, 4.968061, 4.965804, 
    4.964757, 4.964105, 4.965088, 4.967585, 4.971696, 4.977244, 4.98436, 
    4.99191, 5.000689, 5.003982, 5.007212, 5.01007, 5.012156, 5.013031, 
    5.01223, 5.009284, 5.00377, 4.995371, 4.983961, 4.969677, 4.952976, 
    4.93465, 4.915774, 4.897588, 4.881337, 4.868097, 4.85864, 4.853362,
  // momentumY(21,28, 0-49)
    4.928054, 4.936454, 4.944035, 4.950661, 4.956285, 4.960913, 4.964603, 
    4.967442, 4.969531, 4.970989, 4.971935, 4.972499, 4.972823, 4.973068, 
    4.973427, 0, 4.959241, 4.961226, 4.963868, 4.966732, 4.969642, 4.967668, 
    4.96682, 4.966366, 4.967466, 4.969997, 4.974066, 4.979512, 4.986459, 
    4.993795, 5.002191, 5.005653, 5.008963, 5.011804, 5.013775, 5.014439, 
    5.013337, 5.010012, 5.004061, 4.995199, 4.983335, 4.968651, 4.951647, 
    4.933157, 4.914279, 4.896254, 4.880302, 4.867464, 4.858457, 4.853627,
  // momentumY(21,29, 0-49)
    4.92797, 4.936532, 4.944271, 4.951048, 4.956806, 4.961545, 4.965309, 
    4.968172, 4.970227, 4.971584, 4.972364, 4.972703, 4.972755, 4.972694, 
    4.972711, 0, 4.963769, 4.965175, 4.967158, 4.969325, 4.971568, 4.96982, 
    4.969094, 4.968768, 4.969911, 4.972406, 4.976363, 4.981632, 4.988328, 
    4.995357, 5.003223, 5.006826, 5.010169, 5.01293, 5.014711, 5.015079, 
    5.013591, 5.0098, 5.003335, 4.99394, 4.981572, 4.966462, 4.949168, 
    4.930563, 4.911772, 4.894035, 4.878546, 4.866288, 4.85792, 4.853728,
  // momentumY(21,30, 0-49)
    4.926956, 4.934618, 4.941468, 4.947391, 4.952364, 4.956439, 4.959708, 
    4.962296, 4.964333, 4.965935, 4.967184, 4.968123, 4.968738, 4.968968, 
    4.968709, 4.975595, 4.962874, 4.964472, 4.967275, 4.970613, 4.974156, 
    4.97453, 4.975579, 4.976661, 4.978667, 4.98145, 4.985137, 4.989669, 
    4.995262, 5.000958, 5.007199, 5.009936, 5.012409, 5.014312, 5.015257, 
    5.014821, 5.012557, 5.008026, 5.000863, 4.990838, 4.977942, 4.962452, 
    4.944969, 4.926406, 4.9079, 4.890683, 4.875904, 4.864484, 4.857009, 
    4.853695,
  // momentumY(21,31, 0-49)
    4.926929, 4.934672, 4.941601, 4.947601, 4.95264, 4.956754, 4.960025, 
    4.962573, 4.964523, 4.965997, 4.967094, 4.96788, 4.968374, 4.968542, 
    4.968293, 4.975252, 4.964764, 4.96593, 4.968161, 4.970851, 4.97374, 
    4.974269, 4.975286, 4.976324, 4.978278, 4.981052, 4.98479, 4.98941, 
    4.995051, 5.0007, 5.006574, 5.009628, 5.012319, 5.014328, 5.015259, 
    5.014685, 5.012158, 5.007254, 4.999632, 4.989102, 4.975713, 4.959807, 
    4.942053, 4.923415, 4.905064, 4.888221, 4.874006, 4.863276, 4.856546, 
    4.853962,
  // momentumY(21,32, 0-49)
    4.926838, 4.934477, 4.941327, 4.947276, 4.952287, 4.956389, 4.959658, 
    4.962198, 4.964133, 4.965584, 4.966657, 4.967435, 4.967957, 4.968214, 
    4.968139, 4.974419, 4.966065, 4.966943, 4.968725, 4.970888, 4.973237, 
    4.974019, 4.975111, 4.976216, 4.978195, 4.980991, 4.984751, 4.989377, 
    4.994931, 5.000389, 5.005764, 5.009021, 5.011818, 5.013818, 5.014621, 
    5.013795, 5.0109, 5.005525, 4.997361, 4.986272, 4.972367, 4.956063, 
    4.938097, 4.919488, 4.901426, 4.885119, 4.871639, 4.861775, 4.855964, 
    4.854273,
  // momentumY(21,33, 0-49)
    4.926754, 4.934147, 4.940796, 4.946594, 4.951506, 4.955551, 4.958797, 
    4.961343, 4.963299, 4.964785, 4.96591, 4.966764, 4.967407, 4.967854, 
    4.968068, 4.973201, 4.966861, 4.967598, 4.969047, 4.970792, 4.972705, 
    4.973806, 4.97506, 4.976316, 4.978374, 4.981203, 4.984944, 4.989483, 
    4.994825, 4.999962, 5.004738, 5.008092, 5.010881, 5.012757, 5.013318, 
    5.012129, 5.00876, 5.002823, 4.994051, 4.982362, 4.967942, 4.951282, 
    4.93319, 4.914731, 4.897108, 4.881502, 4.868926, 4.86009, 4.855348, 
    4.854691,
  // momentumY(21,34, 0-49)
    4.926736, 4.933774, 4.940129, 4.945702, 4.950455, 4.954404, 4.95761, 
    4.960158, 4.962151, 4.9637, 4.964916, 4.96589, 4.966699, 4.967385, 
    4.967942, 4.971733, 4.967276, 4.967985, 4.969195, 4.970612, 4.972173, 
    4.973621, 4.975093, 4.976563, 4.978733, 4.98159, 4.98526, 4.989622, 
    4.994627, 4.999331, 5.003438, 5.006778, 5.009446, 5.011085, 5.011292, 
    5.009635, 5.005699, 4.999127, 4.989699, 4.977401, 4.962496, 4.945557, 
    4.927455, 4.909292, 4.892269, 4.877531, 4.866017, 4.858353, 4.854806, 
    4.855289,
  // momentumY(21,35, 0-49)
    4.926836, 4.933433, 4.939422, 4.944709, 4.949258, 4.953081, 4.956228, 
    4.95877, 4.960804, 4.96243, 4.96375, 4.964861, 4.965849, 4.966776, 
    4.967676, 4.970145, 4.967444, 4.968202, 4.969242, 4.970393, 4.971665, 
    4.973465, 4.975183, 4.976903, 4.979197, 4.982062, 4.985603, 4.989695, 
    4.994246, 4.998414, 5.001794, 5.005006, 5.007436, 5.008721, 5.008463, 
    5.00624, 5.001657, 4.994396, 4.984295, 4.971416, 4.9561, 4.938995, 
    4.921033, 4.903339, 4.887095, 4.873391, 4.863085, 4.856715, 4.854457, 
    4.856152,
  // momentumY(21,36, 0-49)
    4.927101, 4.933189, 4.938755, 4.943709, 4.948019, 4.951687, 4.954755, 
    4.957284, 4.959356, 4.961058, 4.962487, 4.963735, 4.964891, 4.966037, 
    4.967238, 4.96855, 4.967488, 4.968328, 4.969235, 4.970166, 4.9712, 
    4.973329, 4.975299, 4.977283, 4.979695, 4.982537, 4.985882, 4.989611, 
    4.993591, 4.997127, 4.999732, 5.00269, 5.004757, 5.005571, 5.00474, 
    5.00186, 4.996566, 4.988592, 4.977838, 4.964443, 4.948833, 4.931724, 
    4.91409, 4.897061, 4.881786, 4.869282, 4.860319, 4.855337, 4.85443, 
    4.857368,
  // momentumY(21,37, 0-49)
    4.927572, 4.933101, 4.938197, 4.942782, 4.946818, 4.950309, 4.95328, 
    4.955783, 4.957885, 4.959661, 4.961193, 4.962566, 4.963869, 4.965193, 
    4.966624, 4.967034, 4.967501, 4.96842, 4.969209, 4.969953, 4.970782, 
    4.9732, 4.975408, 4.97765, 4.980156, 4.982931, 4.986008, 4.989279, 
    4.992575, 4.995385, 4.997163, 4.999734, 5.00131, 5.001532, 5.000024, 
    4.996412, 4.990367, 4.981685, 4.970336, 4.956542, 4.940803, 4.923894, 
    4.906811, 4.890669, 4.876559, 4.865418, 4.857912, 4.854388, 4.854856, 
    4.859026,
  // momentumY(21,38, 0-49)
    4.928286, 4.933214, 4.937806, 4.941989, 4.945725, 4.949013, 4.951869, 
    4.954332, 4.956453, 4.95829, 4.959915, 4.9614, 4.962823, 4.964279, 
    4.965862, 4.965644, 4.967535, 4.968503, 4.969175, 4.969752, 4.970407, 
    4.97306, 4.975472, 4.977946, 4.980508, 4.983161, 4.985892, 4.988606, 
    4.991111, 4.993099, 4.993998, 4.996039, 4.99699, 4.996502, 4.994226, 
    4.989821, 4.983016, 4.97367, 4.961834, 4.947803, 4.932146, 4.915679, 
    4.899399, 4.884381, 4.87164, 4.86201, 4.856055, 4.854027, 4.85586, 
    4.861211,
  // momentumY(21,39, 0-49)
    4.929265, 4.933565, 4.937625, 4.941379, 4.944791, 4.947852, 4.950571, 
    4.952974, 4.955095, 4.95698, 4.958681, 4.960257, 4.961775, 4.963317, 
    4.964976, 4.964395, 4.967595, 4.96857, 4.969121, 4.969549, 4.97005, 
    4.972878, 4.975447, 4.978108, 4.980676, 4.983141, 4.985444, 4.987503, 
    4.989108, 4.990186, 4.990143, 4.991511, 4.991702, 4.990395, 4.987274, 
    4.982047, 4.974504, 4.964581, 4.952405, 4.938348, 4.923028, 4.907279, 
    4.892075, 4.878423, 4.867244, 4.859259, 4.854925, 4.8544, 4.857553, 
    4.863996,
  // momentumY(21,40, 0-49)
    4.930509, 4.934163, 4.937672, 4.940976, 4.944041, 4.946851, 4.949409, 
    4.951728, 4.953829, 4.95574, 4.957498, 4.959143, 4.96073, 4.962318, 
    4.963991, 4.96327, 4.967656, 4.968591, 4.969017, 4.969309, 4.969671, 
    4.972606, 4.975278, 4.97807, 4.980577, 4.982781, 4.984569, 4.985875, 
    4.986485, 4.986562, 4.985514, 4.986065, 4.985376, 4.983157, 4.979137, 
    4.973087, 4.964869, 4.954496, 4.942178, 4.928343, 4.913644, 4.898909, 
    4.885057, 4.873009, 4.86357, 4.857339, 4.854666, 4.855622, 4.860014, 
    4.867422,
  // momentumY(21,41, 0-49)
    4.931998, 4.934996, 4.937942, 4.94078, 4.943478, 4.946014, 4.948385, 
    4.950592, 4.952645, 4.954556, 4.956345, 4.958038, 4.959667, 4.961271, 
    4.962908, 4.962221, 4.967657, 4.968509, 4.968806, 4.968975, 4.969211, 
    4.972187, 4.974899, 4.977754, 4.980126, 4.981987, 4.983173, 4.983639, 
    4.983162, 4.982157, 4.980039, 4.979643, 4.977969, 4.974769, 4.969831, 
    4.962996, 4.954207, 4.943558, 4.931327, 4.917993, 4.904217, 4.890792, 
    4.878562, 4.868335, 4.860787, 4.856392, 4.855388, 4.857768, 4.863286, 
    4.8715,
  // momentumY(21,42, 0-49)
    4.933681, 4.93602, 4.938399, 4.940762, 4.943074, 4.945315, 4.947473, 
    4.949539, 4.951512, 4.953393, 4.955186, 4.9569, 4.958545, 4.960138, 
    4.961708, 4.961169, 4.967508, 4.968248, 4.968419, 4.968473, 4.968589, 
    4.971543, 4.97423, 4.977072, 4.979232, 4.980669, 4.981169, 4.980713, 
    4.979079, 4.976922, 4.973677, 4.972228, 4.969491, 4.965276, 4.95944, 
    4.951901, 4.942686, 4.931967, 4.920083, 4.907539, 4.894986, 4.883152, 
    4.872786, 4.864562, 4.859018, 4.856503, 4.857143, 4.860859, 4.867363, 
    4.876194,
  // momentumY(21,43, 0-49)
    4.935478, 4.937166, 4.938977, 4.940857, 4.942774, 4.9447, 4.946618, 
    4.948514, 4.950376, 4.952195, 4.953959, 4.955664, 4.957301, 4.958864, 
    4.960346, 4.960024, 4.967107, 4.967718, 4.967767, 4.967717, 4.967713, 
    4.970584, 4.973182, 4.975931, 4.977798, 4.978734, 4.978477, 4.977031, 
    4.974191, 4.970835, 4.966425, 4.963848, 4.960012, 4.95479, 4.948117, 
    4.939998, 4.930539, 4.919984, 4.908716, 4.897247, 4.886191, 4.876195, 
    4.867887, 4.861801, 4.858331, 4.857696, 4.859924, 4.86486, 4.87218, 
    4.88142,
  // momentumY(21,44, 0-49)
    4.937275, 4.938323, 4.939574, 4.940974, 4.942487, 4.944084, 4.945742, 
    4.947441, 4.949162, 4.950884, 4.95259, 4.954257, 4.955863, 4.957377, 
    4.958764, 4.958681, 4.966344, 4.966816, 4.966756, 4.966607, 4.966479, 
    4.969213, 4.971659, 4.974236, 4.975735, 4.976098, 4.975027, 4.972552, 
    4.968484, 4.96391, 4.958328, 4.954591, 4.949665, 4.943493, 4.936093, 
    4.927554, 4.91806, 4.907915, 4.897525, 4.887393, 4.878069, 4.8701, 
    4.863985, 4.860114, 4.858732, 4.859934, 4.863651, 4.869663, 4.877614, 
    4.887039,
  // momentumY(21,45, 0-49)
    4.938926, 4.939353, 4.940056, 4.940982, 4.942094, 4.943354, 4.944736, 
    4.946219, 4.947771, 4.949369, 4.950988, 4.952592, 4.954145, 4.955598, 
    4.956888, 4.957033, 4.965114, 4.965453, 4.965286, 4.965036, 4.964778, 
    4.967328, 4.969562, 4.97189, 4.972956, 4.972693, 4.970773, 4.967258, 
    4.961981, 4.956205, 4.949481, 4.944608, 4.938652, 4.931637, 4.923662, 
    4.914896, 4.905593, 4.896097, 4.886826, 4.878241, 4.870824, 4.865007, 
    4.861149, 4.859497, 4.860159, 4.863107, 4.868181, 4.875099, 4.883481, 
    4.892863,
  // momentumY(21,46, 0-49)
    4.940262, 4.940084, 4.940259, 4.940728, 4.941444, 4.942371, 4.943476, 
    4.944729, 4.946098, 4.947554, 4.949063, 4.950583, 4.952066, 4.953447, 
    4.954642, 4.95498, 4.963323, 4.963535, 4.963268, 4.96291, 4.962506, 
    4.964828, 4.9668, 4.968812, 4.969393, 4.968471, 4.965699, 4.961167, 
    4.954741, 4.947829, 4.940039, 4.934107, 4.927235, 4.919528, 4.911165, 
    4.902386, 4.893498, 4.884871, 4.876911, 4.870032, 4.864622, 4.861, 
    4.859388, 4.859892, 4.862491, 4.867044, 4.873307, 4.880941, 4.889546, 
    4.898666,
  // momentumY(21,47, 0-49)
    4.941096, 4.940332, 4.939998, 4.940029, 4.940372, 4.940979, 4.941815, 
    4.942842, 4.944026, 4.945332, 4.94672, 4.948144, 4.949549, 4.950854, 
    4.951961, 4.952435, 4.960899, 4.960996, 4.960621, 4.960141, 4.959572, 
    4.961631, 4.963296, 4.964937, 4.965001, 4.963412, 4.959817, 4.954334, 
    4.946867, 4.938931, 4.930195, 4.923338, 4.915718, 4.907512, 4.898972, 
    4.890397, 4.882132, 4.874554, 4.868045, 4.862955, 4.859578, 4.858113, 
    4.858655, 4.861183, 4.865554, 4.871528, 4.878778, 4.886925, 4.895541, 
    4.904192,
  // momentumY(21,48, 0-49)
    4.941243, 4.939906, 4.939085, 4.938703, 4.938699, 4.939013, 4.939602, 
    4.940422, 4.941435, 4.942599, 4.943874, 4.945204, 4.946529, 4.947761, 
    4.948786, 4.949333, 4.957789, 4.957774, 4.957283, 4.956659, 4.955901, 
    4.95767, 4.958993, 4.960226, 4.959764, 4.95753, 4.953178, 4.946849, 
    4.938492, 4.929691, 4.920184, 4.91259, 4.904428, 4.895942, 4.887444, 
    4.879278, 4.871814, 4.865419, 4.860435, 4.857142, 4.855741, 4.856319, 
    4.858856, 4.863209, 4.869135, 4.876301, 4.884318, 4.892757, 4.901187, 
    4.909195,
  // momentumY(21,49, 0-49)
    4.941844, 4.93949, 4.937799, 4.936679, 4.936049, 4.935833, 4.935967, 
    4.936391, 4.937048, 4.937884, 4.938838, 4.939832, 4.94078, 4.941552, 
    4.941981, 4.941836, 4.957452, 4.955976, 4.953788, 4.951624, 4.94955, 
    4.952877, 4.955788, 4.959049, 4.959525, 4.957204, 4.951482, 4.942688, 
    4.930685, 4.918662, 4.906098, 4.898111, 4.889776, 4.881432, 4.873471, 
    4.866293, 4.860284, 4.855782, 4.853061, 4.852297, 4.853556, 4.856781, 
    4.861804, 4.868344, 4.876037, 4.88445, 4.893135, 4.901632, 4.909525, 
    4.916467,
  // momentumY(22,0, 0-49)
    4.880537, 4.886049, 4.892055, 4.89834, 4.90474, 4.911143, 4.917471, 
    4.923685, 4.92976, 4.935697, 4.941501, 4.947173, 4.952713, 4.958113, 
    4.963342, 4.968148, 4.973527, 4.977929, 4.981947, 4.985516, 4.988526, 
    4.991129, 4.992905, 4.993828, 4.99375, 4.992583, 4.990228, 4.986621, 
    4.981689, 4.975449, 4.967793, 4.959002, 4.948776, 4.937156, 4.924249, 
    4.910238, 4.895406, 4.880136, 4.864914, 4.850298, 4.836879, 4.825234, 
    4.815861, 4.809134, 4.805259, 4.804258, 4.805966, 4.810053, 4.816054, 
    4.823408,
  // momentumY(22,1, 0-49)
    4.881404, 4.887128, 4.893311, 4.899741, 4.906262, 4.912758, 4.919157, 
    4.925417, 4.93152, 4.937462, 4.943248, 4.948881, 4.954358, 4.959669, 
    4.964782, 4.969224, 4.975, 4.979175, 4.982958, 4.986339, 4.989226, 
    4.992044, 4.994077, 4.995368, 4.995728, 4.995061, 4.993247, 4.99022, 
    4.985889, 4.980306, 4.973286, 4.96537, 4.95594, 4.94499, 4.932577, 
    4.918843, 4.904028, 4.888497, 4.872729, 4.857299, 4.842846, 4.830007, 
    4.819363, 4.81137, 4.806323, 4.804312, 4.805237, 4.808805, 4.814574, 
    4.821985,
  // momentumY(22,2, 0-49)
    4.882138, 4.888039, 4.894367, 4.900916, 4.907531, 4.914097, 4.920544, 
    4.926829, 4.932936, 4.938857, 4.944596, 4.950159, 4.955542, 4.960733, 
    4.965704, 4.969741, 4.975807, 4.979735, 4.983255, 4.986413, 4.989146, 
    4.992136, 4.994386, 4.996001, 4.99677, 4.996595, 4.995338, 4.992937, 
    4.989284, 4.984453, 4.978187, 4.971295, 4.962846, 4.952787, 4.941124, 
    4.927945, 4.913436, 4.897918, 4.881842, 4.865784, 4.850403, 4.836392, 
    4.824409, 4.815003, 4.808563, 4.805276, 4.805117, 4.807853, 4.813084, 
    4.820271,
  // momentumY(22,3, 0-49)
    4.88286, 4.888899, 4.895341, 4.901977, 4.908658, 4.915267, 4.921736, 
    4.92802, 4.9341, 4.93997, 4.945633, 4.951095, 4.956351, 4.961398, 
    4.966206, 4.969803, 4.976026, 4.979697, 4.982938, 4.98585, 4.988398, 
    4.991513, 4.99393, 4.995817, 4.996953, 4.997241, 4.996539, 4.994784, 
    4.991858, 4.987838, 4.982406, 4.976634, 4.969298, 4.960302, 4.949604, 
    4.937222, 4.923286, 4.908053, 4.891929, 4.875461, 4.859316, 4.844221, 
    4.830904, 4.820007, 4.812023, 4.807248, 4.80575, 4.807377, 4.811787, 
    4.818478,
  // momentumY(22,4, 0-49)
    4.883684, 4.889828, 4.896346, 4.903038, 4.90975, 4.916372, 4.922831, 
    4.929082, 4.935105, 4.940893, 4.946448, 4.951777, 4.956883, 4.96176, 
    4.966392, 4.969527, 4.975749, 4.97916, 4.982116, 4.984766, 4.987107, 
    4.990293, 4.992825, 4.99492, 4.996367, 4.997078, 4.996912, 4.995807, 
    4.993631, 4.990452, 4.985897, 4.981287, 4.975144, 4.96733, 4.957751, 
    4.94637, 4.93324, 4.918549, 4.902637, 4.886006, 4.869302, 4.853272, 
    4.838696, 4.826305, 4.8167, 4.810288, 4.807254, 4.807538, 4.810874, 
    4.816814,
  // momentumY(22,5, 0-49)
    4.884719, 4.890928, 4.897486, 4.904196, 4.910906, 4.917505, 4.92392, 
    4.930103, 4.936036, 4.941709, 4.947129, 4.952298, 4.957226, 4.961914, 
    4.96636, 4.969028, 4.97508, 4.978233, 4.980904, 4.983284, 4.985404, 
    4.98861, 4.991196, 4.993429, 4.995127, 4.99621, 4.996547, 4.996074, 
    4.994657, 4.992321, 4.988653, 4.985206, 4.980282, 4.973714, 4.96536, 
    4.955123, 4.942988, 4.929064, 4.913613, 4.897071, 4.880046, 4.86328, 
    4.847586, 4.833769, 4.822536, 4.814412, 4.809701, 4.80846, 4.81051, 
    4.815478,
  // momentumY(22,6, 0-49)
    4.886049, 4.892287, 4.898846, 4.905535, 4.912204, 4.918742, 4.925076, 
    4.931158, 4.936968, 4.942498, 4.947752, 4.952737, 4.957466, 4.961949, 
    4.9662, 4.968412, 4.974121, 4.97702, 4.979414, 4.981527, 4.983417, 
    4.986587, 4.98917, 4.991468, 4.99335, 4.994747, 4.995544, 4.99568, 
    4.995009, 4.993502, 4.990707, 4.988382, 4.984662, 4.979352, 4.972273, 
    4.963274, 4.952274, 4.9393, 4.924531, 4.908326, 4.89123, 4.873957, 
    4.857336, 4.842224, 4.829421, 4.819574, 4.813116, 4.810222, 4.810823, 
    4.814631,
  // momentumY(22,7, 0-49)
    4.887733, 4.893962, 4.900485, 4.907114, 4.913703, 4.920143, 4.92636, 
    4.932308, 4.937963, 4.94332, 4.948382, 4.953161, 4.957674, 4.961939, 
    4.965983, 4.967781, 4.972977, 4.975623, 4.977752, 4.979605, 4.981266, 
    4.984348, 4.986871, 4.989161, 4.991158, 4.992808, 4.994019, 4.994727, 
    4.994781, 4.994075, 4.992127, 4.990852, 4.98828, 4.984199, 4.978396, 
    4.970678, 4.960901, 4.949014, 4.935112, 4.919465, 4.902544, 4.885012, 
    4.867685, 4.851458, 4.837206, 4.825689, 4.817468, 4.812854, 4.811893, 
    4.814398,
  // momentumY(22,8, 0-49)
    4.88981, 4.895993, 4.902441, 4.908971, 4.915441, 4.921747, 4.927812, 
    4.933593, 4.939067, 4.944226, 4.949075, 4.953628, 4.957908, 4.96194, 
    4.965762, 4.967212, 4.971738, 4.974128, 4.976008, 4.977619, 4.979063, 
    4.982004, 4.98441, 4.986624, 4.988671, 4.990512, 4.992086, 4.993325, 
    4.994076, 4.994135, 4.992996, 4.992678, 4.991173, 4.988257, 4.983695, 
    4.977253, 4.968738, 4.958027, 4.945134, 4.930234, 4.913712, 4.896164, 
    4.878372, 4.86124, 4.845705, 4.832624, 4.822687, 4.816338, 4.813755, 
    4.814858,
  // momentumY(22,9, 0-49)
    4.892284, 4.898389, 4.904727, 4.911123, 4.917439, 4.923574, 4.929457, 
    4.935043, 4.94031, 4.945249, 4.949864, 4.954177, 4.958208, 4.96199, 
    4.965567, 4.966765, 4.970487, 4.972616, 4.974267, 4.975658, 4.976905, 
    4.979655, 4.981893, 4.983966, 4.986002, 4.987977, 4.989863, 4.991588, 
    4.993001, 4.993782, 4.993412, 4.993945, 4.993408, 4.991569, 4.988178, 
    4.982973, 4.975715, 4.966225, 4.954433, 4.940427, 4.924498, 4.90716, 
    4.889142, 4.871335, 4.854712, 4.84022, 4.828661, 4.820616, 4.8164, 
    4.816047,
  // momentumY(22,10, 0-49)
    4.895145, 4.901142, 4.907338, 4.913567, 4.919698, 4.925632, 4.931304, 
    4.93667, 4.941706, 4.946405, 4.950773, 4.95483, 4.958596, 4.96211, 
    4.965409, 4.96648, 4.969285, 4.971148, 4.972591, 4.973794, 4.974871, 
    4.977384, 4.979412, 4.981291, 4.983261, 4.985313, 4.987463, 4.989625, 
    4.991659, 4.993119, 4.993484, 4.99475, 4.995069, 4.994203, 4.991892, 
    4.987855, 4.981818, 4.973549, 4.96291, 4.949902, 4.93472, 4.917789, 
    4.899768, 4.881516, 4.864025, 4.8483, 4.835255, 4.825601, 4.819786, 
    4.817967,
  // momentumY(22,11, 0-49)
    4.898359, 4.904222, 4.910252, 4.916286, 4.922204, 4.927913, 4.93335, 
    4.938472, 4.943258, 4.947702, 4.951809, 4.955594, 4.959082, 4.962301, 
    4.965283, 4.966367, 4.968176, 4.969769, 4.971031, 4.972083, 4.973031, 
    4.975266, 4.977045, 4.978685, 4.980544, 4.98263, 4.984991, 4.987542, 
    4.990149, 4.992247, 4.993314, 4.995196, 4.996253, 4.996246, 4.994911, 
    4.991952, 4.987071, 4.979993, 4.970516, 4.958566, 4.944244, 4.927882, 
    4.910058, 4.891582, 4.873441, 4.856687, 4.842321, 4.831179, 4.823837, 
    4.82058,
  // momentumY(22,12, 0-49)
    4.901878, 4.907592, 4.913434, 4.919252, 4.924936, 4.930398, 4.935579, 
    4.940441, 4.944962, 4.949134, 4.952963, 4.956466, 4.959656, 4.962557, 
    4.965181, 4.966418, 4.967177, 4.968506, 4.96962, 4.970567, 4.97143, 
    4.973352, 4.974858, 4.976231, 4.977943, 4.980022, 4.98255, 4.985436, 
    4.988568, 4.991255, 4.992997, 4.995377, 4.997054, 4.99779, 4.997318, 
    4.995336, 4.991525, 4.98558, 4.977245, 4.966374, 4.952986, 4.937315, 
    4.919857, 4.901359, 4.882782, 4.865209, 4.849709, 4.837227, 4.828466, 
    4.823829,
  // momentumY(22,13, 0-49)
    4.90565, 4.911202, 4.916841, 4.922431, 4.927863, 4.933063, 4.937972, 
    4.942556, 4.946795, 4.950685, 4.954226, 4.957429, 4.960305, 4.962861, 
    4.96509, 4.966601, 4.96628, 4.967366, 4.968375, 4.969272, 4.970106, 
    4.971691, 4.97291, 4.973999, 4.975545, 4.977583, 4.980232, 4.9834, 
    4.986999, 4.990225, 4.992621, 4.995386, 4.997564, 4.998925, 4.999202, 
    4.998087, 4.99525, 4.990359, 4.983118, 4.973319, 4.960899, 4.946009, 
    4.92905, 4.910706, 4.891897, 4.873711, 4.857275, 4.843622, 4.83357, 
    4.827637,
  // momentumY(22,14, 0-49)
    4.909611, 4.915001, 4.920432, 4.925782, 4.930954, 4.935875, 4.940499, 
    4.944792, 4.948737, 4.952328, 4.955569, 4.958461, 4.961009, 4.963201, 
    4.965012, 4.966866, 4.965448, 4.966335, 4.967295, 4.968207, 4.969079, 
    4.970313, 4.971245, 4.97205, 4.973421, 4.975398, 4.978127, 4.981521, 
    4.985519, 4.989235, 4.992261, 4.995299, 4.997867, 4.999737, 5.000646, 
    5.000288, 4.998318, 4.994392, 4.988178, 4.979414, 4.96797, 4.953912, 
    4.937561, 4.919518, 4.900659, 4.882061, 4.864886, 4.850241, 4.839045, 
    4.831921,
  // momentumY(22,15, 0-49)
    4.913706, 4.918937, 4.924161, 4.929266, 4.934164, 4.938797, 4.943122, 
    4.947111, 4.950749, 4.954034, 4.956963, 4.959537, 4.961747, 4.96357, 
    4.964959, 4.967154, 4.964622, 4.965373, 4.966358, 4.967362, 4.968349, 
    4.96923, 4.969894, 4.970437, 4.971638, 4.973541, 4.976313, 4.979875, 
    4.984203, 4.988347, 4.99198, 4.995186, 4.998031, 5.000298, 5.001725, 
    5.002008, 5.000802, 4.997742, 4.992472, 4.984691, 4.974206, 4.96101, 
    4.945339, 4.927721, 4.908974, 4.89015, 4.87243, 4.856977, 4.844789, 
    4.836594,
  // momentumY(22,16, 0-49)
    4.917878, 4.922956, 4.927972, 4.932827, 4.937447, 4.94178, 4.945793, 
    4.949466, 4.952789, 4.95576, 4.958376, 4.960632, 4.962512, 4.963979, 
    4.964971, 4.967404, 4.963717, 4.964427, 4.965526, 4.966713, 4.967906, 
    4.968447, 4.96888, 4.969199, 4.970256, 4.972084, 4.974867, 4.978536, 
    4.983116, 4.987617, 4.991826, 4.995096, 4.998113, 5.000667, 5.002501, 
    5.003314, 5.00276, 5.000465, 4.996054, 4.989187, 4.979626, 4.967295, 
    4.952357, 4.935261, 4.916767, 4.897888, 4.879806, 4.863722, 4.850706, 
    4.841565,
  // momentumY(22,17, 0-49)
    4.92207, 4.926999, 4.931807, 4.936404, 4.940733, 4.944755, 4.948444, 
    4.951794, 4.9548, 4.957461, 4.959776, 4.961733, 4.963308, 4.964456, 
    4.965109, 4.967572, 4.962652, 4.963425, 4.964743, 4.966219, 4.967717, 
    4.967952, 4.96821, 4.968366, 4.96932, 4.971087, 4.973859, 4.977577, 
    4.982324, 4.9871, 4.991838, 4.99507, 4.998154, 5.000888, 5.00302, 
    5.004251, 5.00424, 5.002608, 4.998962, 4.992938, 4.984252, 4.972774, 
    4.9586, 4.942105, 4.923982, 4.905201, 4.886931, 4.870391, 4.856705, 
    4.846749,
  // momentumY(22,18, 0-49)
    4.926219, 4.930993, 4.935577, 4.939902, 4.943923, 4.94762, 4.950982, 
    4.954012, 4.956714, 4.95909, 4.961139, 4.96284, 4.964164, 4.96506, 
    4.965462, 4.967654, 4.961352, 4.962304, 4.963949, 4.965824, 4.967738, 
    4.967719, 4.967881, 4.967954, 4.96887, 4.970606, 4.973351, 4.977064, 
    4.981887, 4.986845, 4.99204, 4.995138, 4.998181, 5.000986, 5.003305, 
    5.004848, 5.005273, 5.004199, 5.001225, 4.995965, 4.988102, 4.977455, 
    4.964059, 4.948224, 4.930574, 4.912029, 4.893728, 4.876899, 4.862697, 
    4.852058,
  // momentumY(22,19, 0-49)
    4.930254, 4.934838, 4.939164, 4.943184, 4.946876, 4.950236, 4.953277, 
    4.95601, 4.958449, 4.960598, 4.962448, 4.963972, 4.965132, 4.96587, 
    4.966131, 4.967701, 4.959782, 4.961017, 4.963089, 4.965472, 4.967917, 
    4.967721, 4.967884, 4.967977, 4.968936, 4.970692, 4.973415, 4.977076, 
    4.981885, 4.986914, 4.992465, 4.995318, 4.998209, 5.000971, 5.003365, 
    5.005108, 5.005862, 5.005246, 5.002851, 4.998276, 4.991178, 4.981333, 
    4.968722, 4.953592, 4.936501, 4.918311, 4.900126, 4.883163, 4.868595, 
    4.857404,
  // momentumY(22,20, 0-49)
    4.935121, 4.940522, 4.945562, 4.95019, 4.954374, 4.958099, 4.961357, 
    4.964148, 4.966482, 4.968373, 4.969851, 4.970959, 4.971753, 4.972302, 
    4.972693, 0, 4.959976, 4.961293, 4.963098, 4.965001, 4.966878, 4.965349, 
    4.964415, 4.963618, 4.964009, 4.965533, 4.968349, 4.972388, 4.97783, 
    4.983681, 4.990357, 4.993667, 4.997002, 5.000195, 5.003012, 5.00518, 
    5.006382, 5.006256, 5.004407, 5.000442, 4.994011, 4.984875, 4.972975, 
    4.958509, 4.941978, 4.924188, 4.906198, 4.8892, 4.874375, 4.862727,
  // momentumY(22,21, 0-49)
    4.939007, 4.944368, 4.949268, 4.953667, 4.957558, 4.960947, 4.963851, 
    4.966298, 4.968316, 4.969938, 4.971203, 4.972163, 4.972878, 4.973427, 
    4.973916, 0, 4.955731, 4.957488, 4.959795, 4.962227, 4.964609, 4.962763, 
    4.96166, 4.960739, 4.961128, 4.962759, 4.965786, 4.970114, 4.975934, 
    4.982237, 4.989596, 4.992975, 4.996485, 4.999949, 5.003128, 5.00574, 
    5.007459, 5.007914, 5.006705, 5.003426, 4.997713, 4.989299, 4.978093, 
    4.964244, 4.948203, 4.930723, 4.912822, 4.895671, 4.880454, 4.868197,
  // momentumY(22,22, 0-49)
    4.942727, 4.948107, 4.952914, 4.957129, 4.960762, 4.96384, 4.966405, 
    4.968505, 4.970191, 4.971513, 4.972527, 4.973292, 4.973882, 4.974389, 
    4.974936, 0, 4.952352, 4.954473, 4.957218, 4.960129, 4.962974, 4.960836, 
    4.959574, 4.958531, 4.958904, 4.960607, 4.963778, 4.968307, 4.974384, 
    4.980988, 4.988835, 4.992147, 4.995678, 4.999262, 5.002652, 5.005566, 
    5.007674, 5.008605, 5.007951, 5.005296, 5.000262, 4.99256, 4.982064, 
    4.968881, 4.953407, 4.936348, 4.918674, 4.901524, 4.886073, 4.873363,
  // momentumY(22,23, 0-49)
    4.946211, 4.951646, 4.956401, 4.960465, 4.963868, 4.966659, 4.968901, 
    4.970664, 4.972017, 4.973031, 4.973774, 4.974321, 4.974754, 4.975182, 
    4.975747, 0, 4.949856, 4.952229, 4.955276, 4.958517, 4.961682, 4.959258, 
    4.957822, 4.956636, 4.956953, 4.958671, 4.961921, 4.966574, 4.97282, 
    4.979625, 4.98781, 4.991016, 4.994521, 4.998165, 5.001703, 5.004858, 
    5.007296, 5.008648, 5.0085, 5.006428, 5.002038, 4.995022, 4.98522, 
    4.972703, 4.957818, 4.94122, 4.923836, 4.906774, 4.891189, 4.878129,
  // momentumY(22,24, 0-49)
    4.949394, 4.954908, 4.959633, 4.963575, 4.966775, 4.969305, 4.971246, 
    4.972689, 4.973722, 4.97443, 4.9749, 4.975216, 4.975473, 4.975791, 
    4.976331, 0, 4.948518, 4.951012, 4.954212, 4.957628, 4.960968, 4.958356, 
    4.95681, 4.955535, 4.955814, 4.957535, 4.960822, 4.965538, 4.971878, 
    4.978793, 4.987182, 4.990316, 4.993803, 4.997482, 5.001118, 5.004433, 
    5.007102, 5.008749, 5.008963, 5.007317, 5.003409, 4.996915, 4.987658, 
    4.975676, 4.961286, 4.945103, 4.928017, 4.911108, 4.895511, 4.882263,
  // momentumY(22,25, 0-49)
    4.952204, 4.957809, 4.962523, 4.966364, 4.969392, 4.971691, 4.973362, 
    4.97451, 4.975244, 4.975662, 4.975863, 4.975944, 4.97601, 4.976191, 
    4.976657, 0, 4.948055, 4.950538, 4.953739, 4.957167, 4.960527, 4.957858, 
    4.956294, 4.955017, 4.955307, 4.957049, 4.960361, 4.965107, 4.971481, 
    4.978438, 4.986895, 4.990032, 4.993546, 4.99728, 5.001002, 5.004436, 
    5.00726, 5.0091, 5.009548, 5.008173, 5.004572, 4.998418, 4.989519, 
    4.977905, 4.96387, 4.948008, 4.931185, 4.914455, 4.898934, 4.885649,
  // momentumY(22,26, 0-49)
    4.95458, 4.960278, 4.964995, 4.96876, 4.971643, 4.973747, 4.975185, 
    4.976077, 4.97654, 4.97669, 4.976631, 4.976472, 4.976333, 4.976344, 
    4.976682, 0, 4.948453, 4.950796, 4.953845, 4.957116, 4.960338, 4.957754, 
    4.956271, 4.955087, 4.95545, 4.95724, 4.960577, 4.965328, 4.97169, 
    4.978623, 4.98702, 4.990255, 4.993862, 4.997688, 5.001496, 5.005016, 
    5.007926, 5.009855, 5.010394, 5.00912, 5.00563, 4.999599, 4.990843, 
    4.979391, 4.965537, 4.949868, 4.933245, 4.916705, 4.901348, 4.888179,
  // momentumY(22,27, 0-49)
    4.95647, 4.962255, 4.966988, 4.970704, 4.973483, 4.975435, 4.976684, 
    4.977357, 4.977584, 4.977483, 4.977173, 4.976769, 4.976398, 4.976196, 
    4.976342, 0, 4.94983, 4.951895, 4.954633, 4.957582, 4.960505, 4.958111, 
    4.956778, 4.955749, 4.956214, 4.95806, 4.961405, 4.966125, 4.972418, 
    4.979264, 4.98748, 4.990894, 4.994651, 4.998594, 5.002487, 5.006057, 
    5.008984, 5.010896, 5.011392, 5.010053, 5.006485, 5.000376, 4.991556, 
    4.98007, 4.96623, 4.950636, 4.934154, 4.917815, 4.902705, 4.889807,
  // momentumY(22,28, 0-49)
    4.957836, 4.963705, 4.968472, 4.972172, 4.974893, 4.976745, 4.977857, 
    4.978356, 4.978376, 4.978041, 4.977476, 4.976804, 4.976159, 4.975689, 
    4.975567, 0, 4.952566, 4.954219, 4.956491, 4.958948, 4.961411, 4.95925, 
    4.958077, 4.957208, 4.95776, 4.959622, 4.962923, 4.967553, 4.973707, 
    4.980392, 4.988312, 4.991958, 4.995893, 4.999952, 5.003895, 5.00745, 
    5.010296, 5.012068, 5.012367, 5.010787, 5.006949, 5.000559, 4.991478, 
    4.979781, 4.965812, 4.950198, 4.933821, 4.917719, 4.90296, 4.890495,
  // momentumY(22,29, 0-49)
    4.95867, 4.964626, 4.969453, 4.973186, 4.975905, 4.977718, 4.978745, 
    4.979113, 4.978947, 4.978374, 4.97753, 4.976545, 4.975567, 4.974751, 
    4.974271, 0, 4.95646, 4.95757, 4.959221, 4.961021, 4.962852, 4.960859, 
    4.959756, 4.958962, 4.95951, 4.961305, 4.96448, 4.968947, 4.974889, 
    4.981332, 4.988841, 4.992712, 4.996807, 5.000953, 5.004909, 5.008403, 
    5.011117, 5.012687, 5.012722, 5.010827, 5.006638, 4.999887, 4.990465, 
    4.978487, 4.964337, 4.94868, 4.932421, 4.916602, 4.902275, 4.890357,
  // momentumY(22,30, 0-49)
    4.958047, 4.963116, 4.967086, 4.970015, 4.972012, 4.973216, 4.973781, 
    4.973852, 4.973566, 4.973029, 4.972315, 4.97146, 4.970461, 4.969284, 
    4.96787, 4.971422, 4.957416, 4.958146, 4.959991, 4.962359, 4.964968, 
    4.964603, 4.964927, 4.965328, 4.966667, 4.968801, 4.971864, 4.975824, 
    4.980929, 4.98633, 4.992523, 4.995769, 4.999239, 5.002778, 5.006158, 
    5.009108, 5.011305, 5.01238, 5.011932, 5.009561, 5.00491, 4.997726, 
    4.987928, 4.975666, 4.961368, 4.945735, 4.929695, 4.914293, 4.900559, 
    4.889373,
  // momentumY(22,31, 0-49)
    4.95789, 4.963067, 4.967144, 4.970172, 4.972244, 4.973488, 4.974046, 
    4.974065, 4.973676, 4.972998, 4.972118, 4.97109, 4.969933, 4.968622, 
    4.967101, 4.971066, 4.959039, 4.959276, 4.960526, 4.96225, 4.964221, 
    4.963971, 4.964255, 4.964615, 4.965906, 4.968037, 4.971161, 4.975234, 
    4.980437, 4.98588, 4.991862, 4.995546, 4.999402, 5.003253, 5.00686, 
    5.009934, 5.012142, 5.013105, 5.012422, 5.009698, 5.004597, 4.9969, 
    4.986571, 4.973823, 4.959142, 4.94329, 4.927226, 4.912013, 4.898664, 
    4.888015,
  // momentumY(22,32, 0-49)
    4.957166, 4.962335, 4.966437, 4.969514, 4.971652, 4.972965, 4.973582, 
    4.97364, 4.973271, 4.972588, 4.971687, 4.970632, 4.969455, 4.968151, 
    4.96666, 4.970359, 4.96031, 4.960156, 4.960892, 4.962051, 4.963462, 
    4.963401, 4.963728, 4.964138, 4.96545, 4.967617, 4.970803, 4.974948, 
    4.980169, 4.985564, 4.991252, 4.995315, 4.999488, 5.003579, 5.007331, 
    5.010444, 5.012566, 5.013313, 5.012284, 5.009094, 5.003433, 4.995127, 
    4.984194, 4.970913, 4.955841, 4.939794, 4.923772, 4.908843, 4.895998, 
    4.886026,
  // momentumY(22,33, 0-49)
    4.955983, 4.961055, 4.965122, 4.968218, 4.970413, 4.971811, 4.972531, 
    4.972694, 4.972424, 4.971832, 4.971011, 4.970033, 4.968942, 4.967745, 
    4.966402, 4.969375, 4.961257, 4.960827, 4.96114, 4.961818, 4.962752, 
    4.962927, 4.963367, 4.963902, 4.965289, 4.967519, 4.970751, 4.974916, 
    4.980073, 4.985337, 4.990673, 4.995048, 4.999469, 5.003721, 5.007534, 
    5.010592, 5.01253, 5.012957, 5.011473, 5.007711, 5.001394, 4.992397, 
    4.980807, 4.966975, 4.951529, 4.935343, 4.919448, 4.904913, 4.892695, 
    4.883534,
  // momentumY(22,34, 0-49)
    4.954448, 4.95936, 4.963346, 4.966434, 4.968682, 4.970178, 4.971027, 
    4.971339, 4.971222, 4.970782, 4.970108, 4.969277, 4.968343, 4.967324, 
    4.966204, 4.968204, 4.961935, 4.961338, 4.961315, 4.96159, 4.962114, 
    4.962554, 4.963157, 4.963874, 4.965377, 4.967681, 4.970933, 4.975061, 
    4.980067, 4.985126, 4.99007, 4.994689, 4.999281, 5.003613, 5.007399, 
    5.010306, 5.01196, 5.011963, 5.009924, 5.005498, 4.998452, 4.988713, 
    4.976445, 4.962076, 4.946308, 4.930067, 4.914408, 4.900389, 4.888928, 
    4.880701,
  // momentumY(22,35, 0-49)
    4.952672, 4.957375, 4.961246, 4.964301, 4.966592, 4.968191, 4.969186, 
    4.969673, 4.969746, 4.969497, 4.969015, 4.968374, 4.967635, 4.966836, 
    4.965979, 4.966949, 4.962429, 4.961751, 4.961463, 4.961401, 4.961579, 
    4.962293, 4.96309, 4.964033, 4.965674, 4.968048, 4.971286, 4.975313, 
    4.980082, 4.984866, 4.989388, 4.994173, 4.99885, 5.00317, 5.006832, 
    5.00949, 5.010759, 5.010242, 5.00756, 5.002398, 4.994569, 4.984073, 
    4.971148, 4.9563, 4.940302, 4.924123, 4.908833, 4.895466, 4.88489, 
    4.877709,
  // momentumY(22,36, 0-49)
    4.950771, 4.955221, 4.958945, 4.961947, 4.96427, 4.965969, 4.967115, 
    4.96779, 4.968071, 4.968041, 4.967778, 4.967352, 4.96683, 4.966259, 
    4.965673, 4.965696, 4.962821, 4.962123, 4.961627, 4.961285, 4.961173, 
    4.96215, 4.963158, 4.96435, 4.96614, 4.968571, 4.97175, 4.975606, 
    4.980051, 4.984489, 4.988561, 4.993416, 4.99808, 5.002285, 5.005719, 
    5.008024, 5.008811, 5.007683, 5.004285, 4.998341, 4.98972, 4.978488, 
    4.96497, 4.949749, 4.933655, 4.917694, 4.902929, 4.890361, 4.880794, 
    4.874759,
  // momentumY(22,37, 0-49)
    4.948856, 4.953017, 4.956562, 4.959488, 4.961827, 4.963615, 4.964911, 
    4.965777, 4.966276, 4.966475, 4.966443, 4.966245, 4.965945, 4.9656, 
    4.965266, 4.964514, 4.963181, 4.962499, 4.961835, 4.961262, 4.960908, 
    4.962128, 4.963348, 4.964801, 4.966734, 4.969196, 4.972267, 4.975879, 
    4.979912, 4.983932, 4.987516, 4.992332, 4.996866, 5.000842, 5.003934, 
    5.005777, 5.005983, 5.004169, 5.000006, 4.993264, 4.983874, 4.971982, 
    4.957987, 4.942545, 4.926535, 4.910977, 4.896918, 4.885301, 4.876864, 
    4.872054,
  // momentumY(22,38, 0-49)
    4.947029, 4.95087, 4.954208, 4.957035, 4.959365, 4.961228, 4.962661, 
    4.96371, 4.964424, 4.964855, 4.965057, 4.965089, 4.965008, 4.964876, 
    4.964758, 4.963451, 4.963553, 4.962902, 4.962105, 4.961343, 4.960793, 
    4.962229, 4.963652, 4.965358, 4.967416, 4.969876, 4.972776, 4.976065, 
    4.979594, 4.983118, 4.98617, 4.990817, 4.995093, 4.99871, 5.00134, 
    5.002613, 5.00215, 4.999588, 4.994634, 4.987115, 4.977029, 4.964597, 
    4.950294, 4.934833, 4.919126, 4.904189, 4.891028, 4.880522, 4.873323, 
    4.869796,
  // momentumY(22,39, 0-49)
    4.945388, 4.948878, 4.95198, 4.954679, 4.956977, 4.958889, 4.960439, 
    4.961655, 4.962572, 4.963227, 4.96366, 4.963917, 4.964046, 4.964107, 
    4.964168, 4.96253, 4.963966, 4.963343, 4.962438, 4.96153, 4.960828, 
    4.962446, 4.964049, 4.965991, 4.968144, 4.970555, 4.973221, 4.976102, 
    4.979031, 4.981975, 4.984433, 4.988768, 4.992643, 4.995764, 4.997804, 
    4.9984, 4.997189, 4.993839, 4.988104, 4.979869, 4.969203, 4.956405, 
    4.94201, 4.926777, 4.911627, 4.89755, 4.885493, 4.876248, 4.870383, 
    4.868177,
  // momentumY(22,40, 0-49)
    4.944005, 4.947119, 4.949958, 4.952499, 4.954735, 4.956668, 4.958309, 
    4.959668, 4.960769, 4.96163, 4.962281, 4.962752, 4.96308, 4.963314, 
    4.963518, 4.961757, 4.964414, 4.963816, 4.962826, 4.961812, 4.960998, 
    4.962762, 4.964519, 4.966666, 4.968871, 4.971179, 4.973535, 4.975921, 
    4.978155, 4.980425, 4.982213, 4.986079, 4.989399, 4.99188, 4.993204, 
    4.993023, 4.991001, 4.986851, 4.980374, 4.971526, 4.960449, 4.947505, 
    4.933281, 4.918559, 4.904246, 4.891278, 4.880527, 4.87269, 4.868237, 
    4.867364,
  // momentumY(22,41, 0-49)
    4.942934, 4.945651, 4.948199, 4.950552, 4.952695, 4.954617, 4.956311, 
    4.957786, 4.959041, 4.960086, 4.960935, 4.961604, 4.962116, 4.962505, 
    4.962822, 4.961109, 4.964873, 4.964289, 4.963243, 4.96216, 4.961271, 
    4.963148, 4.965024, 4.967335, 4.969543, 4.971682, 4.973652, 4.975451, 
    4.976894, 4.978395, 4.979421, 4.98265, 4.985257, 4.986954, 4.987439, 
    4.986394, 4.983522, 4.978585, 4.971448, 4.962138, 4.950858, 4.938031, 
    4.924275, 4.910371, 4.897185, 4.885581, 4.876331, 4.870027, 4.86704, 
    4.867486,
  // momentumY(22,42, 0-49)
    4.942198, 4.944501, 4.946737, 4.948874, 4.950887, 4.952759, 4.954475, 
    4.956024, 4.957401, 4.9586, 4.959621, 4.960468, 4.961146, 4.961676, 
    4.962083, 4.960546, 4.965296, 4.964724, 4.963648, 4.962533, 4.961604, 
    4.963559, 4.96552, 4.967943, 4.970094, 4.971998, 4.973501, 4.974625, 
    4.975183, 4.975811, 4.975973, 4.978401, 4.980134, 4.980906, 4.980445, 
    4.978471, 4.974735, 4.969062, 4.961384, 4.951796, 4.940564, 4.928149, 
    4.91518, 4.90241, 4.890639, 4.880638, 4.873065, 4.868399, 4.866908, 
    4.868633,
  // momentumY(22,43, 0-49)
    4.941798, 4.943673, 4.945574, 4.947466, 4.949317, 4.951102, 4.952796, 
    4.954382, 4.95584, 4.957156, 4.958319, 4.959318, 4.960145, 4.9608, 
    4.961287, 4.960012, 4.965619, 4.965061, 4.963984, 4.962872, 4.961929, 
    4.963934, 4.965942, 4.968421, 4.970454, 4.972047, 4.973005, 4.973367, 
    4.972955, 4.97261, 4.971803, 4.973268, 4.973981, 4.973707, 4.972209, 
    4.969264, 4.964683, 4.958358, 4.950296, 4.940651, 4.929743, 4.918052, 
    4.906193, 4.894865, 4.884781, 4.876598, 4.870849, 4.867894, 4.867904, 
    4.870842,
  // momentumY(22,44, 0-49)
    4.941687, 4.943127, 4.944678, 4.9463, 4.947957, 4.949617, 4.95125, 
    4.952827, 4.954327, 4.955722, 4.956991, 4.958113, 4.959068, 4.959835, 
    4.960393, 4.959428, 4.965758, 4.965227, 4.96418, 4.963101, 4.962169, 
    4.964197, 4.966213, 4.968689, 4.970536, 4.971749, 4.972087, 4.97161, 
    4.970154, 4.968743, 4.966866, 4.967227, 4.966793, 4.965372, 4.962781, 
    4.958857, 4.953483, 4.946626, 4.938364, 4.928908, 4.918612, 4.907955, 
    4.897513, 4.88791, 4.87975, 4.87356, 4.869744, 4.868541, 4.870022, 
    4.874084,
  // momentumY(22,45, 0-49)
    4.941793, 4.942795, 4.943985, 4.945317, 4.946753, 4.948253, 4.949785, 
    4.951314, 4.952811, 4.954244, 4.955584, 4.9568, 4.957859, 4.958724, 
    4.959352, 4.958708, 4.965632, 4.96514, 4.964149, 4.963128, 4.962224, 
    4.964252, 4.966239, 4.96865, 4.97025, 4.971015, 4.97067, 4.969294, 
    4.966736, 4.964185, 4.961152, 4.960292, 4.958618, 4.955986, 4.952279, 
    4.947404, 4.941326, 4.934086, 4.92583, 4.916817, 4.907412, 4.898078, 
    4.889328, 4.881688, 4.875639, 4.87157, 4.869749, 4.870298, 4.873192, 
    4.878266,
  // momentumY(22,46, 0-49)
    4.942007, 4.942574, 4.943394, 4.944422, 4.945613, 4.946927, 4.948323, 
    4.949766, 4.951222, 4.952654, 4.954029, 4.955307, 4.956448, 4.957397, 
    4.958094, 4.957758, 4.965144, 4.964711, 4.963798, 4.962851, 4.961987, 
    4.963995, 4.965917, 4.968205, 4.969499, 4.96976, 4.968681, 4.966363, 
    4.962676, 4.958935, 4.954689, 4.952533, 4.949564, 4.9457, 4.940897, 
    4.935141, 4.928477, 4.921025, 4.91299, 4.904661, 4.896404, 4.888639, 
    4.881803, 4.876304, 4.87249, 4.870608, 4.870795, 4.873055, 4.877275, 
    4.88323,
  // momentumY(22,47, 0-49)
    4.942184, 4.942324, 4.942777, 4.943493, 4.944427, 4.94553, 4.946764, 
    4.948091, 4.949472, 4.950871, 4.952249, 4.95356, 4.954759, 4.955781, 
    4.956546, 4.956481, 4.964205, 4.963849, 4.963029, 4.962167, 4.961345, 
    4.963313, 4.965137, 4.967248, 4.968189, 4.967905, 4.966066, 4.96279, 
    4.957972, 4.953028, 4.947546, 4.944068, 4.939801, 4.934735, 4.928899, 
    4.922368, 4.915265, 4.907782, 4.900171, 4.892743, 4.885846, 4.879838, 
    4.875064, 4.87181, 4.870286, 4.870596, 4.872749, 4.876638, 4.882066, 
    4.888757,
  // momentumY(22,48, 0-49)
    4.942157, 4.941879, 4.941971, 4.942379, 4.943048, 4.943933, 4.94499, 
    4.94618, 4.947465, 4.948805, 4.95016, 4.951481, 4.952719, 4.953801, 
    4.954633, 4.95479, 4.962732, 4.962471, 4.961751, 4.960971, 4.960187, 
    4.962099, 4.963796, 4.965682, 4.966233, 4.965381, 4.962782, 4.958564, 
    4.952653, 4.946531, 4.939835, 4.935065, 4.929556, 4.923367, 4.916611, 
    4.909441, 4.902061, 4.894722, 4.887719, 4.881363, 4.875974, 4.871838, 
    4.869196, 4.86821, 4.868954, 4.871396, 4.875418, 4.880815, 4.887309, 
    4.894578,
  // momentumY(22,49, 0-49)
    4.942302, 4.941273, 4.940712, 4.94055, 4.940726, 4.94118, 4.941866, 
    4.942734, 4.943739, 4.944835, 4.945973, 4.947086, 4.948108, 4.94893, 
    4.949424, 4.949001, 4.964243, 4.962885, 4.960816, 4.958843, 4.957083, 
    4.960893, 4.964464, 4.968607, 4.970275, 4.969415, 4.9654, 4.958524, 
    4.948629, 4.938767, 4.928291, 4.922237, 4.915466, 4.908151, 4.900531, 
    4.892879, 4.885505, 4.878732, 4.872895, 4.868293, 4.865188, 4.863756, 
    4.864096, 4.866197, 4.869948, 4.875145, 4.881518, 4.888731, 4.896425, 
    4.904231,
  // momentumY(23,0, 0-49)
    4.895426, 4.901486, 4.90759, 4.913628, 4.919533, 4.92527, 4.930825, 
    4.936199, 4.941404, 4.946454, 4.951359, 4.956124, 4.960742, 4.965197, 
    4.969453, 4.973246, 4.977482, 4.980842, 4.983828, 4.986425, 4.988595, 
    4.990544, 4.991959, 4.992893, 4.993297, 4.993151, 4.992422, 4.991085, 
    4.989092, 4.986431, 4.982956, 4.978846, 4.973688, 4.967337, 4.959653, 
    4.950525, 4.939891, 4.927777, 4.914315, 4.899775, 4.884562, 4.869212, 
    4.85435, 4.840641, 4.828725, 4.819151, 4.812321, 4.808452, 4.807563, 
    4.809484,
  // momentumY(23,1, 0-49)
    4.896116, 4.90232, 4.908538, 4.914664, 4.920634, 4.92641, 4.931978, 
    4.937342, 4.942514, 4.947505, 4.952327, 4.956984, 4.961471, 4.965774, 
    4.969862, 4.97324, 4.977746, 4.980855, 4.983581, 4.985966, 4.987989, 
    4.990112, 4.991745, 4.993001, 4.993792, 4.994096, 4.993859, 4.993059, 
    4.991638, 4.989619, 4.986797, 4.983615, 4.979371, 4.973888, 4.966999, 
    4.958545, 4.948429, 4.936629, 4.923249, 4.908527, 4.892865, 4.876808, 
    4.861016, 4.846209, 4.8331, 4.822316, 4.814339, 4.809461, 4.807758, 
    4.809104,
  // momentumY(23,2, 0-49)
    4.896848, 4.903163, 4.909467, 4.915654, 4.921661, 4.927448, 4.933006, 
    4.938334, 4.943444, 4.948349, 4.953061, 4.957585, 4.961919, 4.966052, 
    4.96996, 4.972911, 4.977615, 4.980476, 4.982946, 4.985118, 4.986993, 
    4.989272, 4.991097, 4.992633, 4.993772, 4.994483, 4.9947, 4.994403, 
    4.993524, 4.99211, 4.989905, 4.987619, 4.98428, 4.979692, 4.973659, 
    4.965992, 4.956553, 4.945277, 4.932223, 4.917595, 4.901763, 4.885261, 
    4.868759, 4.853016, 4.838797, 4.826807, 4.81761, 4.81158, 4.808866, 
    4.809398,
  // momentumY(23,3, 0-49)
    4.897707, 4.904102, 4.910461, 4.91668, 4.922695, 4.928468, 4.933987, 
    4.939251, 4.944274, 4.949068, 4.953646, 4.958017, 4.962181, 4.966132, 
    4.969855, 4.972373, 4.977182, 4.979805, 4.98203, 4.983992, 4.985715, 
    4.988125, 4.990106, 4.991872, 4.993307, 4.994374, 4.994997, 4.99516, 
    4.994784, 4.993926, 4.992285, 4.990835, 4.988363, 4.984661, 4.979513, 
    4.972706, 4.964067, 4.953493, 4.940991, 4.926718, 4.910996, 4.894328, 
    4.877372, 4.860893, 4.845701, 4.832562, 4.822122, 4.814842, 4.810956, 
    4.810467,
  // momentumY(23,4, 0-49)
    4.898767, 4.905207, 4.911588, 4.917809, 4.923801, 4.929531, 4.934984, 
    4.940162, 4.945074, 4.949735, 4.954161, 4.958361, 4.962342, 4.966105, 
    4.969644, 4.971735, 4.976532, 4.978934, 4.980926, 4.982686, 4.984258, 
    4.986763, 4.988861, 4.990802, 4.992469, 4.993831, 4.994809, 4.995383, 
    4.99547, 4.995112, 4.993973, 4.993282, 4.991616, 4.988761, 4.984494, 
    4.978585, 4.970834, 4.9611, 4.949344, 4.935659, 4.920317, 4.903763, 
    4.886617, 4.869635, 4.853644, 4.839461, 4.827805, 4.819223, 4.814049, 
    4.812364,
  // momentumY(23,5, 0-49)
    4.900073, 4.906525, 4.912896, 4.919085, 4.925028, 4.930689, 4.93605, 
    4.941118, 4.945899, 4.950413, 4.95467, 4.958691, 4.962481, 4.966052, 
    4.969409, 4.971094, 4.975749, 4.977942, 4.979719, 4.981287, 4.982709, 
    4.985273, 4.987438, 4.989486, 4.991323, 4.992917, 4.994195, 4.995135, 
    4.995642, 4.995732, 4.995035, 4.995014, 4.994076, 4.992012, 4.988597, 
    4.983593, 4.976781, 4.967987, 4.957124, 4.94423, 4.929503, 4.913324, 
    4.896254, 4.879013, 4.862425, 4.847337, 4.834532, 4.824646, 4.818106, 
    4.815096,
  // momentumY(23,6, 0-49)
    4.901654, 4.908082, 4.914409, 4.920537, 4.926403, 4.931969, 4.937221, 
    4.94216, 4.946796, 4.951147, 4.95523, 4.959061, 4.962658, 4.966038, 
    4.969217, 4.970532, 4.974907, 4.976904, 4.978485, 4.979873, 4.981148, 
    4.983724, 4.985905, 4.987993, 4.989932, 4.991693, 4.993219, 4.994479, 
    4.995372, 4.995861, 4.995553, 4.996108, 4.995815, 4.994474, 4.991864, 
    4.987747, 4.98189, 4.974093, 4.964232, 4.952282, 4.938368, 4.922791, 
    4.906042, 4.888782, 4.87181, 4.855984, 4.842136, 4.830983, 4.823049, 
    4.818624,
  // momentumY(23,7, 0-49)
    4.903516, 4.909886, 4.916139, 4.922179, 4.927942, 4.933392, 4.938515, 
    4.943311, 4.947791, 4.951973, 4.955874, 4.959517, 4.96292, 4.966109, 
    4.96911, 4.97011, 4.974067, 4.975875, 4.977278, 4.9785, 4.979634, 
    4.982173, 4.984315, 4.986372, 4.988348, 4.990219, 4.991941, 4.99348, 
    4.994731, 4.995581, 4.995622, 4.996662, 4.996929, 4.996234, 4.994371, 
    4.991102, 4.986189, 4.979417, 4.970619, 4.959719, 4.946767, 4.931982, 
    4.915766, 4.898709, 4.881564, 4.86518, 4.85042, 4.838073, 4.82876, 4.82288,
  // momentumY(23,8, 0-49)
    4.905653, 4.911932, 4.918082, 4.924006, 4.929646, 4.934963, 4.939943, 
    4.944586, 4.948904, 4.952912, 4.956631, 4.960085, 4.963297, 4.966295, 
    4.969112, 4.969871, 4.973276, 4.974898, 4.97614, 4.977212, 4.978214, 
    4.980665, 4.982713, 4.984673, 4.986623, 4.988544, 4.990419, 4.992204, 
    4.99379, 4.994974, 4.995334, 4.996774, 4.997522, 4.997402, 4.996218, 
    4.993746, 4.989747, 4.98399, 4.976279, 4.966488, 4.954601, 4.940746, 
    4.925236, 4.908576, 4.891455, 4.874695, 4.859173, 4.845736, 4.835096, 
    4.827761,
  // momentumY(23,9, 0-49)
    4.908045, 4.914205, 4.920225, 4.926012, 4.931508, 4.936678, 4.941504, 
    4.945988, 4.95014, 4.953975, 4.957514, 4.960781, 4.963801, 4.966605, 
    4.969224, 4.969835, 4.972563, 4.973999, 4.975098, 4.976038, 4.976922, 
    4.979229, 4.981129, 4.982932, 4.984797, 4.986721, 4.988709, 4.99071, 
    4.992615, 4.994116, 4.994787, 4.996551, 4.997704, 4.998085, 4.997517, 
    4.995781, 4.992645, 4.987872, 4.981241, 4.972581, 4.961812, 4.948979, 
    4.934303, 4.918199, 4.901276, 4.884313, 4.868188, 4.853786, 4.841904, 
    4.833155,
  // momentumY(23,10, 0-49)
    4.910669, 4.916684, 4.922551, 4.928182, 4.93352, 4.938529, 4.943195, 
    4.947515, 4.951498, 4.955161, 4.958521, 4.961602, 4.96443, 4.967033, 
    4.969435, 4.969999, 4.971944, 4.973189, 4.97416, 4.974993, 4.975775, 
    4.977887, 4.979592, 4.981181, 4.982915, 4.984797, 4.986864, 4.989058, 
    4.991269, 4.993081, 4.994066, 4.996086, 4.997576, 4.998394, 4.998374, 
    4.997312, 4.994981, 4.991141, 4.985553, 4.978009, 4.968371, 4.956611, 
    4.942855, 4.927424, 4.910847, 4.893844, 4.877275, 4.862051, 4.849038, 
    4.838949,
  // momentumY(23,11, 0-49)
    4.9135, 4.919349, 4.925044, 4.930502, 4.935669, 4.94051, 4.945008, 
    4.94916, 4.952974, 4.956462, 4.959645, 4.96254, 4.965172, 4.967559, 
    4.969719, 4.970341, 4.971409, 4.972464, 4.973328, 4.974075, 4.974782, 
    4.976649, 4.978117, 4.979452, 4.981015, 4.982821, 4.984939, 4.9873, 
    4.989808, 4.991928, 4.993247, 4.995461, 4.997231, 4.998425, 4.998889, 
    4.998437, 4.996847, 4.993878, 4.989277, 4.98281, 4.974285, 4.963607, 
    4.950817, 4.936144, 4.92003, 4.903127, 4.886267, 4.870369, 4.856357, 
    4.845033,
  // momentumY(23,12, 0-49)
    4.916521, 4.922186, 4.927694, 4.932967, 4.937951, 4.942612, 4.946934, 
    4.950913, 4.954554, 4.957866, 4.960867, 4.963572, 4.965996, 4.968154, 
    4.970044, 4.970819, 4.970935, 4.971805, 4.972583, 4.973278, 4.97394, 
    4.975521, 4.976722, 4.97777, 4.979136, 4.98084, 4.982984, 4.985491, 
    4.988282, 4.990713, 4.99239, 4.994746, 4.996741, 4.998255, 4.999147, 
    4.999241, 4.998323, 4.996156, 4.992476, 4.987025, 4.97957, 4.969954, 
    4.958146, 4.944283, 4.928721, 4.912042, 4.895033, 4.878615, 4.863748, 
    4.851315,
  // momentumY(23,13, 0-49)
    4.919718, 4.925189, 4.930497, 4.935571, 4.940359, 4.944829, 4.948966, 
    4.952762, 4.956221, 4.95935, 4.962162, 4.964666, 4.966873, 4.968783, 
    4.970378, 4.971375, 4.97047, 4.971176, 4.971901, 4.972583, 4.97324, 
    4.9745, 4.975414, 4.976161, 4.977314, 4.978903, 4.981051, 4.983681, 
    4.98674, 4.989478, 4.991546, 4.993996, 4.996167, 4.997951, 4.999214, 
    4.999793, 4.999481, 4.998042, 4.995209, 4.990702, 4.984257, 4.975666, 
    4.964827, 4.951798, 4.936854, 4.920501, 4.903476, 4.886686, 4.871117, 
    4.857717,
  // momentumY(23,14, 0-49)
    4.92309, 4.928356, 4.933453, 4.938313, 4.942891, 4.947155, 4.95109, 
    4.954689, 4.957953, 4.960886, 4.963496, 4.96579, 4.967766, 4.969412, 
    4.970696, 4.97194, 4.96995, 4.970529, 4.971247, 4.971963, 4.972665, 
    4.973577, 4.974202, 4.97465, 4.975592, 4.977057, 4.979191, 4.981923, 
    4.985222, 4.988264, 4.990751, 4.99325, 4.995551, 4.997555, 4.999138, 
    5.000143, 5.000372, 4.999589, 4.997525, 4.993887, 4.988383, 4.980763, 
    4.970865, 4.958676, 4.944394, 4.928452, 4.91153, 4.894514, 4.878398, 
    4.864184,
  // momentumY(23,15, 0-49)
    4.926639, 4.931692, 4.936564, 4.941194, 4.945542, 4.949579, 4.95329, 
    4.956672, 4.959722, 4.962442, 4.964838, 4.966904, 4.968638, 4.970015, 
    4.970989, 4.972441, 4.969296, 4.969801, 4.970569, 4.97138, 4.972188, 
    4.972746, 4.973093, 4.973263, 4.974007, 4.975351, 4.977458, 4.980263, 
    4.983772, 4.9871, 4.99003, 4.992534, 4.99492, 4.997099, 4.99895, 
    5.000324, 5.001028, 5.000831, 4.999461, 4.996616, 4.99198, 4.985271, 
    4.976275, 4.96492, 4.95133, 4.93587, 4.919161, 4.902054, 4.885547, 
    4.870674,
  // momentumY(23,16, 0-49)
    4.93037, 4.935199, 4.939828, 4.944206, 4.948298, 4.952079, 4.95554, 
    4.958678, 4.961491, 4.96398, 4.966144, 4.967977, 4.969463, 4.970573, 
    4.971258, 4.972813, 4.968417, 4.968924, 4.969812, 4.970793, 4.971777, 
    4.971989, 4.972089, 4.97202, 4.972597, 4.973833, 4.975907, 4.978754, 
    4.982432, 4.986019, 4.989403, 4.991866, 4.994292, 4.996596, 4.998665, 
    5.000351, 5.00147, 5.001792, 5.001044, 4.998916, 4.995078, 4.989218, 
    4.981081, 4.970545, 4.957668, 4.942747, 4.926349, 4.909281, 4.892532, 
    4.877156,
  // momentumY(23,17, 0-49)
    4.934283, 4.938868, 4.943231, 4.947325, 4.951125, 4.954617, 4.957797, 
    4.960662, 4.963215, 4.965456, 4.967381, 4.968978, 4.970225, 4.971089, 
    4.971526, 4.973015, 4.967241, 4.967832, 4.968923, 4.970154, 4.971397, 
    4.971285, 4.971189, 4.970938, 4.971395, 4.972552, 4.974586, 4.97745, 
    4.981249, 4.985054, 4.988883, 4.991256, 4.99367, 4.99605, 4.998283, 
    5.000228, 5.001703, 5.002481, 5.002286, 5.000806, 4.997698, 4.992626, 
    4.985308, 4.975571, 4.96342, 4.94909, 4.933088, 4.91618, 4.89933, 4.883603,
  // momentumY(23,18, 0-49)
    4.938361, 4.942673, 4.946726, 4.950492, 4.953959, 4.957124, 4.95999, 
    4.962561, 4.964844, 4.966834, 4.968524, 4.969899, 4.970932, 4.971589, 
    4.971833, 4.973045, 4.96572, 4.966478, 4.967849, 4.969416, 4.971005, 
    4.970614, 4.970387, 4.970029, 4.97043, 4.971549, 4.973553, 4.976407, 
    4.980273, 4.98424, 4.988482, 4.990712, 4.993061, 4.995459, 4.9978, 
    4.999946, 5.001716, 5.002888, 5.003185, 5.00229, 4.99985, 4.995514, 
    4.988973, 4.980016, 4.968597, 4.9549, 4.939373, 4.922735, 4.905919, 
    4.889985,
  // momentumY(23,19, 0-49)
    4.942561, 4.94654, 4.950226, 4.953609, 4.956694, 4.959494, 4.962023, 
    4.964293, 4.96631, 4.96807, 4.969558, 4.970748, 4.971611, 4.972114, 
    4.972234, 4.972956, 4.963853, 4.964847, 4.966568, 4.968548, 4.970571, 
    4.969965, 4.969689, 4.969313, 4.969736, 4.970868, 4.972862, 4.97569, 
    4.979569, 4.98363, 4.988221, 4.990247, 4.992464, 4.994816, 4.9972, 
    4.999482, 5.001488, 5.002994, 5.003723, 5.003355, 5.001528, 4.99788, 
    4.992079, 4.983882, 4.973204, 4.960176, 4.945191, 4.928922, 4.912266, 
    4.896266,
  // momentumY(23,20, 0-49)
    4.947812, 4.952392, 4.956592, 4.960402, 4.963821, 4.966853, 4.969504, 
    4.971782, 4.973697, 4.975266, 4.976511, 4.977463, 4.978164, 4.978666, 
    4.97904, 0, 4.962282, 4.963513, 4.965213, 4.966989, 4.9687, 4.967034, 
    4.965853, 4.964697, 4.964581, 4.965442, 4.967443, 4.970533, 4.974926, 
    4.979701, 4.98531, 4.987769, 4.990425, 4.993213, 4.996024, 4.998729, 
    5.001162, 5.003111, 5.004313, 5.004456, 5.003191, 5.000156, 4.995014, 
    4.987504, 4.977509, 4.965121, 4.950686, 4.934827, 4.918398, 4.902422,
  // momentumY(23,21, 0-49)
    4.952321, 4.956649, 4.960524, 4.963956, 4.966967, 4.969578, 4.971817, 
    4.973706, 4.975272, 4.97654, 4.977539, 4.978305, 4.978885, 4.979341, 
    4.979759, 0, 4.957336, 4.958926, 4.96105, 4.963284, 4.965437, 4.96349, 
    4.962173, 4.960936, 4.960859, 4.961868, 4.964108, 4.967514, 4.972302, 
    4.977538, 4.983817, 4.986392, 4.989252, 4.992331, 4.995506, 4.998638, 
    5.001549, 5.004018, 5.005775, 5.006501, 5.005841, 5.003427, 4.99891, 
    4.992016, 4.982603, 4.970729, 4.956704, 4.941106, 4.924758, 4.90866,
  // momentumY(23,22, 0-49)
    4.956862, 4.960968, 4.964542, 4.967612, 4.970216, 4.972399, 4.974205, 
    4.975675, 4.97685, 4.977767, 4.978467, 4.978996, 4.979407, 4.979776, 
    4.98021, 0, 4.953183, 4.955079, 4.957577, 4.960221, 4.962775, 4.960561, 
    4.959106, 4.957771, 4.957701, 4.958802, 4.961205, 4.96483, 4.969896, 
    4.975457, 4.982234, 4.984813, 4.987763, 4.991016, 4.994449, 4.997913, 
    5.001224, 5.004153, 5.00642, 5.0077, 5.007632, 5.005837, 5.001956, 
    4.995699, 4.986902, 4.975594, 4.962046, 4.946799, 4.930641, 4.914544,
  // momentumY(23,23, 0-49)
    4.961319, 4.96523, 4.968522, 4.971242, 4.973449, 4.975204, 4.976571, 
    4.977608, 4.978371, 4.97891, 4.979281, 4.979536, 4.979744, 4.979992, 
    4.980406, 0, 4.949828, 4.951932, 4.954688, 4.957613, 4.960438, 4.957965, 
    4.956351, 4.954892, 4.954782, 4.955913, 4.958411, 4.962177, 4.967437, 
    4.973226, 4.980362, 4.982919, 4.985924, 4.989314, 4.992963, 4.996723, 
    5.000404, 5.00377, 5.006535, 5.008361, 5.008878, 5.007699, 5.004451, 
    4.998827, 4.990645, 4.979904, 4.966846, 4.951975, 4.936047, 4.920007,
  // momentumY(23,24, 0-49)
    4.965569, 4.969304, 4.972334, 4.974724, 4.976551, 4.977893, 4.978831, 
    4.979438, 4.979786, 4.97994, 4.979965, 4.979927, 4.979905, 4.98, 4.98035, 
    0, 4.947584, 4.949786, 4.952665, 4.955732, 4.958699, 4.956051, 4.954333, 
    4.952793, 4.952653, 4.953795, 4.956342, 4.960189, 4.965566, 4.971498, 
    4.97887, 4.981437, 4.984508, 4.988023, 4.991858, 4.995862, 4.999844, 
    5.003561, 5.006723, 5.008988, 5.009978, 5.009296, 5.006564, 5.001464, 
    4.993795, 4.983542, 4.970922, 4.956411, 4.940742, 4.924834,
  // momentumY(23,25, 0-49)
    4.969476, 4.973059, 4.975853, 4.977944, 4.97942, 4.980377, 4.980908, 
    4.981107, 4.981056, 4.98083, 4.980508, 4.980166, 4.979897, 4.979808, 
    4.980052, 0, 4.946215, 4.948393, 4.951257, 4.954316, 4.95728, 4.954575, 
    4.95283, 4.951283, 4.951154, 4.952318, 4.9549, 4.958794, 4.96423, 
    4.970243, 4.97773, 4.980377, 4.983562, 4.987227, 4.991247, 4.995472, 
    4.999707, 5.003707, 5.007178, 5.009773, 5.011113, 5.010795, 5.008437, 
    5.003716, 4.996426, 4.986541, 4.974265, 4.960062, 4.944643, 4.928911,
  // momentumY(23,26, 0-49)
    4.972922, 4.976376, 4.97897, 4.980797, 4.981965, 4.982578, 4.982746, 
    4.982569, 4.982144, 4.981558, 4.980897, 4.980248, 4.979712, 4.979408, 
    4.979493, 0, 4.945743, 4.947777, 4.950482, 4.953379, 4.956195, 4.95355, 
    4.951866, 4.950394, 4.950324, 4.951531, 4.954144, 4.95806, 4.963513, 
    4.969546, 4.977036, 4.979848, 4.983212, 4.987065, 4.991282, 4.995709, 
    5.000151, 5.00436, 5.008039, 5.010841, 5.012385, 5.012269, 5.010112, 
    5.005596, 4.998515, 4.988846, 4.976793, 4.962817, 4.947624, 4.932106,
  // momentumY(23,27, 0-49)
    4.975794, 4.979151, 4.981586, 4.983203, 4.984118, 4.984444, 4.9843, 
    4.983793, 4.983029, 4.982104, 4.981112, 4.980152, 4.979331, 4.978775, 
    4.978641, 0, 4.946302, 4.948066, 4.950467, 4.953045, 4.955564, 4.953069, 
    4.9515, 4.950153, 4.950165, 4.951417, 4.954041, 4.957945, 4.963362, 
    4.969354, 4.976735, 4.979789, 4.983385, 4.987454, 4.991872, 4.996479, 
    5.001076, 5.005418, 5.009205, 5.012092, 5.013698, 5.013628, 5.011506, 
    5.007021, 4.999983, 4.990378, 4.978427, 4.964598, 4.9496, 4.934321,
  // momentumY(23,28, 0-49)
    4.978009, 4.981311, 4.983644, 4.985114, 4.985842, 4.985948, 4.985551, 
    4.984766, 4.983699, 4.982455, 4.981137, 4.979851, 4.978716, 4.977863, 
    4.977447, 0, 4.948286, 4.949656, 4.951609, 4.953715, 4.955791, 4.953478, 
    4.952028, 4.950802, 4.950869, 4.952122, 4.9547, 4.958529, 4.963839, 
    4.969721, 4.97689, 4.98023, 4.984081, 4.988367, 4.992958, 4.997692, 
    5.002371, 5.006748, 5.010526, 5.01336, 5.014878, 5.014691, 5.012437, 
    5.007819, 5.000664, 4.990985, 4.979025, 4.965273, 4.950454, 4.935455,
  // momentumY(23,29, 0-49)
    4.979519, 4.98282, 4.985117, 4.98652, 4.987142, 4.987102, 4.986516, 
    4.985497, 4.984156, 4.982601, 4.980945, 4.979306, 4.977814, 4.976609, 
    4.975844, 0, 4.951502, 4.952365, 4.95373, 4.955213, 4.956685, 4.954491, 
    4.953069, 4.951875, 4.951902, 4.953065, 4.955513, 4.959191, 4.964319, 
    4.970014, 4.976858, 4.980478, 4.984567, 4.989044, 4.993778, 4.998605, 
    5.003326, 5.007692, 5.011411, 5.01414, 5.015511, 5.015141, 5.012679, 
    5.007847, 5.000496, 4.990666, 4.978632, 4.964911, 4.95025, 4.93554,
  // momentumY(23,30, 0-49)
    4.979384, 4.981814, 4.983278, 4.983901, 4.98382, 4.983175, 4.9821, 
    4.980711, 4.979107, 4.977366, 4.975537, 4.973642, 4.971686, 4.969653, 
    4.967526, 4.968501, 4.95388, 4.953983, 4.955086, 4.956669, 4.958492, 
    4.957497, 4.95718, 4.956963, 4.957675, 4.959179, 4.961603, 4.964932, 
    4.969421, 4.974288, 4.980054, 4.983217, 4.986848, 4.990884, 4.995209, 
    4.999662, 5.004045, 5.008105, 5.011535, 5.013987, 5.015082, 5.014435, 
    5.011695, 5.006598, 4.999016, 4.98902, 4.976917, 4.96326, 4.948817, 
    4.934488,
  // momentumY(23,31, 0-49)
    4.979453, 4.981999, 4.983564, 4.984265, 4.984229, 4.983586, 4.982464, 
    4.980983, 4.979244, 4.977332, 4.97531, 4.973215, 4.971061, 4.968839, 
    4.966521, 4.968116, 4.955175, 4.954739, 4.955228, 4.956167, 4.957366, 
    4.956451, 4.956088, 4.955835, 4.956506, 4.958014, 4.960509, 4.963962, 
    4.96857, 4.97352, 4.979156, 4.9828, 4.986884, 4.991324, 4.995992, 
    5.000715, 5.005282, 5.009428, 5.012842, 5.01517, 5.016033, 5.015054, 
    5.011901, 5.006335, 4.99827, 4.987822, 4.975352, 4.961461, 4.94695, 
    4.932743,
  // momentumY(23,32, 0-49)
    4.978727, 4.981336, 4.98298, 4.983766, 4.983811, 4.983236, 4.982162, 
    4.980702, 4.978957, 4.977013, 4.974936, 4.972773, 4.970546, 4.968249, 
    4.965855, 4.967472, 4.956299, 4.9554, 4.955333, 4.955686, 4.956318, 
    4.955542, 4.955204, 4.95499, 4.955684, 4.95724, 4.959817, 4.963375, 
    4.968049, 4.97302, 4.978463, 4.982544, 4.987028, 4.991814, 4.996756, 
    5.001674, 5.006341, 5.010485, 5.013781, 5.015877, 5.016394, 5.014968, 
    5.011288, 5.00515, 4.996514, 4.985552, 4.97268, 4.958555, 4.944016, 
    4.929998,
  // momentumY(23,33, 0-49)
    4.977302, 4.979942, 4.981656, 4.982538, 4.982697, 4.982244, 4.981289, 
    4.979935, 4.97828, 4.976404, 4.974379, 4.972252, 4.970052, 4.967782, 
    4.965415, 4.966619, 4.957237, 4.955972, 4.955427, 4.955264, 4.955398, 
    4.954807, 4.954551, 4.954451, 4.955221, 4.956857, 4.959517, 4.963147, 
    4.967824, 4.972751, 4.977959, 4.982429, 4.987256, 4.992321, 4.997468, 
    5.002501, 5.007183, 5.011227, 5.014306, 5.01606, 5.016119, 5.014136, 
    5.009826, 5.003026, 4.99375, 4.982231, 4.968952, 4.954619, 4.940107, 
    4.926363,
  // momentumY(23,34, 0-49)
    4.975289, 4.977936, 4.979716, 4.98071, 4.981011, 4.98072, 4.979937, 
    4.978752, 4.977258, 4.975528, 4.97363, 4.971616, 4.969521, 4.967354, 
    4.965097, 4.965625, 4.958004, 4.956473, 4.955529, 4.954925, 4.954628, 
    4.954253, 4.954134, 4.954203, 4.955094, 4.956829, 4.959558, 4.963218, 
    4.967833, 4.972657, 4.977599, 4.982405, 4.987512, 4.992789, 4.998067, 
    5.003136, 5.007743, 5.011593, 5.01435, 5.015658, 5.015156, 5.012516, 
    5.007489, 4.99996, 4.990002, 4.977917, 4.964249, 4.94976, 4.935356, 
    4.921988,
  // momentumY(23,35, 0-49)
    4.972805, 4.975446, 4.977287, 4.978399, 4.978864, 4.978765, 4.978192, 
    4.977223, 4.97594, 4.97441, 4.972696, 4.970852, 4.968914, 4.966905, 
    4.964818, 4.964561, 4.958642, 4.956938, 4.955672, 4.954696, 4.954036, 
    4.953892, 4.953948, 4.954236, 4.955279, 4.957119, 4.959894, 4.963537, 
    4.96802, 4.972685, 4.977338, 4.982416, 4.987737, 4.993151, 4.998478, 
    5.003494, 5.007935, 5.011493, 5.013832, 5.014596, 5.013438, 5.010059, 
    5.004251, 4.995952, 4.985302, 4.972674, 4.958676, 4.944117, 4.929926, 
    4.917049,
  // momentumY(23,36, 0-49)
    4.969972, 4.972589, 4.974487, 4.975722, 4.97636, 4.976475, 4.976136, 
    4.975414, 4.974378, 4.973086, 4.971597, 4.969959, 4.968216, 4.966397, 
    4.964516, 4.963494, 4.959198, 4.957397, 4.955878, 4.954597, 4.953636, 
    4.953732, 4.95399, 4.954529, 4.955745, 4.957692, 4.960482, 4.964052, 
    4.968329, 4.972781, 4.977126, 4.9824, 4.987854, 4.993322, 4.99861, 
    5.00348, 5.007657, 5.010827, 5.01265, 5.01278, 5.01089, 5.006711, 
    5.000083, 4.991011, 4.979698, 4.966591, 4.952356, 4.937846, 4.924, 
    4.911744,
  // momentumY(23,37, 0-49)
    4.966919, 4.969494, 4.971436, 4.972788, 4.973604, 4.973938, 4.973849, 
    4.973393, 4.972626, 4.971597, 4.970358, 4.968953, 4.967428, 4.965818, 
    4.964155, 4.96248, 4.959714, 4.957877, 4.956165, 4.954644, 4.953441, 
    4.953775, 4.954249, 4.955064, 4.95646, 4.9585, 4.961268, 4.964707, 
    4.968708, 4.972888, 4.976903, 4.982288, 4.987783, 4.99321, 4.998359, 
    5.002985, 5.006799, 5.009483, 5.010701, 5.010118, 5.007432, 5.002418, 
    4.994967, 4.985151, 4.973249, 4.959768, 4.945435, 4.931123, 4.917774, 
    4.906282,
  // momentumY(23,38, 0-49)
    4.963768, 4.966279, 4.968248, 4.969707, 4.970693, 4.971244, 4.971407, 
    4.971223, 4.970736, 4.969985, 4.969013, 4.967857, 4.966562, 4.96517, 
    4.963725, 4.96156, 4.96023, 4.958398, 4.956545, 4.954842, 4.953458, 
    4.95402, 4.954714, 4.955815, 4.95739, 4.959505, 4.962207, 4.965453, 
    4.969102, 4.972951, 4.976608, 4.982003, 4.987434, 4.992712, 4.997617, 
    5.001892, 5.005239, 5.007343, 5.007872, 5.006511, 5.002993, 4.997136, 
    4.988894, 4.978408, 4.96603, 4.952328, 4.938067, 4.924137, 4.911459, 
    4.90088,
  // momentumY(23,39, 0-49)
    4.960637, 4.963058, 4.965035, 4.96658, 4.967719, 4.968476, 4.968884, 
    4.968968, 4.968763, 4.968296, 4.967598, 4.966702, 4.965645, 4.964471, 
    4.963233, 4.960762, 4.96077, 4.958971, 4.957023, 4.955193, 4.953681, 
    4.954453, 4.955369, 4.956755, 4.958495, 4.960657, 4.963246, 4.966229, 
    4.969455, 4.972909, 4.976169, 4.981458, 4.986709, 4.99172, 4.996265, 
    5.000077, 5.002857, 5.00429, 5.004058, 5.001873, 4.997508, 4.990834, 
    4.981874, 4.970839, 4.958142, 4.944409, 4.930429, 4.917086, 4.905265, 
    4.895751,
  // momentumY(23,40, 0-49)
    4.95763, 4.959937, 4.961891, 4.963499, 4.964767, 4.965711, 4.966346, 
    4.966689, 4.966758, 4.96657, 4.966147, 4.965512, 4.964697, 4.963742, 
    4.962697, 4.960098, 4.961344, 4.959596, 4.957597, 4.95569, 4.954103, 
    4.95507, 4.956193, 4.957851, 4.959733, 4.961905, 4.964325, 4.966981, 
    4.969707, 4.972701, 4.975508, 4.980567, 4.98551, 4.990129, 4.99419, 
    4.997423, 4.999531, 5.000209, 4.99916, 4.996129, 4.990932, 4.983507, 
    4.973942, 4.962516, 4.949704, 4.936168, 4.922704, 4.910172, 4.8994, 
    4.891098,
  // momentumY(23,41, 0-49)
    4.95484, 4.957002, 4.958905, 4.960543, 4.961915, 4.963018, 4.963856, 
    4.964436, 4.964763, 4.964844, 4.96469, 4.964315, 4.963742, 4.963002, 
    4.962139, 4.959574, 4.961953, 4.96027, 4.958256, 4.956322, 4.954705, 
    4.955848, 4.957162, 4.959065, 4.961057, 4.963192, 4.965388, 4.967646, 
    4.9698, 4.972257, 4.974547, 4.979238, 4.983736, 4.987826, 4.991275, 
    4.993814, 4.995153, 4.995003, 4.993098, 4.989223, 4.983247, 4.975173, 
    4.965159, 4.953546, 4.940858, 4.927775, 4.915082, 4.903592, 4.89406, 
    4.887104,
  // momentumY(23,42, 0-49)
    4.952335, 4.954322, 4.956143, 4.957779, 4.959219, 4.960448, 4.961461, 
    4.962251, 4.962814, 4.963148, 4.963252, 4.963131, 4.962798, 4.962269, 
    4.961581, 4.959179, 4.962581, 4.960975, 4.958985, 4.95707, 4.955463, 
    4.956761, 4.958241, 4.960354, 4.962413, 4.964461, 4.966369, 4.96816, 
    4.96967, 4.971512, 4.973205, 4.977383, 4.981291, 4.984713, 4.987421, 
    4.989151, 4.989631, 4.988597, 4.985819, 4.981133, 4.974466, 4.965889, 
    4.955624, 4.944065, 4.931768, 4.919414, 4.907753, 4.897533, 4.889417, 
    4.883925,
  // momentumY(23,43, 0-49)
    4.950162, 4.951948, 4.953654, 4.955253, 4.956722, 4.958042, 4.959195, 
    4.960165, 4.960937, 4.9615, 4.961845, 4.961969, 4.961868, 4.961549, 
    4.961031, 4.958889, 4.963201, 4.961686, 4.959754, 4.957897, 4.956337, 
    4.957767, 4.959386, 4.961664, 4.963741, 4.965644, 4.967198, 4.968454, 
    4.96925, 4.970394, 4.971401, 4.97492, 4.97809, 4.980704, 4.982542, 
    4.983356, 4.982902, 4.980946, 4.977309, 4.971876, 4.964646, 4.955748, 
    4.945463, 4.934228, 4.922611, 4.91127, 4.900899, 4.892162, 4.885618, 
    4.881681,
  // momentumY(23,44, 0-49)
    4.948341, 4.9499, 4.951458, 4.952984, 4.954449, 4.955821, 4.957075, 
    4.958187, 4.959137, 4.959904, 4.96047, 4.960821, 4.960945, 4.960835, 
    4.960487, 4.958665, 4.963771, 4.962362, 4.960526, 4.958759, 4.957273, 
    4.958815, 4.960539, 4.962932, 4.96497, 4.966668, 4.967808, 4.968459, 
    4.968475, 4.968838, 4.96906, 4.971774, 4.974064, 4.975734, 4.976582, 
    4.976389, 4.974941, 4.972054, 4.967598, 4.961523, 4.953889, 4.944887, 
    4.934844, 4.92422, 4.913573, 4.903521, 4.894681, 4.887616, 4.882772, 
    4.88045,
  // momentumY(23,45, 0-49)
    4.946861, 4.948171, 4.949554, 4.950976, 4.952395, 4.95378, 4.955097, 
    4.956316, 4.957407, 4.958346, 4.959108, 4.95967, 4.960007, 4.960099, 
    4.959925, 4.958453, 4.964239, 4.962955, 4.961242, 4.959595, 4.958201, 
    4.959833, 4.961634, 4.964084, 4.966026, 4.967455, 4.968119, 4.968105, 
    4.967281, 4.966781, 4.966122, 4.967893, 4.969166, 4.96977, 4.969526, 
    4.968252, 4.96578, 4.961977, 4.956776, 4.950191, 4.942346, 4.933481, 
    4.923957, 4.914234, 4.904842, 4.896333, 4.889235, 4.883993, 4.880938, 
    4.880261,
  // momentumY(23,46, 0-49)
    4.945683, 4.946728, 4.947913, 4.949197, 4.950539, 4.951898, 4.953238, 
    4.954524, 4.955721, 4.9568, 4.957727, 4.958476, 4.959012, 4.959301, 
    4.959304, 4.958188, 4.964537, 4.963399, 4.961836, 4.96033, 4.959041, 
    4.960747, 4.962584, 4.965035, 4.966822, 4.967922, 4.968055, 4.967322, 
    4.965609, 4.964171, 4.962538, 4.963241, 4.963384, 4.962819, 4.961406, 
    4.959006, 4.955505, 4.950835, 4.944994, 4.938061, 4.930218, 4.921744, 
    4.913013, 4.904469, 4.896591, 4.889844, 4.884655, 4.881347, 4.88013, 
    4.881088,
  // momentumY(23,47, 0-49)
    4.944736, 4.945503, 4.946472, 4.947594, 4.948827, 4.950127, 4.951453, 
    4.952766, 4.954033, 4.955215, 4.956281, 4.957191, 4.957909, 4.958385, 
    4.958569, 4.957788, 4.964588, 4.96362, 4.962227, 4.960876, 4.959701, 
    4.961462, 4.963302, 4.965695, 4.96727, 4.967989, 4.967543, 4.96605, 
    4.96341, 4.960971, 4.958283, 4.957822, 4.956746, 4.954939, 4.952308, 
    4.948769, 4.944271, 4.938815, 4.932464, 4.925364, 4.917743, 4.909908, 
    4.902228, 4.895111, 4.888963, 4.884154, 4.880991, 4.879674, 4.8803, 
    4.882845,
  // momentumY(23,48, 0-49)
    4.943918, 4.9444, 4.945139, 4.946082, 4.947184, 4.948393, 4.949674, 
    4.950984, 4.952284, 4.953536, 4.954707, 4.955752, 4.956629, 4.957283, 
    4.957647, 4.957171, 4.964309, 4.96353, 4.962326, 4.961139, 4.960081, 
    4.961879, 4.963689, 4.965969, 4.967283, 4.967573, 4.966515, 4.964235, 
    4.960649, 4.957168, 4.953364, 4.951672, 4.949322, 4.946239, 4.942382, 
    4.93773, 4.932302, 4.926166, 4.919459, 4.91238, 4.905197, 4.898226, 
    4.891818, 4.886326, 4.882068, 4.87931, 4.878233, 4.878918, 4.881347, 
    4.885399,
  // momentumY(23,49, 0-49)
    4.943139, 4.943075, 4.943346, 4.94389, 4.944658, 4.945593, 4.946653, 
    4.94779, 4.948959, 4.950121, 4.951228, 4.952226, 4.953055, 4.953636, 
    4.953867, 4.95286, 4.96727, 4.965607, 4.963223, 4.960995, 4.959105, 
    4.962934, 4.966742, 4.971398, 4.97398, 4.974425, 4.972114, 4.967323, 
    4.959898, 4.952757, 4.94517, 4.942115, 4.938286, 4.93369, 4.928385, 
    4.922455, 4.916029, 4.909282, 4.902445, 4.895787, 4.889615, 4.884236, 
    4.879951, 4.877014, 4.875607, 4.87583, 4.877696, 4.881118, 4.885932, 
    4.8919,
  // momentumY(24,0, 0-49)
    4.910848, 4.916671, 4.922301, 4.927701, 4.932858, 4.937772, 4.942453, 
    4.946915, 4.951171, 4.955228, 4.959091, 4.962752, 4.9662, 4.969418, 
    4.972382, 4.974842, 4.97764, 4.97967, 4.981387, 4.98284, 4.984052, 
    4.985279, 4.986291, 4.987188, 4.987974, 4.988667, 4.989259, 4.989744, 
    4.990077, 4.99023, 4.990046, 4.989658, 4.988633, 4.986763, 4.983824, 
    4.979576, 4.973786, 4.966261, 4.95687, 4.945582, 4.932493, 4.917852, 
    4.902067, 4.8857, 4.869432, 4.854009, 4.840175, 4.8286, 4.81981, 4.81415,
  // momentumY(24,1, 0-49)
    4.911695, 4.917596, 4.923278, 4.928706, 4.933865, 4.938758, 4.943394, 
    4.94779, 4.951956, 4.955903, 4.959635, 4.963151, 4.96644, 4.969491, 
    4.972285, 4.974345, 4.977362, 4.979176, 4.980673, 4.981947, 4.983039, 
    4.984436, 4.985643, 4.986808, 4.987906, 4.988943, 4.989892, 4.990752, 
    4.991471, 4.992055, 4.9923, 4.992604, 4.992283, 4.991125, 4.988891, 
    4.985327, 4.980186, 4.973246, 4.964348, 4.95343, 4.940554, 4.92594, 
    4.909973, 4.89321, 4.876342, 4.860144, 4.845407, 4.832861, 4.823102, 
    4.816533,
  // momentumY(24,2, 0-49)
    4.912669, 4.91862, 4.924327, 4.929756, 4.934893, 4.93974, 4.944309, 
    4.948617, 4.952674, 4.956494, 4.960084, 4.963445, 4.966572, 4.969456, 
    4.972089, 4.973764, 4.97696, 4.978581, 4.979879, 4.980993, 4.981977, 
    4.983537, 4.984918, 4.986313, 4.987674, 4.988997, 4.990244, 4.99141, 
    4.992443, 4.993364, 4.993931, 4.994814, 4.995092, 4.994552, 4.992957, 
    4.990049, 4.985571, 4.979286, 4.97101, 4.96065, 4.948229, 4.933926, 
    4.918087, 4.901238, 4.884052, 4.867312, 4.851837, 4.8384, 4.827665, 
    4.820106,
  // momentumY(24,3, 0-49)
    4.91381, 4.919782, 4.925487, 4.93089, 4.935981, 4.940762, 4.945244, 
    4.949446, 4.953381, 4.957063, 4.960503, 4.963704, 4.966669, 4.969393, 
    4.971877, 4.973185, 4.976495, 4.977949, 4.979077, 4.98005, 4.980939, 
    4.982646, 4.984173, 4.98575, 4.987319, 4.988866, 4.990348, 4.991757, 
    4.993032, 4.994204, 4.994997, 4.996337, 4.997099, 4.997078, 4.996046, 
    4.993749, 4.98993, 4.984341, 4.976785, 4.967137, 4.955381, 4.941644, 
    4.92622, 4.909581, 4.892362, 4.875326, 4.859296, 4.845084, 4.833405, 
    4.824807,
  // momentumY(24,4, 0-49)
    4.915136, 4.921102, 4.926778, 4.932133, 4.937155, 4.941853, 4.946233, 
    4.950315, 4.954117, 4.957655, 4.960942, 4.963984, 4.966791, 4.969364, 
    4.971712, 4.972683, 4.976027, 4.977337, 4.978322, 4.979175, 4.979979, 
    4.981809, 4.983449, 4.985155, 4.986871, 4.988581, 4.990238, 4.991829, 
    4.993289, 4.994633, 4.995562, 4.997245, 4.998381, 4.99878, 4.998229, 
    4.996487, 4.993301, 4.988431, 4.98166, 4.972841, 4.961918, 4.948961, 
    4.934201, 4.918041, 4.901056, 4.883966, 4.867583, 4.852731, 4.840173, 
    4.830526,
  // momentumY(24,5, 0-49)
    4.916652, 4.922581, 4.928205, 4.933492, 4.938432, 4.943027, 4.947294, 
    4.951252, 4.954916, 4.958307, 4.961441, 4.964331, 4.966985, 4.969419, 
    4.971646, 4.972317, 4.975591, 4.976784, 4.977652, 4.978406, 4.979137, 
    4.981061, 4.982773, 4.984549, 4.986351, 4.988163, 4.989937, 4.99166, 
    4.993255, 4.994709, 4.995702, 4.997621, 4.999029, 4.999756, 4.999607, 
    4.99836, 4.995777, 4.99162, 4.985671, 4.977759, 4.967791, 4.95578, 
    4.941885, 4.926431, 4.909919, 4.893005, 4.876468, 4.861129, 4.847784, 
    4.837109,
  // momentumY(24,6, 0-49)
    4.918346, 4.924214, 4.929765, 4.934965, 4.939806, 4.944293, 4.948441, 
    4.952268, 4.955794, 4.959041, 4.962029, 4.96477, 4.967284, 4.969589, 
    4.971706, 4.972129, 4.975222, 4.976313, 4.97709, 4.977765, 4.978433, 
    4.980412, 4.982152, 4.983939, 4.985767, 4.98762, 4.989464, 4.991274, 
    4.992972, 4.994491, 4.995498, 4.997561, 4.999152, 5.000124, 5.000306, 
    4.999494, 4.997471, 4.994012, 4.988893, 4.98193, 4.972991, 4.96204, 
    4.949162, 4.934595, 4.918754, 4.902222, 4.885718, 4.870051, 4.856028, 
    4.844377,
  // momentumY(24,7, 0-49)
    4.920202, 4.925986, 4.931444, 4.936544, 4.941278, 4.945648, 4.949674, 
    4.953372, 4.956764, 4.959872, 4.962719, 4.965323, 4.967707, 4.969892, 
    4.971903, 4.972137, 4.97493, 4.975934, 4.976643, 4.977257, 4.977875, 
    4.979867, 4.981587, 4.983323, 4.985119, 4.986961, 4.988832, 4.990698, 
    4.992476, 4.994034, 4.995025, 4.997155, 4.998858, 5.000006, 5.000455, 
    5.000026, 4.99852, 4.995724, 4.991423, 4.985418, 4.977546, 4.96772, 
    4.955954, 4.942404, 4.92739, 4.911408, 4.89511, 4.879266, 4.864686, 
    4.852138,
  // momentumY(24,8, 0-49)
    4.922203, 4.927882, 4.933229, 4.938216, 4.942835, 4.947088, 4.95099, 
    4.954564, 4.957827, 4.960806, 4.963521, 4.965996, 4.968257, 4.970326, 
    4.972233, 4.972349, 4.97472, 4.975642, 4.976302, 4.976875, 4.977454, 
    4.979413, 4.981066, 4.982692, 4.984403, 4.986189, 4.988052, 4.989952, 
    4.991802, 4.993388, 4.994358, 4.996493, 4.998249, 4.999518, 5.000184, 
    5.000089, 4.999055, 4.996887, 4.993373, 4.988306, 4.981501, 4.972822, 
    4.962221, 4.949767, 4.935689, 4.92039, 4.904442, 4.888564, 4.873551, 
    4.860202,
  // momentumY(24,9, 0-49)
    4.924329, 4.929885, 4.935111, 4.939977, 4.944474, 4.948607, 4.95239, 
    4.955841, 4.958982, 4.961837, 4.964429, 4.966784, 4.968927, 4.970881, 
    4.972672, 4.972748, 4.974584, 4.975426, 4.976051, 4.9766, 4.977153, 
    4.97903, 4.980568, 4.982034, 4.983612, 4.985303, 4.987132, 4.989051, 
    4.990974, 4.992595, 4.993559, 4.995654, 4.997419, 4.998772, 4.999612, 
    4.999809, 4.999207, 4.997621, 4.994853, 4.990687, 4.98492, 4.977376, 
    4.967946, 4.956625, 4.943548, 4.929025, 4.913544, 4.897759, 4.88244, 
    4.868397,
  // momentumY(24,10, 0-49)
    4.926576, 4.931991, 4.937082, 4.941818, 4.946189, 4.950202, 4.953865, 
    4.957198, 4.960221, 4.962958, 4.965433, 4.967671, 4.969696, 4.971531, 
    4.973192, 4.97331, 4.974496, 4.975257, 4.975863, 4.976406, 4.976948, 
    4.978693, 4.980071, 4.981329, 4.982737, 4.984304, 4.98608, 4.98801, 
    4.990017, 4.99169, 4.992681, 4.994704, 4.996451, 4.997856, 4.998842, 
    4.999298, 4.999086, 4.998041, 4.995966, 4.992651, 4.98787, 4.981419, 
    4.973136, 4.962947, 4.9509, 4.937212, 4.922284, 4.906702, 4.891196, 
    4.876576,
  // momentumY(24,11, 0-49)
    4.928943, 4.934204, 4.939147, 4.943745, 4.947984, 4.95187, 4.955413, 
    4.958628, 4.961534, 4.964156, 4.966515, 4.968637, 4.97054, 4.972244, 
    4.973755, 4.973986, 4.97442, 4.975101, 4.975702, 4.976256, 4.976806, 
    4.978368, 4.97955, 4.980563, 4.981774, 4.983195, 4.984904, 4.986845, 
    4.988947, 4.990697, 4.991765, 4.993696, 4.995408, 4.996849, 4.997957, 
    4.998643, 4.998786, 4.998235, 4.996804, 4.994276, 4.990419, 4.985002, 
    4.977817, 4.968729, 4.957708, 4.944883, 4.930571, 4.91528, 4.899696, 
    4.884621,
  // momentumY(24,12, 0-49)
    4.931442, 4.936534, 4.941318, 4.945765, 4.949864, 4.953617, 4.957031, 
    4.960122, 4.962908, 4.965411, 4.967651, 4.969649, 4.971423, 4.972981, 
    4.974318, 4.974725, 4.974307, 4.974916, 4.975528, 4.976114, 4.976694, 
    4.978027, 4.978982, 4.979725, 4.98072, 4.981984, 4.983621, 4.985569, 
    4.98778, 4.989639, 4.990843, 4.992671, 4.994336, 4.995801, 4.997019, 
    4.997913, 4.998381, 4.998281, 4.997436, 4.995634, 4.992631, 4.988174, 
    4.982021, 4.973984, 4.963962, 4.952005, 4.938346, 4.923423, 4.907864, 
    4.892451,
  // momentumY(24,13, 0-49)
    4.934093, 4.939003, 4.943612, 4.947893, 4.951836, 4.955441, 4.958715, 
    4.961672, 4.964326, 4.966701, 4.968812, 4.970676, 4.972308, 4.973703, 
    4.974848, 4.975464, 4.974095, 4.974648, 4.975296, 4.975943, 4.976576, 
    4.977641, 4.978346, 4.978808, 4.97958, 4.980684, 4.982246, 4.984205, 
    4.986533, 4.988531, 4.989935, 4.991654, 4.993267, 4.994752, 4.996068, 
    4.997155, 4.997918, 4.99823, 4.997921, 4.996779, 4.994556, 4.990984, 
    4.985788, 4.978738, 4.969673, 4.958571, 4.94559, 4.931089, 4.915645, 
    4.900013,
  // momentumY(24,14, 0-49)
    4.936921, 4.94163, 4.946046, 4.950143, 4.953909, 4.957345, 4.96046, 
    4.963262, 4.96577, 4.968, 4.969966, 4.971681, 4.973152, 4.974371, 
    4.975314, 4.976134, 4.973717, 4.97424, 4.974955, 4.975695, 4.976418, 
    4.977182, 4.977629, 4.977811, 4.978366, 4.979317, 4.980805, 4.982772, 
    4.985224, 4.987384, 4.989049, 4.990658, 4.992219, 4.993719, 4.995128, 
    4.996392, 4.997429, 4.998117, 4.998294, 4.997752, 4.996239, 4.993473, 
    4.989157, 4.983024, 4.974865, 4.964593, 4.952296, 4.938266, 4.923021, 
    4.907284,
  // momentumY(24,15, 0-49)
    4.939954, 4.944445, 4.948641, 4.952525, 4.956085, 4.959326, 4.962252, 
    4.964876, 4.967212, 4.969275, 4.971076, 4.972627, 4.973923, 4.974956, 
    4.975694, 4.976676, 4.973099, 4.973635, 4.974455, 4.975329, 4.976182, 
    4.976626, 4.976819, 4.976738, 4.977095, 4.977906, 4.979325, 4.981301, 
    4.983872, 4.986211, 4.988193, 4.98969, 4.991199, 4.992713, 4.994207, 
    4.995636, 4.996924, 4.997959, 4.998579, 4.99858, 4.99771, 4.995675, 
    4.992167, 4.986881, 4.979572, 4.970099, 4.958487, 4.944963, 4.929991, 
    4.914255,
  // momentumY(24,16, 0-49)
    4.943211, 4.947452, 4.951399, 4.955036, 4.958356, 4.961365, 4.964069, 
    4.966485, 4.968622, 4.970495, 4.972114, 4.973482, 4.974594, 4.975438, 
    4.975983, 4.977036, 4.972176, 4.972776, 4.97375, 4.974805, 4.975837, 
    4.975954, 4.975911, 4.9756, 4.975791, 4.976484, 4.977843, 4.979822, 
    4.982503, 4.985028, 4.98737, 4.988751, 4.990204, 4.991729, 4.993303, 
    4.994886, 4.996407, 4.997757, 4.998783, 4.999278, 4.99899, 4.997621, 
    4.994846, 4.990343, 4.983829, 4.97512, 4.964186, 4.9512, 4.936568, 
    4.920935,
  // momentumY(24,17, 0-49)
    4.946694, 4.950654, 4.95431, 4.957654, 4.960692, 4.963429, 4.965877, 
    4.968051, 4.969965, 4.971627, 4.973047, 4.974223, 4.975149, 4.97581, 
    4.976184, 4.977188, 4.970901, 4.971617, 4.972795, 4.974083, 4.975348, 
    4.975148, 4.974903, 4.974407, 4.974476, 4.975085, 4.976398, 4.978378, 
    4.981153, 4.983857, 4.986584, 4.987842, 4.989233, 4.990761, 4.992407, 
    4.994132, 4.995866, 4.997506, 4.998901, 4.999847, 5.000089, 4.999326, 
    4.997222, 4.993437, 4.987666, 4.979686, 4.969424, 4.956998, 4.942767, 
    4.927331,
  // momentumY(24,18, 0-49)
    4.950392, 4.954015, 4.957329, 4.960334, 4.963038, 4.965462, 4.96762, 
    4.969528, 4.9712, 4.972644, 4.973861, 4.974846, 4.975591, 4.976085, 
    4.976321, 4.97714, 4.969261, 4.970144, 4.971568, 4.973141, 4.974692, 
    4.974195, 4.973797, 4.973176, 4.973178, 4.973746, 4.975035, 4.977013, 
    4.97986, 4.982726, 4.985838, 4.986964, 4.988281, 4.9898, 4.991502, 
    4.99335, 4.99528, 4.997187, 4.998922, 5.000279, 5.001005, 5.000793, 
    4.999304, 4.996184, 4.991109, 4.983826, 4.974225, 4.962378, 4.948599, 
    4.933446,
  // momentumY(24,19, 0-49)
    4.954257, 4.957479, 4.960381, 4.962982, 4.965306, 4.967378, 4.969222, 
    4.970854, 4.972284, 4.973517, 4.974545, 4.975358, 4.975943, 4.976294, 
    4.976423, 4.976936, 4.967296, 4.968376, 4.970076, 4.971971, 4.973859, 
    4.973104, 4.972607, 4.971929, 4.971931, 4.972509, 4.973804, 4.975785, 
    4.978683, 4.981678, 4.985153, 4.986128, 4.987349, 4.988836, 4.990572, 
    4.992523, 4.994625, 4.996772, 4.998816, 5.000549, 5.001719, 5.002016, 
    5.001093, 4.99859, 4.994166, 4.98755, 4.978599, 4.967349, 4.954068, 
    4.939276,
  // momentumY(24,20, 0-49)
    4.959174, 4.962858, 4.966164, 4.969108, 4.971708, 4.973982, 4.975949, 
    4.977625, 4.979029, 4.980179, 4.981099, 4.981818, 4.982371, 4.982801, 
    4.983164, 0, 4.964798, 4.966055, 4.967796, 4.969609, 4.971327, 4.969703, 
    4.968443, 4.967083, 4.966592, 4.9669, 4.968161, 4.970348, 4.973696, 
    4.977341, 4.981765, 4.983172, 4.984841, 4.986776, 4.988951, 4.991327, 
    4.993841, 4.996396, 4.998845, 5.000997, 5.002602, 5.003364, 5.002938, 
    5.000969, 4.997112, 4.991087, 4.982724, 4.972033, 4.959246, 4.944842,
  // momentumY(24,21, 0-49)
    4.963408, 4.966722, 4.969628, 4.972158, 4.974346, 4.976221, 4.977811, 
    4.979146, 4.980244, 4.981132, 4.981833, 4.982378, 4.982804, 4.983163, 
    4.983527, 0, 4.959586, 4.9611, 4.963162, 4.96533, 4.967396, 4.965482, 
    4.964082, 4.96265, 4.96222, 4.962704, 4.964239, 4.966779, 4.970561, 
    4.974705, 4.979818, 4.98141, 4.983339, 4.985602, 4.98816, 4.990963, 
    4.993931, 4.996956, 4.999882, 5.002509, 5.004585, 5.00581, 5.005842, 
    5.004326, 5.000915, 4.995324, 4.987371, 4.97705, 4.964567, 4.950371,
  // momentumY(24,22, 0-49)
    4.967702, 4.970664, 4.973182, 4.975305, 4.977076, 4.978538, 4.979732, 
    4.980693, 4.981451, 4.982034, 4.982473, 4.982803, 4.983067, 4.983329, 
    4.983677, 0, 4.955086, 4.956829, 4.959173, 4.961654, 4.964025, 4.961829, 
    4.960271, 4.958739, 4.958321, 4.95891, 4.960636, 4.963431, 4.967537, 
    4.97206, 4.977712, 4.979404, 4.981507, 4.984018, 4.986888, 4.990057, 
    4.993435, 4.9969, 5.000288, 5.003388, 5.00594, 5.007639, 5.008145, 
    5.007098, 5.004148, 4.999008, 4.99149, 4.981569, 4.969436, 4.955513,
  // momentumY(24,23, 0-49)
    4.971951, 4.974577, 4.976721, 4.978443, 4.979802, 4.980852, 4.98164, 
    4.982214, 4.98261, 4.982863, 4.983012, 4.983098, 4.983173, 4.983312, 
    4.983619, 0, 4.951283, 4.953178, 4.955709, 4.958392, 4.960952, 4.958478, 
    4.956745, 4.95508, 4.954624, 4.955256, 4.957099, 4.960074, 4.964422, 
    4.969233, 4.975299, 4.977072, 4.979327, 4.982063, 4.985225, 4.988744, 
    4.992522, 4.996426, 5.000281, 5.003865, 5.006908, 5.009098, 5.010088, 
    5.009516, 5.007031, 5.002338, 4.995245, 4.985715, 4.973922, 4.960277,
  // momentumY(24,24, 0-49)
    4.976042, 4.978349, 4.980137, 4.981477, 4.982438, 4.983085, 4.983476, 
    4.983662, 4.983689, 4.983603, 4.983446, 4.983268, 4.98313, 4.983118, 
    4.983349, 0, 4.948518, 4.95047, 4.953073, 4.955839, 4.958478, 4.955807, 
    4.953943, 4.952183, 4.951692, 4.952342, 4.954256, 4.957346, 4.961858, 
    4.966876, 4.973243, 4.975129, 4.977551, 4.980509, 4.98394, 4.987772, 
    4.991901, 4.996183, 5.000436, 5.004429, 5.007885, 5.010486, 5.011881, 
    5.011705, 5.009609, 5.005295, 4.998567, 4.989384, 4.97791, 4.964542,
  // momentumY(24,25, 0-49)
    4.979859, 4.981875, 4.983335, 4.984321, 4.984909, 4.985174, 4.985183, 
    4.984993, 4.984659, 4.984231, 4.983762, 4.983307, 4.982939, 4.982748, 
    4.982862, 0, 4.94658, 4.948485, 4.951038, 4.953754, 4.956346, 4.953585, 
    4.951666, 4.949878, 4.949385, 4.95006, 4.952026, 4.955197, 4.959819, 
    4.964978, 4.971531, 4.973589, 4.976222, 4.979423, 4.983128, 4.987259, 
    4.991705, 4.996318, 5.000906, 5.005232, 5.009016, 5.011939, 5.013646, 
    5.013772, 5.011967, 5.007938, 5.00149, 4.992584, 4.981378, 4.968261,
  // momentumY(24,26, 0-49)
    4.983298, 4.98506, 4.986228, 4.986894, 4.987146, 4.987062, 4.986718, 
    4.986174, 4.985493, 4.984731, 4.983946, 4.983204, 4.982584, 4.982186, 
    4.982136, 0, 4.945513, 4.947264, 4.949642, 4.952173, 4.954591, 4.951852, 
    4.949958, 4.948216, 4.947764, 4.948481, 4.95049, 4.953713, 4.958396, 
    4.963634, 4.970265, 4.972566, 4.975461, 4.978936, 4.982924, 4.987339, 
    4.992069, 4.996956, 5.001805, 5.006377, 5.010392, 5.013525, 5.015426, 
    5.015734, 5.014105, 5.01025, 5.003979, 4.99526, 4.984254, 4.97135,
  // momentumY(24,27, 0-49)
    4.986259, 4.987812, 4.988739, 4.989136, 4.989098, 4.988709, 4.988045, 
    4.987175, 4.986165, 4.985077, 4.983976, 4.982936, 4.982043, 4.9814, 
    4.981136, 0, 4.94546, 4.946948, 4.949024, 4.951235, 4.95335, 4.950716, 
    4.948902, 4.947252, 4.946861, 4.947614, 4.949643, 4.952878, 4.957563, 
    4.962814, 4.969408, 4.972008, 4.975201, 4.978966, 4.983234, 4.987912, 
    4.99288, 4.997982, 5.003019, 5.007753, 5.011899, 5.015141, 5.017131, 
    5.017511, 5.015946, 5.012156, 5.005963, 4.997341, 4.986464, 4.973726,
  // momentumY(24,28, 0-49)
    4.988665, 4.990068, 4.990814, 4.991004, 4.990735, 4.990089, 4.989146, 
    4.98798, 4.986658, 4.985248, 4.983824, 4.982468, 4.981272, 4.980346, 
    4.979819, 0, 4.946815, 4.947936, 4.949587, 4.951346, 4.953032, 4.950542, 
    4.948813, 4.947252, 4.946893, 4.947637, 4.949623, 4.952797, 4.957403, 
    4.962586, 4.969032, 4.971952, 4.975448, 4.97949, 4.984002, 4.98889, 
    4.994031, 4.999268, 5.004402, 5.0092, 5.013378, 5.016623, 5.018593, 
    5.018941, 5.017337, 5.013512, 5.007304, 4.998701, 4.987891, 4.975283,
  // momentumY(24,29, 0-49)
    4.990462, 4.991789, 4.992432, 4.992489, 4.992052, 4.991203, 4.990024, 
    4.988585, 4.986959, 4.985222, 4.983455, 4.981752, 4.980217, 4.978965, 
    4.978124, 0, 4.949393, 4.950053, 4.951162, 4.952341, 4.953464, 4.951066, 
    4.949343, 4.947788, 4.947369, 4.948007, 4.949859, 4.952889, 4.957327, 
    4.96235, 4.968523, 4.971735, 4.9755, 4.97978, 4.984496, 4.989554, 
    4.994829, 5.000166, 5.005371, 5.010205, 5.014393, 5.01762, 5.019548, 
    5.019832, 5.018151, 5.014245, 5.007967, 4.999325, 4.988527, 4.976,
  // momentumY(24,30, 0-49)
    4.990738, 4.99121, 4.991029, 4.990311, 4.989165, 4.987687, 4.985961, 
    4.984056, 4.982023, 4.979897, 4.977703, 4.975448, 4.973134, 4.970758, 
    4.968334, 4.967433, 4.952801, 4.952506, 4.95306, 4.954014, 4.955168, 
    4.953628, 4.952737, 4.951961, 4.952108, 4.953052, 4.954916, 4.957685, 
    4.961609, 4.965942, 4.971194, 4.974047, 4.977447, 4.981374, 4.985769, 
    4.990544, 4.995582, 5.000725, 5.005774, 5.010484, 5.014568, 5.017704, 
    5.019542, 5.019734, 5.017958, 5.013961, 5.007609, 4.998928, 4.988154, 
    4.975735,
  // momentumY(24,31, 0-49)
    4.991224, 4.991782, 4.991659, 4.990963, 4.989799, 4.988257, 4.986423, 
    4.984369, 4.982151, 4.979816, 4.977396, 4.974913, 4.972373, 4.969775, 
    4.967119, 4.966956, 4.953699, 4.952859, 4.952815, 4.953157, 4.953729, 
    4.952262, 4.951339, 4.950546, 4.950665, 4.951616, 4.953545, 4.956422, 
    4.960444, 4.964846, 4.969977, 4.973281, 4.977116, 4.981448, 4.986209, 
    4.991305, 4.996608, 5.001957, 5.007145, 5.011923, 5.016, 5.01905, 
    5.020725, 5.020681, 5.018607, 5.014267, 5.007555, 4.998531, 4.987468, 
    4.97485,
  // momentumY(24,32, 0-49)
    4.990952, 4.991582, 4.991526, 4.990881, 4.989748, 4.988213, 4.986357, 
    4.984251, 4.981956, 4.979523, 4.976988, 4.974381, 4.971712, 4.968981, 
    4.966177, 4.966247, 4.954534, 4.953211, 4.952619, 4.952398, 4.952437, 
    4.951101, 4.950212, 4.94947, 4.949618, 4.950622, 4.952628, 4.955601, 
    4.959674, 4.964085, 4.969033, 4.97274, 4.976955, 4.98163, 4.986691, 
    4.992035, 4.99753, 5.003008, 5.008257, 5.013021, 5.017007, 5.019885, 
    5.02131, 5.020944, 5.018488, 5.013731, 5.006595, 4.997181, 4.985804, 
    4.972989,
  // momentumY(24,33, 0-49)
    4.989976, 4.990683, 4.990708, 4.990148, 4.98909, 4.987619, 4.985811, 
    4.983734, 4.981448, 4.979006, 4.976447, 4.973802, 4.971087, 4.968307, 
    4.965442, 4.965351, 4.955271, 4.953551, 4.952481, 4.951764, 4.95134, 
    4.950182, 4.949387, 4.948767, 4.949002, 4.950088, 4.952173, 4.955213, 
    4.959281, 4.96364, 4.968359, 4.972418, 4.976954, 4.981907, 4.987197, 
    4.992716, 4.998327, 5.003853, 5.00908, 5.013745, 5.017552, 5.020169, 
    5.021256, 5.020481, 5.017564, 5.012319, 5.004707, 4.994871, 4.983172, 
    4.970181,
  // momentumY(24,34, 0-49)
    4.988362, 4.989154, 4.989285, 4.98884, 4.9879, 4.986543, 4.984841, 
    4.982858, 4.980649, 4.978268, 4.975753, 4.973141, 4.970451, 4.967691, 
    4.964846, 4.964324, 4.955907, 4.953883, 4.95241, 4.951271, 4.950449, 
    4.949511, 4.948865, 4.948426, 4.948793, 4.949985, 4.952144, 4.955214, 
    4.959218, 4.96347, 4.967926, 4.972286, 4.977082, 4.982247, 4.987697, 
    4.993318, 4.998965, 5.004459, 5.009578, 5.014056, 5.017594, 5.019861, 
    5.020521, 5.019255, 5.015803, 5.010012, 5.001885, 4.991614, 4.979609, 
    4.96648,
  // momentumY(24,35, 0-49)
    4.986187, 4.987076, 4.987331, 4.987029, 4.986242, 4.985043, 4.983495, 
    4.981658, 4.979582, 4.977318, 4.974906, 4.972382, 4.969771, 4.967087, 
    4.964324, 4.963235, 4.956457, 4.954219, 4.952422, 4.950934, 4.949782, 
    4.94909, 4.948639, 4.948434, 4.94897, 4.950284, 4.952501, 4.955562, 
    4.959439, 4.963533, 4.967704, 4.972306, 4.977299, 4.98261, 4.988148, 
    4.993796, 4.9994, 5.004778, 5.009702, 5.013903, 5.017081, 5.018907, 
    5.019053, 5.017218, 5.013171, 5.006792, 4.998133, 4.987436, 4.975163, 
    4.961967,
  // momentumY(24,36, 0-49)
    4.983537, 4.98453, 4.984925, 4.98479, 4.984187, 4.983179, 4.981824, 
    4.980174, 4.978276, 4.976174, 4.973908, 4.971516, 4.969026, 4.966462, 
    4.963827, 4.962144, 4.956951, 4.95458, 4.952532, 4.950767, 4.949354, 
    4.948923, 4.9487, 4.948773, 4.949505, 4.950946, 4.953201, 4.956208, 
    4.959899, 4.963787, 4.967659, 4.972442, 4.977566, 4.982953, 4.988503, 
    4.994096, 4.999576, 5.004749, 5.009388, 5.013221, 5.015947, 5.017244, 
    5.016798, 5.014329, 5.009636, 5.002648, 4.993464, 4.982381, 4.969909, 
    4.956739,
  // momentumY(24,37, 0-49)
    4.980508, 4.981606, 4.982151, 4.982196, 4.981798, 4.981007, 4.979875, 
    4.978444, 4.976758, 4.974855, 4.972772, 4.970547, 4.968214, 4.965799, 
    4.963324, 4.9611, 4.957419, 4.954983, 4.952751, 4.950772, 4.949162, 
    4.949, 4.949028, 4.949411, 4.950358, 4.951927, 4.954195, 4.957103, 
    4.96055, 4.96419, 4.967753, 4.97265, 4.977834, 4.983218, 4.988704, 
    4.99416, 4.999428, 5.004307, 5.008569, 5.01194, 5.014123, 5.014809, 
    5.013699, 5.010541, 5.005176, 4.997579, 4.987903, 4.976503, 4.963933, 
    4.950914,
  // momentumY(24,38, 0-49)
    4.977201, 4.978397, 4.979091, 4.979325, 4.979144, 4.978589, 4.977698, 
    4.976512, 4.975065, 4.97339, 4.971519, 4.969489, 4.967337, 4.965096, 
    4.962796, 4.960145, 4.957889, 4.955441, 4.953079, 4.950952, 4.949204, 
    4.949308, 4.949604, 4.950312, 4.951482, 4.953172, 4.955426, 4.958192, 
    4.96134, 4.964695, 4.967939, 4.972879, 4.978047, 4.983353, 4.988689, 
    4.993921, 4.998884, 5.003378, 5.007168, 5.009984, 5.011538, 5.011535, 
    5.0097, 5.005819, 4.999774, 4.991597, 4.981497, 4.96988, 4.957343, 
    4.944621,
  // momentumY(24,39, 0-49)
    4.973715, 4.974999, 4.975837, 4.976258, 4.976297, 4.975984, 4.975348, 
    4.974423, 4.973234, 4.971807, 4.970172, 4.968362, 4.966412, 4.964359, 
    4.962245, 4.959305, 4.958379, 4.955961, 4.953523, 4.9513, 4.949468, 
    4.949832, 4.950396, 4.951439, 4.95283, 4.954629, 4.956837, 4.959415, 
    4.962219, 4.965253, 4.968168, 4.973073, 4.978147, 4.983289, 4.988388, 
    4.993306, 4.997871, 5.001883, 5.005105, 5.007277, 5.00812, 5.007362, 
    5.004759, 5.000136, 4.993432, 4.984732, 4.974305, 4.962605, 4.950256, 
    4.938003,
  // momentumY(24,40, 0-49)
    4.970154, 4.971507, 4.972474, 4.973073, 4.973326, 4.973255, 4.972881, 
    4.972223, 4.971304, 4.970143, 4.968762, 4.967189, 4.965458, 4.963606, 
    4.96168, 4.958601, 4.958908, 4.956546, 4.954076, 4.951808, 4.949941, 
    4.950551, 4.951377, 4.952746, 4.95435, 4.956237, 4.958365, 4.960715, 
    4.96313, 4.96581, 4.968381, 4.973172, 4.978065, 4.982956, 4.987728, 
    4.992238, 4.996309, 4.999742, 5.002305, 5.003745, 5.003803, 5.002235, 
    4.998837, 4.993484, 4.986167, 4.977036, 4.966411, 4.954787, 4.942811, 
    4.931215,
  // momentumY(24,41, 0-49)
    4.966611, 4.968009, 4.969085, 4.969845, 4.970301, 4.970465, 4.970348, 
    4.969962, 4.969318, 4.968431, 4.967318, 4.965998, 4.964501, 4.962861, 
    4.961126, 4.958048, 4.959484, 4.957199, 4.954734, 4.952466, 4.950603, 
    4.951441, 4.952514, 4.954194, 4.955987, 4.957934, 4.959948, 4.96203, 
    4.964015, 4.966311, 4.968513, 4.973105, 4.977732, 4.982281, 4.98663, 
    4.990634, 4.994115, 4.996872, 4.998685, 4.999315, 4.998528, 4.996117, 
    4.99192, 4.985871, 4.978022, 4.96858, 4.957916, 4.946559, 4.935153, 
    4.924411,
  // momentumY(24,42, 0-49)
    4.963175, 4.964589, 4.965748, 4.966649, 4.96729, 4.967675, 4.967805, 
    4.967684, 4.967317, 4.966709, 4.96587, 4.964814, 4.963562, 4.962146, 
    4.960603, 4.957645, 4.960103, 4.957912, 4.955489, 4.953257, 4.951434, 
    4.952474, 4.953773, 4.955733, 4.957686, 4.959659, 4.961521, 4.963294, 
    4.964817, 4.966691, 4.968498, 4.972802, 4.977069, 4.98118, 4.985012, 
    4.988411, 4.991204, 4.993195, 4.994174, 4.993927, 4.992252, 4.988981, 
    4.984013, 4.977334, 4.969066, 4.959468, 4.948955, 4.938068, 4.927447, 
    4.917754,
  // momentumY(24,43, 0-49)
    4.959915, 4.961318, 4.962533, 4.963548, 4.964352, 4.964938, 4.965301, 
    4.965435, 4.965337, 4.965007, 4.964446, 4.963661, 4.962666, 4.96148, 
    4.960136, 4.957391, 4.960761, 4.95868, 4.956325, 4.954162, 4.952404, 
    4.953622, 4.955115, 4.957315, 4.959389, 4.961347, 4.963018, 4.964441, 
    4.965469, 4.966885, 4.968258, 4.972181, 4.975993, 4.979571, 4.982786, 
    4.985485, 4.987495, 4.988636, 4.988711, 4.987537, 4.984951, 4.980837, 
    4.97515, 4.967946, 4.959401, 4.94983, 4.939674, 4.929479, 4.919853, 
    4.911402,
  // momentumY(24,44, 0-49)
    4.956895, 4.958255, 4.959497, 4.960596, 4.961537, 4.962301, 4.962876, 
    4.963249, 4.963411, 4.963352, 4.963067, 4.962556, 4.961821, 4.960875, 
    4.959737, 4.957268, 4.961443, 4.959482, 4.957224, 4.955157, 4.953481, 
    4.954848, 4.956501, 4.958893, 4.961037, 4.962934, 4.964368, 4.965406, 
    4.965909, 4.966825, 4.967713, 4.971162, 4.974424, 4.97737, 4.979871, 
    4.981776, 4.98292, 4.983132, 4.98225, 4.98012, 4.976628, 4.971716, 
    4.965401, 4.957804, 4.949159, 4.93982, 4.930246, 4.920966, 4.912542, 
    4.905505,
  // momentumY(24,45, 0-49)
    4.954153, 4.955442, 4.956679, 4.957835, 4.958883, 4.959798, 4.960562, 
    4.961154, 4.961558, 4.961758, 4.961742, 4.961503, 4.961034, 4.960333, 
    4.959406, 4.957256, 4.962121, 4.960298, 4.958159, 4.956203, 4.954621, 
    4.95611, 4.957882, 4.960408, 4.962569, 4.964353, 4.96551, 4.966124, 
    4.966069, 4.96644, 4.966787, 4.969665, 4.972278, 4.974496, 4.976191, 
    4.977215, 4.977416, 4.976646, 4.974771, 4.971683, 4.967322, 4.961689, 
    4.95487, 4.947047, 4.938503, 4.929619, 4.920855, 4.912706, 4.905671, 
    4.900196,
  // momentumY(24,46, 0-49)
    4.951709, 4.952902, 4.954107, 4.955286, 4.956411, 4.957448, 4.958375, 
    4.959161, 4.959786, 4.960229, 4.960472, 4.960496, 4.96029, 4.959839, 
    4.959132, 4.957314, 4.962758, 4.961088, 4.95909, 4.957263, 4.955777, 
    4.957358, 4.959206, 4.961804, 4.963924, 4.965539, 4.966373, 4.966525, 
    4.965885, 4.965662, 4.965401, 4.967614, 4.969483, 4.970881, 4.971683, 
    4.97175, 4.970951, 4.969162, 4.966289, 4.962273, 4.957111, 4.950871, 
    4.943702, 4.935844, 4.927619, 4.919419, 4.911686, 4.904869, 4.899387, 
    4.895587,
  // momentumY(24,47, 0-49)
    4.949562, 4.950633, 4.951778, 4.952954, 4.954126, 4.955256, 4.956315, 
    4.957269, 4.95809, 4.958755, 4.959237, 4.959513, 4.959562, 4.959362, 
    4.958882, 4.957393, 4.963307, 4.961806, 4.959966, 4.958274, 4.956888, 
    4.958531, 4.960414, 4.963019, 4.965039, 4.966431, 4.966897, 4.96655, 
    4.965296, 4.964425, 4.963489, 4.964943, 4.965979, 4.966473, 4.966308, 
    4.965361, 4.963523, 4.960705, 4.956856, 4.951973, 4.946115, 4.939414, 
    4.932077, 4.924395, 4.916712, 4.90942, 4.902925, 4.897609, 4.893805, 
    4.891757,
  // momentumY(24,48, 0-49)
    4.94768, 4.948614, 4.949677, 4.950824, 4.952013, 4.953206, 4.954365, 
    4.955455, 4.956445, 4.957305, 4.958005, 4.958517, 4.958811, 4.958855, 
    4.958607, 4.95743, 4.963704, 4.962394, 4.960724, 4.959174, 4.957884, 
    4.959568, 4.961443, 4.963991, 4.965849, 4.966964, 4.967022, 4.966144, 
    4.964246, 4.962679, 4.960994, 4.961605, 4.961727, 4.961245, 4.960056, 
    4.958057, 4.95517, 4.951344, 4.946577, 4.940922, 4.934504, 4.927511, 
    4.920208, 4.912917, 4.905994, 4.899813, 4.894729, 4.891049, 4.889009, 
    4.888746,
  // momentumY(24,49, 0-49)
    4.945692, 4.946275, 4.947063, 4.948007, 4.949056, 4.950163, 4.951286, 
    4.952384, 4.953416, 4.954346, 4.955135, 4.95574, 4.956119, 4.956212, 
    4.955952, 4.954215, 4.967573, 4.965439, 4.962609, 4.960008, 4.957872, 
    4.961558, 4.965416, 4.970356, 4.973582, 4.975026, 4.974078, 4.971011, 
    4.965668, 4.960866, 4.955824, 4.955507, 4.954542, 4.952848, 4.950368, 
    4.947054, 4.942887, 4.937885, 4.932127, 4.925748, 4.918957, 4.912019, 
    4.905252, 4.899001, 4.89361, 4.88939, 4.886611, 4.885452, 4.886003, 
    4.888259,
  // momentumY(25,0, 0-49)
    4.925933, 4.931124, 4.936015, 4.940607, 4.944907, 4.948923, 4.952667, 
    4.956147, 4.959369, 4.962331, 4.965029, 4.967461, 4.969619, 4.971503, 
    4.973116, 4.974247, 4.975694, 4.976534, 4.977195, 4.977763, 4.978303, 
    4.97908, 4.979904, 4.98088, 4.98202, 4.983343, 4.984835, 4.986478, 
    4.988221, 4.990023, 4.991735, 4.993485, 4.994883, 4.995748, 4.995881, 
    4.995065, 4.993076, 4.989686, 4.984684, 4.977894, 4.969201, 4.95857, 
    4.946083, 4.931956, 4.916556, 4.9004, 4.884132, 4.868479, 4.854189, 
    4.841959,
  // momentumY(25,1, 0-49)
    4.927026, 4.932236, 4.937124, 4.941692, 4.945944, 4.949895, 4.953556, 
    4.956938, 4.960046, 4.962883, 4.965448, 4.967741, 4.96976, 4.971508, 
    4.972995, 4.97379, 4.975451, 4.976137, 4.976635, 4.977072, 4.977521, 
    4.978458, 4.979441, 4.980615, 4.981967, 4.983503, 4.985191, 4.98702, 
    4.988934, 4.99092, 4.992792, 4.994941, 4.996752, 4.998055, 4.998661, 
    4.998352, 4.996904, 4.994087, 4.98968, 4.983487, 4.975367, 4.965255, 
    4.953193, 4.939358, 4.924083, 4.907857, 4.891315, 4.875189, 4.860251, 
    4.847242,
  // momentumY(25,2, 0-49)
    4.928236, 4.933441, 4.938304, 4.942826, 4.947015, 4.950887, 4.954455, 
    4.95773, 4.960721, 4.963433, 4.965869, 4.968032, 4.969925, 4.971556, 
    4.972939, 4.973425, 4.975278, 4.975841, 4.976205, 4.97653, 4.976901, 
    4.977989, 4.979106, 4.980435, 4.981947, 4.983635, 4.985459, 4.987404, 
    4.989417, 4.991495, 4.993425, 4.995854, 4.997965, 4.999597, 5.000571, 
    5.000686, 4.999723, 4.997451, 4.993648, 4.988107, 4.980661, 4.97122, 
    4.959781, 4.946479, 4.931597, 4.91558, 4.899025, 4.882655, 4.867242, 
    4.853558,
  // momentumY(25,3, 0-49)
    4.929566, 4.934745, 4.939562, 4.944022, 4.948135, 4.951917, 4.955383, 
    4.958548, 4.961421, 4.964013, 4.966328, 4.968372, 4.970154, 4.971688, 
    4.972991, 4.973203, 4.975204, 4.975671, 4.975931, 4.976166, 4.976469, 
    4.977692, 4.978915, 4.980353, 4.981971, 4.983752, 4.985653, 4.987656, 
    4.989704, 4.991798, 4.993697, 4.996298, 4.998598, 5.000453, 5.001705, 
    5.00216, 5.001616, 4.99985, 4.996643, 4.991779, 4.985082, 4.976425, 
    4.965772, 4.953203, 4.938946, 4.923386, 4.907069, 4.890676, 4.874971, 
    4.860731,
  // momentumY(25,4, 0-49)
    4.931008, 4.93614, 4.940896, 4.945281, 4.949308, 4.952993, 4.956354, 
    4.959407, 4.962167, 4.964643, 4.966847, 4.968788, 4.970478, 4.971931, 
    4.973177, 4.973155, 4.975237, 4.975637, 4.975821, 4.975992, 4.976242, 
    4.977576, 4.978874, 4.98037, 4.982038, 4.983856, 4.98578, 4.987794, 
    4.98983, 4.991879, 4.993676, 4.996348, 4.998741, 5.000727, 5.002164, 
    5.002882, 5.002693, 5.001389, 4.998754, 4.994576, 4.988664, 4.980871, 
    4.971121, 4.959445, 4.946002, 4.931112, 4.915251, 4.899047, 4.883229, 
    4.868569,
  // momentumY(25,5, 0-49)
    4.932553, 4.937619, 4.942299, 4.9466, 4.950532, 4.954118, 4.957373, 
    4.960318, 4.962967, 4.965339, 4.967442, 4.969292, 4.970905, 4.9723, 
    4.973505, 4.973295, 4.975376, 4.975733, 4.975873, 4.975999, 4.976211, 
    4.977631, 4.978968, 4.980473, 4.982137, 4.983939, 4.985843, 4.987827, 
    4.98982, 4.991777, 4.993423, 4.996082, 4.998482, 5.000516, 5.002064, 
    5.002976, 5.003079, 5.002186, 5.000093, 4.996589, 4.991478, 4.984593, 
    4.975825, 4.965151, 4.952667, 4.938615, 4.923396, 4.907567, 4.891808, 
    4.876867,
  // momentumY(25,6, 0-49)
    4.934185, 4.93917, 4.943763, 4.94797, 4.951805, 4.955288, 4.95844, 
    4.961281, 4.963829, 4.966102, 4.968116, 4.96989, 4.97144, 4.97279, 
    4.973968, 4.973625, 4.975606, 4.975941, 4.976063, 4.97617, 4.976358, 
    4.977833, 4.979174, 4.980636, 4.982246, 4.983988, 4.985836, 4.987762, 
    4.989691, 4.991532, 4.992995, 4.995569, 4.997908, 4.999924, 5.001517, 
    5.00256, 5.002903, 5.002374, 5.000784, 4.997931, 4.993614, 4.987652, 
    4.979905, 4.970301, 4.958872, 4.945784, 4.931354, 4.916058, 4.900511, 
    4.885429,
  // momentumY(25,7, 0-49)
    4.935893, 4.940784, 4.94528, 4.949388, 4.953124, 4.956505, 4.959556, 
    4.962297, 4.964751, 4.966934, 4.968871, 4.970577, 4.972075, 4.973391, 
    4.974547, 4.974128, 4.975905, 4.976233, 4.976362, 4.976471, 4.976653, 
    4.97815, 4.979456, 4.980828, 4.98234, 4.983981, 4.985743, 4.987593, 
    4.989452, 4.991168, 4.992439, 4.994873, 4.997096, 4.999042, 5.000629, 
    5.001756, 5.002291, 5.002082, 5.000955, 4.998718, 4.995172, 4.990123, 
    4.983405, 4.974901, 4.964583, 4.952542, 4.939005, 4.924366, 4.909166, 
    4.894073,
  // momentumY(25,8, 0-49)
    4.937671, 4.942457, 4.946848, 4.950853, 4.954486, 4.957766, 4.960718, 
    4.963364, 4.965728, 4.96783, 4.969694, 4.971343, 4.972795, 4.974077, 
    4.975214, 4.97478, 4.976242, 4.976571, 4.97673, 4.976866, 4.977058, 
    4.97854, 4.979775, 4.981012, 4.982388, 4.983896, 4.985551, 4.987316, 
    4.98911, 4.990705, 4.991796, 4.994046, 4.996115, 4.997952, 4.999499, 
    5.00067, 5.001359, 5.001431, 5.000728, 4.999069, 4.996257, 4.992092, 
    4.986383, 4.978979, 4.969792, 4.958836, 4.946263, 4.932373, 4.91763, 
    4.902642,
  // momentumY(25,9, 0-49)
    4.939522, 4.944192, 4.948471, 4.952366, 4.955894, 4.959072, 4.961926, 
    4.964479, 4.966755, 4.96878, 4.970574, 4.972166, 4.973575, 4.974823, 
    4.975928, 4.975544, 4.976576, 4.976916, 4.977123, 4.977306, 4.977529, 
    4.978956, 4.980087, 4.981149, 4.982355, 4.983707, 4.985243, 4.986919, 
    4.988662, 4.990154, 4.991093, 4.993133, 4.995021, 4.996726, 4.998206, 
    4.999397, 5.00021, 5.000529, 5.000213, 4.999092, 4.996973, 4.993648, 
    4.988911, 4.982576, 4.974506, 4.964649, 4.953072, 4.939991, 4.92579, 
    4.911009,
  // momentumY(25,10, 0-49)
    4.941456, 4.945998, 4.950157, 4.953936, 4.957352, 4.960425, 4.963178, 
    4.965636, 4.967824, 4.96977, 4.971497, 4.973028, 4.974387, 4.975594, 
    4.976652, 4.976379, 4.976869, 4.977222, 4.977496, 4.977747, 4.978018, 
    4.979352, 4.980344, 4.981201, 4.982213, 4.983394, 4.984804, 4.986394, 
    4.988105, 4.989521, 4.990354, 4.992166, 4.993861, 4.99542, 4.99682, 
    4.998015, 4.998931, 4.999473, 4.999509, 4.998883, 4.997409, 4.994874, 
    4.991057, 4.985744, 4.978755, 4.969977, 4.959402, 4.947165, 4.933567, 
    4.919079,
  // momentumY(25,11, 0-49)
    4.943488, 4.947892, 4.951918, 4.955572, 4.958869, 4.961828, 4.964473, 
    4.96683, 4.968925, 4.970785, 4.972435, 4.973901, 4.975202, 4.976351, 
    4.977344, 4.977236, 4.977071, 4.977445, 4.9778, 4.978139, 4.978481, 
    4.979679, 4.980506, 4.981133, 4.981936, 4.982936, 4.984219, 4.985733, 
    4.98743, 4.988805, 4.98959, 4.991169, 4.992666, 4.994079, 4.995396, 
    4.996587, 4.997594, 4.998336, 4.998695, 4.998528, 4.99765, 4.995848, 
    4.992891, 4.988542, 4.982579, 4.97484, 4.96525, 4.953867, 4.940912, 
    4.926785,
  // momentumY(25,12, 0-49)
    4.94564, 4.949892, 4.953773, 4.957288, 4.960452, 4.963284, 4.965809, 
    4.968053, 4.970044, 4.971808, 4.973372, 4.974759, 4.975985, 4.977059, 
    4.97797, 4.978063, 4.977129, 4.977533, 4.97799, 4.978438, 4.978873, 
    4.979895, 4.980533, 4.980914, 4.981503, 4.982321, 4.983479, 4.984927, 
    4.986634, 4.988007, 4.988809, 4.990157, 4.991462, 4.992733, 4.993971, 
    4.995159, 4.996251, 4.997179, 4.997838, 4.998092, 4.997764, 4.996637, 
    4.994474, 4.991019, 4.986021, 4.979267, 4.970627, 4.960088, 4.947798, 
    4.934089,
  // momentumY(25,13, 0-49)
    4.947933, 4.952016, 4.955732, 4.959089, 4.962103, 4.964792, 4.967181, 
    4.969296, 4.971166, 4.972819, 4.97428, 4.975571, 4.976707, 4.977689, 
    4.978497, 4.978809, 4.976994, 4.977444, 4.978021, 4.978601, 4.979153, 
    4.979963, 4.980396, 4.980526, 4.980901, 4.981544, 4.982584, 4.983975, 
    4.985711, 4.987123, 4.988012, 4.989138, 4.990263, 4.991405, 4.992577, 
    4.993766, 4.994943, 4.996046, 4.996986, 4.997628, 4.997803, 4.997297, 
    4.995863, 4.99323, 4.989122, 4.983292, 4.975555, 4.965837, 4.95422, 
    4.94097,
  // momentumY(25,14, 0-49)
    4.950387, 4.954278, 4.957808, 4.960986, 4.963825, 4.966348, 4.968579, 
    4.970545, 4.972275, 4.973796, 4.975134, 4.976312, 4.977338, 4.97821, 
    4.978907, 4.979425, 4.97661, 4.97713, 4.977851, 4.978589, 4.979284, 
    4.979852, 4.980071, 4.979954, 4.980126, 4.980606, 4.981539, 4.982883, 
    4.984664, 4.98615, 4.987199, 4.988118, 4.989079, 4.990109, 4.991226, 
    4.99243, 4.993695, 4.994971, 4.996171, 4.997174, 4.99781, 4.99787, 
    4.997099, 4.995217, 4.991927, 4.98695, 4.980062, 4.971135, 4.960188, 
    4.947428,
  // momentumY(25,15, 0-49)
    4.953012, 4.956685, 4.960002, 4.96297, 4.965608, 4.967937, 4.969985, 
    4.971778, 4.973346, 4.974717, 4.975914, 4.976958, 4.977856, 4.978607, 
    4.979187, 4.979874, 4.975935, 4.976555, 4.977448, 4.97837, 4.979236, 
    4.979536, 4.979541, 4.979192, 4.97918, 4.979517, 4.980358, 4.981665, 
    4.983503, 4.985093, 4.986369, 4.987097, 4.987914, 4.988852, 4.989933, 
    4.991162, 4.992521, 4.993965, 4.995416, 4.996754, 4.997815, 4.998388, 
    4.998218, 4.997016, 4.99447, 4.990279, 4.98418, 4.976004, 4.965717, 
    4.95347,
  // momentumY(25,16, 0-49)
    4.955808, 4.959229, 4.9623, 4.965026, 4.967431, 4.969538, 4.971376, 
    4.972972, 4.974357, 4.975558, 4.976596, 4.97749, 4.978249, 4.978869, 
    4.979337, 4.980128, 4.974936, 4.975688, 4.976779, 4.977916, 4.978982, 
    4.978996, 4.978796, 4.978239, 4.978075, 4.978295, 4.979061, 4.980342, 
    4.982244, 4.983959, 4.98552, 4.986079, 4.986772, 4.987638, 4.9887, 
    4.989968, 4.99143, 4.993042, 4.994732, 4.996383, 4.997833, 4.998872, 
    4.999245, 4.998656, 4.996783, 4.993306, 4.987936, 4.98047, 4.970826, 
    4.959108,
  // momentumY(25,17, 0-49)
    4.958763, 4.961892, 4.964672, 4.96712, 4.969258, 4.971113, 4.972718, 
    4.974096, 4.975282, 4.976298, 4.977165, 4.9779, 4.978511, 4.979, 
    4.979367, 4.980179, 4.9736, 4.974513, 4.975829, 4.977204, 4.978499, 
    4.97822, 4.977831, 4.977103, 4.976825, 4.976961, 4.977675, 4.978942, 
    4.980911, 4.982769, 4.984655, 4.985065, 4.985654, 4.986466, 4.987527, 
    4.988847, 4.990417, 4.992199, 4.994118, 4.99606, 4.997868, 4.99933, 
    5.000191, 5.000153, 4.998885, 4.996056, 4.991358, 4.984556, 4.975537, 
    4.964358,
  // momentumY(25,18, 0-49)
    4.961843, 4.964629, 4.967072, 4.969197, 4.971034, 4.972611, 4.973962, 
    4.975113, 4.976092, 4.976921, 4.977616, 4.97819, 4.978654, 4.979015, 
    4.979291, 4.980046, 4.971954, 4.973047, 4.974599, 4.976233, 4.977781, 
    4.977211, 4.976659, 4.975799, 4.975451, 4.975545, 4.976236, 4.977504, 
    4.979541, 4.981548, 4.983785, 4.984062, 4.984563, 4.985336, 4.986408, 
    4.98779, 4.989474, 4.991421, 4.993559, 4.995777, 4.997911, 4.999756, 
    5.001056, 5.001511, 5.000786, 4.998543, 4.99446, 4.988282, 4.979865, 
    4.969234,
  // momentumY(25,19, 0-49)
    4.965, 4.967378, 4.969427, 4.971184, 4.972685, 4.973964, 4.975053, 
    4.975977, 4.976758, 4.977411, 4.977946, 4.978371, 4.978695, 4.978937, 
    4.979131, 4.97977, 4.970062, 4.97134, 4.973125, 4.975019, 4.976834, 
    4.975983, 4.975299, 4.974353, 4.973983, 4.974082, 4.974786, 4.976074, 
    4.978185, 4.980337, 4.982932, 4.983087, 4.983509, 4.98425, 4.985336, 
    4.986781, 4.988577, 4.990685, 4.993031, 4.995503, 4.99794, 5.000132, 
    5.001826, 5.002723, 5.002485, 5.000772, 4.997253, 4.991659, 4.983825, 
    4.973745,
  // momentumY(25,20, 0-49)
    4.96907, 4.971853, 4.97428, 4.976379, 4.978179, 4.979703, 4.980981, 
    4.982036, 4.982894, 4.983582, 4.984131, 4.98457, 4.984934, 4.985262, 
    4.9856, 0, 4.967362, 4.968657, 4.970433, 4.97227, 4.973977, 4.972389, 
    4.971055, 4.969516, 4.968708, 4.968553, 4.969211, 4.970665, 4.973172, 
    4.975917, 4.979388, 4.979959, 4.980811, 4.981984, 4.98349, 4.985337, 
    4.98751, 4.989974, 4.992662, 4.995465, 4.99823, 5.000757, 5.002801, 
    5.00407, 5.004237, 5.002963, 4.999919, 4.994827, 4.987511, 4.977941,
  // momentumY(25,21, 0-49)
    4.972409, 4.974806, 4.976856, 4.978595, 4.980055, 4.981269, 4.982268, 
    4.983077, 4.983721, 4.984225, 4.984614, 4.984921, 4.985179, 4.985434, 
    4.985746, 0, 4.962254, 4.963721, 4.965726, 4.967824, 4.969792, 4.9679, 
    4.966414, 4.964807, 4.964072, 4.964111, 4.965068, 4.966903, 4.969873, 
    4.97314, 4.977301, 4.978094, 4.979231, 4.980741, 4.982622, 4.984862, 
    4.987442, 4.990312, 4.993392, 4.996568, 4.999682, 5.002536, 5.004883, 
    5.006442, 5.00689, 5.005895, 5.003135, 4.998338, 4.991322, 4.982051,
  // momentumY(25,22, 0-49)
    4.97575, 4.977777, 4.979461, 4.980845, 4.981971, 4.982874, 4.983584, 
    4.984133, 4.984543, 4.984839, 4.985049, 4.985203, 4.985339, 4.98551, 
    4.985789, 0, 4.957802, 4.959422, 4.961627, 4.96395, 4.966136, 4.963939, 
    4.962275, 4.960557, 4.959836, 4.959994, 4.961162, 4.963283, 4.966613, 
    4.970295, 4.975018, 4.975973, 4.977332, 4.97912, 4.981323, 4.983923, 
    4.986884, 4.990145, 4.993617, 4.997175, 5.000654, 5.003854, 5.006526, 
    5.008392, 5.009137, 5.008434, 5.005967, 5.001472, 4.994767, 4.985815,
  // momentumY(25,23, 0-49)
    4.97903, 4.9807, 4.98203, 4.983072, 4.98387, 4.984463, 4.984885, 
    4.985168, 4.985334, 4.985412, 4.985426, 4.985411, 4.985411, 4.985483, 
    4.985715, 0, 4.953951, 4.955665, 4.95799, 4.960441, 4.962743, 4.960247, 
    4.958386, 4.956528, 4.955769, 4.955982, 4.957291, 4.959627, 4.96324, 
    4.967253, 4.972426, 4.973531, 4.9751, 4.977151, 4.979666, 4.982618, 
    4.98596, 4.98962, 4.993496, 4.997456, 5.001327, 5.004899, 5.007923, 
    5.010116, 5.011169, 5.010761, 5.00858, 5.00437, 4.997954, 4.989296,
  // momentumY(25,24, 0-49)
    4.982182, 4.983513, 4.984507, 4.985221, 4.985703, 4.985996, 4.986135, 
    4.98615, 4.98607, 4.985919, 4.985728, 4.985533, 4.98538, 4.985335, 
    4.985494, 0, 4.951048, 4.95278, 4.955128, 4.957605, 4.959929, 4.957211, 
    4.9552, 4.953234, 4.952438, 4.952682, 4.954084, 4.956569, 4.960389, 
    4.964658, 4.970174, 4.971457, 4.973247, 4.975561, 4.978374, 4.98165, 
    4.985334, 4.989345, 4.993575, 4.997882, 5.002086, 5.005975, 5.009296, 
    5.011769, 5.013084, 5.012925, 5.010993, 5.007029, 5.000869, 4.992476,
  // momentumY(25,25, 0-49)
    4.985147, 4.986164, 4.986844, 4.98725, 4.987433, 4.987438, 4.9873, 
    4.987053, 4.986725, 4.986343, 4.985937, 4.985548, 4.985225, 4.98504, 
    4.985095, 0, 4.948891, 4.950555, 4.952825, 4.955217, 4.957455, 4.95462, 
    4.952531, 4.950522, 4.949719, 4.949996, 4.95147, 4.954067, 4.958037, 
    4.962492, 4.968243, 4.969755, 4.971803, 4.974401, 4.977515, 4.981103, 
    4.985105, 4.989431, 4.993968, 4.998568, 5.003051, 5.007197, 5.010757, 
    5.013449, 5.014969, 5.015006, 5.013266, 5.009499, 5.003544, 4.99537,
  // momentumY(25,26, 0-49)
    4.987865, 4.9886, 4.988998, 4.98912, 4.989028, 4.98876, 4.988358, 
    4.987854, 4.987276, 4.986655, 4.986023, 4.985425, 4.98491, 4.984558, 
    4.98447, 0, 4.947531, 4.949038, 4.951124, 4.95332, 4.955368, 4.952527, 
    4.950438, 4.948456, 4.947687, 4.948007, 4.94954, 4.952215, 4.956279, 
    4.960855, 4.966729, 4.968522, 4.970867, 4.97377, 4.97719, 4.98108, 
    4.985371, 4.989972, 4.994764, 4.999599, 5.004291, 5.008625, 5.01235, 
    5.015193, 5.01685, 5.017016, 5.015405, 5.011773, 5.005966, 4.997958,
  // momentumY(25,27, 0-49)
    4.990288, 4.990781, 4.990932, 4.990807, 4.990461, 4.989943, 4.989286, 
    4.988528, 4.987698, 4.986828, 4.985954, 4.985124, 4.984395, 4.983844, 
    4.983571, 0, 4.947104, 4.948366, 4.950164, 4.952053, 4.953806, 4.951047, 
    4.949018, 4.947112, 4.946393, 4.946748, 4.948308, 4.951011, 4.9551, 
    4.959718, 4.965595, 4.967705, 4.970366, 4.973579, 4.977294, 4.981462, 
    4.986007, 4.990837, 4.995832, 5.000842, 5.005686, 5.010149, 5.013985, 
    5.016919, 5.018657, 5.018899, 5.017364, 5.013811, 5.008099, 5.000204,
  // momentumY(25,28, 0-49)
    4.992364, 4.99267, 4.992622, 4.992288, 4.991722, 4.990971, 4.990073, 
    4.989061, 4.987968, 4.986831, 4.985691, 4.984602, 4.983626, 4.982843, 
    4.982348, 0, 4.947995, 4.94893, 4.950346, 4.951824, 4.953187, 4.950557, 
    4.948601, 4.946773, 4.946075, 4.946415, 4.947931, 4.950579, 4.954597, 
    4.959157, 4.964909, 4.967333, 4.970298, 4.97379, 4.977762, 4.982154, 
    4.986895, 4.991891, 4.997024, 5.002145, 5.00708, 5.011614, 5.015508, 
    5.018489, 5.020265, 5.020542, 5.019038, 5.015524, 5.009858, 5.002028,
  // momentumY(25,29, 0-49)
    4.99406, 4.994244, 4.994057, 4.993563, 4.992815, 4.991854, 4.990718, 
    4.989445, 4.98807, 4.986638, 4.985197, 4.983812, 4.982553, 4.981504, 
    4.980756, 0, 4.950003, 4.95055, 4.951498, 4.952468, 4.953333, 4.950801, 
    4.948859, 4.947036, 4.946271, 4.946498, 4.947872, 4.950364, 4.954204, 
    4.958596, 4.964083, 4.966768, 4.969983, 4.973703, 4.97788, 4.982456, 
    4.98736, 4.992499, 4.997761, 5.002997, 5.008034, 5.012661, 5.016634, 
    5.019682, 5.021515, 5.021831, 5.020354, 5.016856, 5.011202, 5.003389,
  // momentumY(25,30, 0-49)
    4.994519, 4.993861, 4.992861, 4.991597, 4.990131, 4.988516, 4.986785, 
    4.984964, 4.983063, 4.981089, 4.979038, 4.976903, 4.974685, 4.97239, 
    4.970056, 4.968032, 4.954024, 4.95362, 4.953893, 4.954456, 4.955149, 
    4.953227, 4.951905, 4.950692, 4.950378, 4.950848, 4.952226, 4.954489, 
    4.957869, 4.961644, 4.966294, 4.968657, 4.97154, 4.974941, 4.978828, 
    4.983158, 4.987868, 4.99287, 4.998047, 5.00325, 5.008296, 5.012966, 
    5.017006, 5.020132, 5.02204, 5.022424, 5.021001, 5.017544, 5.01192, 
    5.004138,
  // momentumY(25,31, 0-49)
    4.995345, 4.994719, 4.99372, 4.992418, 4.990875, 4.98914, 4.98725, 
    4.985236, 4.983119, 4.98091, 4.978617, 4.976248, 4.9738, 4.97128, 
    4.968707, 4.967444, 4.954495, 4.953582, 4.953315, 4.953332, 4.953514, 
    4.951689, 4.950369, 4.949167, 4.948839, 4.949316, 4.950732, 4.953062, 
    4.956487, 4.960275, 4.964766, 4.967505, 4.970757, 4.974515, 4.978742, 
    4.983388, 4.988389, 4.993653, 4.999059, 5.004455, 5.009655, 5.014433, 
    5.018531, 5.02166, 5.023511, 5.023779, 5.022181, 5.018497, 5.012614, 
    5.004563,
  // momentumY(25,32, 0-49)
    4.995613, 4.995025, 4.99404, 4.992726, 4.991141, 4.989335, 4.987347, 
    4.985208, 4.982944, 4.980573, 4.978112, 4.975571, 4.972955, 4.970267, 
    4.967512, 4.966613, 4.954969, 4.953597, 4.952828, 4.952345, 4.952063, 
    4.950393, 4.949138, 4.948009, 4.947721, 4.948237, 4.949703, 4.952083, 
    4.955504, 4.959243, 4.96351, 4.966569, 4.97013, 4.97418, 4.978678, 
    4.983575, 4.988803, 4.994267, 4.999846, 5.005381, 5.010685, 5.015527, 
    5.019639, 5.022727, 5.024477, 5.024584, 5.022766, 5.018817, 5.01264, 
    5.00429,
  // momentumY(25,33, 0-49)
    4.995334, 4.994799, 4.993851, 4.992554, 4.990967, 4.989133, 4.987097, 
    4.984889, 4.982537, 4.980067, 4.977499, 4.97485, 4.972124, 4.969328, 
    4.966456, 4.965581, 4.955402, 4.953644, 4.952435, 4.951514, 4.95083, 
    4.949367, 4.948236, 4.947248, 4.947051, 4.947638, 4.949155, 4.951556, 
    4.954919, 4.958547, 4.962534, 4.96586, 4.96967, 4.973946, 4.978648, 
    4.983727, 4.989114, 4.994714, 5.000402, 5.006021, 5.011372, 5.016219, 
    5.020291, 5.023284, 5.024884, 5.024779, 5.022697, 5.01844, 5.011938, 
    5.003271,
  // momentumY(25,34, 0-49)
    4.994516, 4.994058, 4.993176, 4.991931, 4.990377, 4.98856, 4.986521, 
    4.984294, 4.981909, 4.979394, 4.976773, 4.974064, 4.971285, 4.968438, 
    4.965515, 4.964412, 4.955777, 4.953714, 4.952136, 4.950844, 4.949824, 
    4.94861, 4.947661, 4.946874, 4.946813, 4.947495, 4.949058, 4.95145, 
    4.954698, 4.95816, 4.961833, 4.965373, 4.969373, 4.97381, 4.978651, 
    4.983845, 4.989325, 4.994994, 5.000727, 5.006361, 5.011694, 5.016483, 
    5.020451, 5.02329, 5.024677, 5.024305, 5.02191, 5.017309, 5.010454, 
    5.001464,
  // momentumY(25,35, 0-49)
    4.993182, 4.992826, 4.992038, 4.990879, 4.989397, 4.987638, 4.985642, 
    4.983441, 4.98107, 4.978556, 4.975928, 4.97321, 4.970424, 4.967576, 
    4.96466, 4.963175, 4.9561, 4.953816, 4.951942, 4.95035, 4.949063, 
    4.948124, 4.947401, 4.946869, 4.946983, 4.94778, 4.949381, 4.95173, 
    4.954807, 4.958058, 4.961395, 4.965098, 4.969231, 4.97377, 4.978685, 
    4.983928, 4.989433, 4.995101, 5.000806, 5.006383, 5.011625, 5.016284, 
    5.020075, 5.022686, 5.023796, 5.023099, 5.02034, 5.015363, 5.008144, 
    4.998838,
  // momentumY(25,36, 0-49)
    4.99136, 4.991127, 4.990465, 4.989424, 4.988052, 4.986389, 4.984475, 
    4.982344, 4.980028, 4.97756, 4.974968, 4.972284, 4.969531, 4.966724, 
    4.963866, 4.961936, 4.956396, 4.953965, 4.951863, 4.950037, 4.948545, 
    4.947903, 4.94744, 4.947205, 4.947526, 4.948452, 4.950078, 4.95235, 
    4.955209, 4.958213, 4.961207, 4.965024, 4.969234, 4.973816, 4.978744, 
    4.983969, 4.989426, 4.995021, 5.000623, 5.006064, 5.011133, 5.01558, 
    5.019113, 5.02142, 5.022179, 5.021094, 5.017928, 5.012548, 5.004965, 
    4.995371,
  // momentumY(25,37, 0-49)
    4.989093, 4.989005, 4.988489, 4.987594, 4.986362, 4.984831, 4.983038, 
    4.981017, 4.9788, 4.976418, 4.973905, 4.97129, 4.968606, 4.965876, 
    4.963112, 4.960749, 4.956685, 4.954175, 4.951907, 4.949906, 4.948266, 
    4.947929, 4.947752, 4.947848, 4.9484, 4.949461, 4.951101, 4.953265, 
    4.955864, 4.958595, 4.961247, 4.96513, 4.969367, 4.973936, 4.978812, 
    4.983953, 4.989293, 4.994737, 5.000153, 5.005373, 5.010181, 5.014324, 
    5.01751, 5.019426, 5.01976, 5.018228, 5.014614, 5.008818, 5.000887, 
    4.991054,
  // momentumY(25,38, 0-49)
    4.986433, 4.986499, 4.986148, 4.985423, 4.98436, 4.982993, 4.981357, 
    4.979482, 4.977402, 4.975144, 4.972745, 4.970237, 4.967655, 4.965031, 
    4.962386, 4.959657, 4.956991, 4.954454, 4.952072, 4.949954, 4.948216, 
    4.948183, 4.948303, 4.948752, 4.949552, 4.950753, 4.952391, 4.954421, 
    4.956728, 4.959168, 4.961491, 4.965396, 4.969607, 4.974107, 4.978873, 
    4.983865, 4.989013, 4.994225, 4.999371, 5.004277, 5.008728, 5.012469, 
    5.015213, 5.016651, 5.016483, 5.014445, 5.010352, 5.00414, 4.995898, 
    4.985897,
  // momentumY(25,39, 0-49)
    4.98344, 4.983667, 4.983495, 4.982955, 4.982084, 4.980909, 4.979459, 
    4.977764, 4.975853, 4.973757, 4.971507, 4.969138, 4.966689, 4.964193, 
    4.961687, 4.95869, 4.957332, 4.954806, 4.952355, 4.950166, 4.948378, 
    4.948637, 4.949059, 4.949871, 4.950925, 4.952264, 4.953889, 4.955763, 
    4.957753, 4.959896, 4.961904, 4.965787, 4.969928, 4.974308, 4.978906, 
    4.983677, 4.988561, 4.99346, 4.998243, 5.002738, 5.006731, 5.009968, 
    5.01217, 5.013039, 5.012294, 5.0097, 5.00511, 4.998499, 4.990002, 4.97993,
  // momentumY(25,40, 0-49)
    4.980185, 4.980569, 4.980579, 4.980239, 4.979576, 4.978613, 4.977376, 
    4.975892, 4.974182, 4.972278, 4.970209, 4.96801, 4.96572, 4.963377, 
    4.961021, 4.957868, 4.957716, 4.955232, 4.952751, 4.950531, 4.948729, 
    4.949263, 4.949982, 4.951154, 4.952459, 4.953933, 4.955529, 4.957229, 
    4.95889, 4.960732, 4.962445, 4.966266, 4.970292, 4.974501, 4.978872, 
    4.983361, 4.987904, 4.992404, 4.996732, 5.000714, 5.004144, 5.006771, 
    5.008329, 5.008542, 5.007154, 5.003967, 4.998874, 4.9919, 4.983227, 
    4.973203,
  // momentumY(25,41, 0-49)
    4.976741, 4.977275, 4.977466, 4.97733, 4.976886, 4.976152, 4.975149, 
    4.973896, 4.972416, 4.970734, 4.968876, 4.966875, 4.964769, 4.962596, 
    4.960401, 4.957204, 4.958153, 4.95573, 4.953249, 4.951032, 4.949247, 
    4.950036, 4.951032, 4.952551, 4.954097, 4.955692, 4.957246, 4.958759, 
    4.960083, 4.96163, 4.963066, 4.966787, 4.970655, 4.974645, 4.978733, 
    4.982875, 4.987002, 4.991017, 4.994792, 4.998161, 5.000918, 5.00283, 
    5.003649, 5.003125, 5.001037, 4.997231, 4.991654, 4.984376, 4.975628, 
    4.965791,
  // momentumY(25,42, 0-49)
    4.973186, 4.973859, 4.974224, 4.97429, 4.974071, 4.973577, 4.972821, 
    4.971821, 4.970592, 4.969154, 4.967532, 4.965755, 4.963854, 4.96187, 
    4.959843, 4.956702, 4.958642, 4.956295, 4.953839, 4.951653, 4.949909, 
    4.950922, 4.952172, 4.954015, 4.955778, 4.957478, 4.958976, 4.96029, 
    4.961278, 4.962534, 4.963706, 4.967291, 4.970962, 4.974685, 4.978436, 
    4.982165, 4.985803, 4.989247, 4.992375, 4.995026, 4.997008, 4.998106, 
    4.998096, 4.996766, 4.993938, 4.989511, 4.983484, 4.975986, 4.967286, 
    4.957791,
  // momentumY(25,43, 0-49)
    4.969604, 4.970394, 4.970921, 4.971184, 4.971187, 4.970936, 4.970438, 
    4.969702, 4.968741, 4.967569, 4.966205, 4.964672, 4.962998, 4.961216, 
    4.959366, 4.956364, 4.959184, 4.95692, 4.954512, 4.952376, 4.950689, 
    4.951897, 4.953369, 4.955495, 4.957449, 4.959227, 4.960651, 4.961758, 
    4.962413, 4.963387, 4.964305, 4.967716, 4.971148, 4.97456, 4.977921, 
    4.981175, 4.984247, 4.987039, 4.989427, 4.991263, 4.992372, 4.992564, 
    4.99165, 4.989461, 4.985876, 4.980847, 4.974436, 4.966821, 4.958312, 
    4.949332,
  // momentumY(25,44, 0-49)
    4.966064, 4.966953, 4.967626, 4.968073, 4.968293, 4.968284, 4.968047, 
    4.967584, 4.966902, 4.966008, 4.964917, 4.963645, 4.962215, 4.960651, 
    4.958984, 4.956183, 4.95977, 4.9576, 4.955254, 4.953185, 4.951562, 
    4.952929, 4.954587, 4.956951, 4.959055, 4.960881, 4.962212, 4.963103, 
    4.963431, 4.964125, 4.96479, 4.967986, 4.971137, 4.974195, 4.977112, 
    4.979828, 4.982265, 4.984324, 4.98589, 4.986822, 4.986973, 4.986184, 
    4.984309, 4.981235, 4.976897, 4.971315, 4.964608, 4.957005, 4.948846, 
    4.940559,
  // momentumY(25,45, 0-49)
    4.962638, 4.963603, 4.964401, 4.965019, 4.965446, 4.965672, 4.965693, 
    4.965505, 4.965105, 4.964497, 4.96369, 4.962691, 4.961516, 4.960183, 
    4.958711, 4.95615, 4.96039, 4.958319, 4.956052, 4.954056, 4.952502, 
    4.953992, 4.955791, 4.95834, 4.960548, 4.962384, 4.963598, 4.964264, 
    4.96427, 4.96468, 4.965085, 4.968025, 4.97085, 4.973502, 4.975922, 
    4.978043, 4.97978, 4.981034, 4.9817, 4.981656, 4.98078, 4.978958, 
    4.976094, 4.972135, 4.967084, 4.961026, 4.954139, 4.946698, 4.939058, 
    4.931637,
  // momentumY(25,46, 0-49)
    4.959384, 4.960401, 4.961304, 4.962074, 4.962692, 4.963142, 4.963412, 
    4.963494, 4.963376, 4.963057, 4.962538, 4.961819, 4.96091, 4.959814, 
    4.958544, 4.956244, 4.961024, 4.959065, 4.956888, 4.954971, 4.95348, 
    4.955057, 4.95695, 4.959622, 4.961882, 4.963686, 4.964756, 4.965185, 
    4.964869, 4.964985, 4.965108, 4.967745, 4.970198, 4.972394, 4.974265, 
    4.975734, 4.97671, 4.977099, 4.976804, 4.975729, 4.973786, 4.970906, 
    4.967056, 4.962245, 4.956552, 4.950125, 4.9432, 4.936079, 4.92913, 
    4.922746,
  // momentumY(25,47, 0-49)
    4.95635, 4.957393, 4.95838, 4.959281, 4.960072, 4.960729, 4.961237, 
    4.961576, 4.961733, 4.961699, 4.961466, 4.961028, 4.960386, 4.959536, 
    4.958477, 4.956443, 4.961648, 4.959813, 4.957735, 4.955901, 4.954465, 
    4.956092, 4.958033, 4.960762, 4.963014, 4.964739, 4.965635, 4.965809, 
    4.965172, 4.964973, 4.964783, 4.967062, 4.969089, 4.970776, 4.972046, 
    4.972809, 4.972975, 4.972452, 4.971157, 4.969021, 4.966, 4.962074, 
    4.957274, 4.951685, 4.945455, 4.938794, 4.931985, 4.925356, 4.919264, 
    4.914069,
  // momentumY(25,48, 0-49)
    4.953563, 4.954612, 4.955658, 4.956668, 4.957611, 4.958456, 4.959181, 
    4.959764, 4.960183, 4.96042, 4.960465, 4.960305, 4.959929, 4.959326, 
    4.958488, 4.956709, 4.96223, 4.960528, 4.958559, 4.956808, 4.955421, 
    4.957064, 4.959004, 4.961722, 4.963907, 4.965501, 4.966192, 4.966093, 
    4.965123, 4.964581, 4.964033, 4.965894, 4.967434, 4.968557, 4.969174, 
    4.969187, 4.968502, 4.967037, 4.964726, 4.961534, 4.957456, 4.952534, 
    4.946867, 4.940608, 4.933976, 4.927238, 4.920715, 4.914744, 4.909664, 
    4.90578,
  // momentumY(25,49, 0-49)
    4.95051, 4.9514, 4.952364, 4.953356, 4.954337, 4.95527, 4.956123, 
    4.956862, 4.957456, 4.957881, 4.95811, 4.958118, 4.957881, 4.957365, 
    4.956535, 4.954092, 4.966395, 4.963832, 4.960638, 4.957756, 4.955451, 
    4.959006, 4.962871, 4.96796, 4.971593, 4.973686, 4.973638, 4.971708, 
    4.96775, 4.964478, 4.961112, 4.962604, 4.963628, 4.964084, 4.963889, 
    4.962953, 4.961198, 4.958563, 4.95502, 4.950583, 4.945317, 4.939349, 
    4.932869, 4.926122, 4.919407, 4.91305, 4.907397, 4.902774, 4.899466, 
    4.897687,
  // momentumY(26,0, 0-49)
    4.94, 4.944391, 4.94844, 4.952157, 4.95555, 4.958627, 4.961393, 4.963849, 
    4.965998, 4.96784, 4.969378, 4.970623, 4.97159, 4.972304, 4.9728, 
    4.972906, 4.973375, 4.973431, 4.973461, 4.973564, 4.973804, 4.974427, 
    4.975248, 4.976345, 4.977716, 4.979355, 4.981232, 4.983315, 4.985551, 
    4.987894, 4.990223, 4.992686, 4.994967, 4.996955, 4.998531, 4.999562, 
    4.999901, 4.999391, 4.997859, 4.995126, 4.991014, 4.985359, 4.978026, 
    4.968945, 4.958121, 4.945682, 4.931883, 4.917126, 4.901945, 4.886976,
  // momentumY(26,1, 0-49)
    4.941255, 4.945621, 4.949628, 4.95329, 4.956614, 4.959611, 4.962287, 
    4.96465, 4.966698, 4.96844, 4.96988, 4.971029, 4.971907, 4.972544, 
    4.972975, 4.97282, 4.973508, 4.973464, 4.973378, 4.973377, 4.973534, 
    4.974285, 4.975206, 4.976415, 4.977892, 4.979619, 4.981553, 4.983666, 
    4.985904, 4.988244, 4.990533, 4.993175, 4.995648, 4.997859, 4.999695, 
    5.00104, 5.001753, 5.001679, 5.000646, 4.998471, 4.994966, 4.989946, 
    4.983253, 4.97478, 4.964502, 4.952498, 4.938988, 4.924335, 4.909052, 
    4.893767,
  // momentumY(26,2, 0-49)
    4.942569, 4.946893, 4.950846, 4.954443, 4.957692, 4.960606, 4.963196, 
    4.965467, 4.967426, 4.969079, 4.970437, 4.971511, 4.972326, 4.97291, 
    4.973302, 4.972916, 4.973806, 4.973686, 4.973504, 4.973412, 4.973489, 
    4.974351, 4.975346, 4.976624, 4.978158, 4.979918, 4.981861, 4.983953, 
    4.986146, 4.988422, 4.990607, 4.993344, 4.995931, 4.998283, 5.000306, 
    5.001887, 5.002901, 5.0032, 5.002613, 5.00096, 4.998045, 4.993671, 
    4.987662, 4.979883, 4.970272, 4.958864, 4.945834, 4.931497, 4.916326, 
    4.900925,
  // momentumY(26,3, 0-49)
    4.943935, 4.948204, 4.952092, 4.955615, 4.958785, 4.961618, 4.964122, 
    4.966311, 4.968189, 4.969768, 4.97106, 4.97208, 4.972853, 4.973409, 
    4.973786, 4.973205, 4.974256, 4.974084, 4.97383, 4.973662, 4.973668, 
    4.974619, 4.975657, 4.976962, 4.978502, 4.98025, 4.982156, 4.984193, 
    4.986302, 4.988472, 4.990499, 4.99326, 4.995889, 4.99831, 5.000443, 
    5.002193, 5.003439, 5.004045, 5.003849, 5.002671, 5.000317, 4.996583, 
    4.991277, 4.984245, 4.975389, 4.964705, 4.952313, 4.938476, 4.923614, 
    4.908288,
  // momentumY(26,4, 0-49)
    4.945349, 4.949549, 4.953363, 4.956806, 4.959896, 4.962646, 4.96507, 
    4.967181, 4.96899, 4.970509, 4.97175, 4.972735, 4.973485, 4.974032, 
    4.974418, 4.973681, 4.974834, 4.974633, 4.974329, 4.974107, 4.97405, 
    4.975069, 4.976121, 4.977407, 4.978909, 4.980601, 4.982437, 4.984389, 
    4.986394, 4.988424, 4.990258, 4.992982, 4.995586, 4.998013, 5.000195, 
    5.002046, 5.003461, 5.004312, 5.004447, 5.003695, 5.001862, 4.998744, 
    4.994145, 4.987888, 4.979846, 4.969979, 4.958351, 4.945166, 4.930783, 
    4.915707,
  // momentumY(26,5, 0-49)
    4.946802, 4.950924, 4.954657, 4.958016, 4.961022, 4.96369, 4.966037, 
    4.968078, 4.969824, 4.971294, 4.9725, 4.973464, 4.974208, 4.974766, 
    4.975174, 4.974328, 4.975505, 4.975296, 4.974972, 4.974713, 4.974607, 
    4.97567, 4.976707, 4.977932, 4.979356, 4.980954, 4.982691, 4.984538, 
    4.986431, 4.988306, 4.989924, 4.992555, 4.995082, 4.997459, 4.999632, 
    5.001528, 5.003053, 5.004092, 5.004505, 5.004128, 5.002773, 5.000243, 
    4.996334, 4.99086, 4.983668, 4.974679, 4.963905, 4.951492, 4.937729, 
    4.923054,
  // momentumY(26,6, 0-49)
    4.948296, 4.952331, 4.955975, 4.959248, 4.962167, 4.964754, 4.967025, 
    4.969, 4.97069, 4.972117, 4.973296, 4.974251, 4.975002, 4.975583, 
    4.976024, 4.975116, 4.97623, 4.976032, 4.975711, 4.975441, 4.975303, 
    4.976385, 4.977377, 4.978502, 4.979811, 4.981283, 4.982903, 4.984636, 
    4.986417, 4.988131, 4.989528, 4.992019, 4.994424, 4.996704, 4.998821, 
    5.000714, 5.002299, 5.003477, 5.004117, 5.004066, 5.00315, 5.001173, 
    4.997931, 4.99323, 4.986898, 4.978821, 4.968964, 4.957409, 4.944374, 
    4.930231,
  // momentumY(26,7, 0-49)
    4.949835, 4.953774, 4.957324, 4.960505, 4.963335, 4.965837, 4.968033, 
    4.96994, 4.971579, 4.972966, 4.974124, 4.975074, 4.97584, 4.976448, 
    4.976927, 4.976012, 4.976964, 4.976792, 4.976501, 4.976244, 4.976095, 
    4.977169, 4.97809, 4.97908, 4.980241, 4.981565, 4.983052, 4.984669, 
    4.986344, 4.987903, 4.98909, 4.991405, 4.993648, 4.995795, 4.997818, 
    4.999667, 5.001273, 5.002547, 5.003373, 5.003607, 5.003088, 5.001628, 
    4.999024, 4.995079, 4.989602, 4.982448, 4.97354, 4.962898, 4.950672, 
    4.93716,
  // momentumY(26,8, 0-49)
    4.951429, 4.955265, 4.958713, 4.961794, 4.96453, 4.966943, 4.969059, 
    4.970898, 4.97248, 4.97383, 4.974967, 4.975914, 4.976696, 4.977333, 
    4.977845, 4.976974, 4.97766, 4.977527, 4.977291, 4.977073, 4.976935, 
    4.977974, 4.978799, 4.979623, 4.980614, 4.98177, 4.983119, 4.98462, 
    4.986207, 4.987626, 4.988623, 4.99073, 4.992783, 4.994769, 4.996668, 
    4.998445, 5.000041, 5.001379, 5.002355, 5.002841, 5.002684, 5.001705, 
    4.99971, 4.99649, 4.991849, 4.985611, 4.97766, 4.967961, 4.956597, 
    4.943792,
  // momentumY(26,9, 0-49)
    4.953088, 4.956812, 4.96015, 4.963123, 4.965757, 4.968074, 4.970102, 
    4.971866, 4.973389, 4.974695, 4.975805, 4.976745, 4.977537, 4.978196, 
    4.978734, 4.97796, 4.97827, 4.978189, 4.978033, 4.97788, 4.97778, 
    4.978755, 4.97946, 4.980095, 4.980895, 4.981874, 4.98308, 4.984471, 
    4.985987, 4.987292, 4.988131, 4.990008, 4.991851, 4.993655, 4.995411, 
    4.997094, 4.998659, 5.000037, 5.00114, 5.001849, 5.002026, 5.001497, 
    5.000074, 4.99755, 4.993714, 4.988372, 4.981369, 4.972619, 4.962144, 
    4.950095,
  // momentumY(26,10, 0-49)
    4.954827, 4.958428, 4.961646, 4.964502, 4.967022, 4.969234, 4.971165, 
    4.972841, 4.974293, 4.975544, 4.97662, 4.977544, 4.978334, 4.979006, 
    4.979555, 4.97893, 4.97875, 4.978733, 4.978679, 4.978618, 4.978583, 
    4.979466, 4.980032, 4.980456, 4.981056, 4.981851, 4.982915, 4.984207, 
    4.985671, 4.986889, 4.987614, 4.989247, 4.990867, 4.992477, 4.99408, 
    4.995658, 4.997178, 4.998582, 4.999794, 5.000707, 5.001192, 5.001086, 
    5.000204, 4.998339, 4.995272, 4.990792, 4.98471, 4.976898, 4.967317, 
    4.956054,
  // momentumY(26,11, 0-49)
    4.956657, 4.960123, 4.963208, 4.965933, 4.968327, 4.970419, 4.972239, 
    4.973818, 4.975185, 4.976367, 4.977395, 4.978288, 4.979064, 4.97973, 
    4.980277, 4.979839, 4.979058, 4.979119, 4.979188, 4.979247, 4.979304, 
    4.980065, 4.980476, 4.980678, 4.981071, 4.981682, 4.982608, 4.983808, 
    4.985242, 4.986406, 4.987069, 4.98845, 4.989841, 4.991255, 4.992701, 
    4.994172, 4.995643, 4.997068, 4.998378, 4.99948, 5.000252, 5.000543, 
    5.00017, 4.998927, 4.996589, 4.992929, 4.987732, 4.98083, 4.972133, 
    4.961664,
  // momentumY(26,12, 0-49)
    4.958586, 4.961901, 4.964838, 4.967417, 4.96967, 4.971628, 4.973322, 
    4.974786, 4.976053, 4.977152, 4.978113, 4.978957, 4.9797, 4.980344, 
    4.98087, 4.980648, 4.979154, 4.979307, 4.979526, 4.97973, 4.979906, 
    4.980518, 4.980759, 4.980734, 4.980921, 4.981354, 4.982149, 4.983266, 
    4.984689, 4.985831, 4.986491, 4.987618, 4.988783, 4.990006, 4.9913, 
    4.992667, 4.994092, 4.995536, 4.996943, 4.998224, 4.99927, 4.999934, 
    5.000038, 4.999378, 4.997725, 4.994837, 4.990478, 4.984446, 4.976607, 
    4.966925,
  // momentumY(26,13, 0-49)
    4.960617, 4.963764, 4.966533, 4.968949, 4.971044, 4.97285, 4.974402, 
    4.975734, 4.976882, 4.97788, 4.978757, 4.979533, 4.980224, 4.980828, 
    4.981322, 4.981328, 4.979001, 4.979272, 4.979662, 4.980037, 4.98036, 
    4.980793, 4.980856, 4.980605, 4.980595, 4.980857, 4.981531, 4.982577, 
    4.984003, 4.985156, 4.985874, 4.986757, 4.987704, 4.988744, 4.989898, 
    4.991172, 4.992559, 4.994028, 4.99553, 4.996988, 4.998293, 4.999307, 
    4.999858, 4.999741, 4.998724, 4.996556, 4.992984, 4.987775, 4.980757, 
    4.971845,
  // momentumY(26,14, 0-49)
    4.962743, 4.965701, 4.968283, 4.970517, 4.972435, 4.974072, 4.975463, 
    4.976647, 4.977662, 4.978541, 4.979313, 4.980003, 4.980623, 4.981172, 
    4.981625, 4.981853, 4.978575, 4.978984, 4.97957, 4.980143, 4.980638, 
    4.980866, 4.980747, 4.980277, 4.980084, 4.980192, 4.980755, 4.98174, 
    4.983183, 4.984377, 4.985216, 4.985863, 4.986608, 4.987482, 4.988513, 
    4.989711, 4.991073, 4.992577, 4.994179, 4.995807, 4.99736, 4.998702, 
    4.999669, 5.000055, 4.999626, 4.998124, 4.995279, 4.99084, 4.984598, 
    4.976427,
  // momentumY(26,15, 0-49)
    4.96495, 4.967693, 4.970068, 4.972099, 4.973822, 4.975271, 4.976488, 
    4.977509, 4.978373, 4.979118, 4.979771, 4.980357, 4.980891, 4.98137, 
    4.981779, 4.982203, 4.977856, 4.978431, 4.979234, 4.980026, 4.980718, 
    4.98072, 4.98042, 4.979746, 4.97939, 4.979363, 4.979831, 4.980763, 
    4.982235, 4.983498, 4.984517, 4.984947, 4.985507, 4.986237, 4.987163, 
    4.988302, 4.989655, 4.991206, 4.992913, 4.99471, 4.996499, 4.998151, 
    4.999502, 5.000349, 5.000455, 4.999561, 4.997384, 4.993657, 4.98814, 
    4.980677,
  // momentumY(26,16, 0-49)
    4.967216, 4.969719, 4.971859, 4.973665, 4.975173, 4.97642, 4.977448, 
    4.978295, 4.979, 4.979597, 4.98012, 4.98059, 4.981026, 4.981429, 4.98179, 
    4.98237, 4.976842, 4.977604, 4.978645, 4.979676, 4.980588, 4.980343, 
    4.979868, 4.979012, 4.978518, 4.978383, 4.978773, 4.979663, 4.981173, 
    4.982527, 4.983779, 4.984013, 4.984412, 4.98502, 4.985863, 4.986963, 
    4.988326, 4.989933, 4.991749, 4.993711, 4.995725, 4.997665, 4.999369, 
    5.000635, 5.001229, 5.000884, 4.999315, 4.996238, 4.991397, 4.984601,
  // momentumY(26,17, 0-49)
    4.969512, 4.97174, 4.973618, 4.975176, 4.976452, 4.977484, 4.978314, 
    4.97898, 4.979518, 4.979966, 4.980352, 4.980701, 4.981031, 4.981352, 
    4.981671, 4.982362, 4.975548, 4.976512, 4.977801, 4.979086, 4.980233, 
    4.979731, 4.979088, 4.978076, 4.977477, 4.977263, 4.977597, 4.978462, 
    4.980017, 4.981482, 4.98301, 4.983071, 4.983333, 4.983841, 4.984626, 
    4.985706, 4.987091, 4.988766, 4.990695, 4.99282, 4.995048, 4.997253, 
    4.999278, 5.000922, 5.001952, 5.002101, 5.001079, 4.998593, 4.994374, 
    4.988206,
  // momentumY(26,18, 0-49)
    4.971802, 4.973717, 4.975297, 4.976582, 4.977609, 4.978417, 4.979047, 
    4.979535, 4.979914, 4.980217, 4.98047, 4.980698, 4.980921, 4.981159, 
    4.981435, 4.982197, 4.974019, 4.975191, 4.976727, 4.978267, 4.979657, 
    4.978886, 4.978089, 4.97695, 4.976281, 4.976023, 4.97633, 4.977189, 
    4.978799, 4.980386, 4.982221, 4.982135, 4.982282, 4.982712, 4.983455, 
    4.984532, 4.985951, 4.9877, 4.989746, 4.992026, 4.994454, 4.996904, 
    4.999218, 5.001203, 5.002622, 5.003211, 5.00268, 5.00073, 4.99708, 
    4.991498,
  // momentumY(26,19, 0-49)
    4.974044, 4.975593, 4.976839, 4.977823, 4.978588, 4.979169, 4.979604, 
    4.979926, 4.980161, 4.980335, 4.98047, 4.980588, 4.98071, 4.980864, 
    4.981096, 4.981905, 4.972337, 4.973706, 4.975469, 4.977249, 4.978876, 
    4.977831, 4.976893, 4.975658, 4.974956, 4.974691, 4.975004, 4.975879, 
    4.977556, 4.979274, 4.981433, 4.981222, 4.981273, 4.981641, 4.982354, 
    4.983438, 4.984897, 4.986722, 4.98888, 4.991309, 4.993922, 4.996593, 
    4.999171, 5.001457, 5.003224, 5.004207, 5.004115, 5.00265, 4.999523, 
    4.994492,
  // momentumY(26,20, 0-49)
    4.977043, 4.979004, 4.980653, 4.982024, 4.983145, 4.984046, 4.984755, 
    4.985302, 4.985719, 4.986032, 4.986275, 4.986479, 4.986677, 4.986904, 
    4.987205, 0, 4.969875, 4.971127, 4.972816, 4.974531, 4.976083, 4.974407, 
    4.972915, 4.971169, 4.97008, 4.969584, 4.969836, 4.970838, 4.972848, 
    4.975082, 4.978014, 4.978158, 4.978577, 4.979314, 4.980385, 4.981804, 
    4.983576, 4.985689, 4.988112, 4.990792, 4.993645, 4.996556, 4.999379, 
    5.001928, 5.003983, 5.005283, 5.005549, 5.004485, 5.001798, 4.997241,
  // momentumY(26,21, 0-49)
    4.97925, 4.980883, 4.98223, 4.983332, 4.984216, 4.984912, 4.985448, 
    4.985849, 4.986141, 4.98635, 4.9865, 4.986621, 4.986745, 4.986916, 
    4.987184, 0, 4.965111, 4.966493, 4.968369, 4.970301, 4.97207, 4.970103, 
    4.968467, 4.966664, 4.965661, 4.965364, 4.965918, 4.967295, 4.969753, 
    4.972483, 4.976055, 4.976404, 4.977072, 4.978096, 4.979475, 4.981217, 
    4.983313, 4.985742, 4.988464, 4.991421, 4.994527, 4.997666, 5.000692, 
    5.003428, 5.005657, 5.007132, 5.007581, 5.006714, 5.004252, 4.999951,
  // momentumY(26,22, 0-49)
    4.981404, 4.982722, 4.983783, 4.984627, 4.985284, 4.985783, 4.986148, 
    4.986403, 4.986568, 4.986663, 4.986715, 4.986749, 4.986797, 4.986908, 
    4.98714, 0, 4.96099, 4.962482, 4.964514, 4.966624, 4.968567, 4.966304, 
    4.964496, 4.962591, 4.961608, 4.961434, 4.962199, 4.963859, 4.966667, 
    4.969792, 4.973887, 4.974385, 4.975251, 4.976512, 4.978163, 4.980196, 
    4.982597, 4.985335, 4.988364, 4.991613, 4.994995, 4.998389, 5.00165, 
    5.004604, 5.007035, 5.008707, 5.009351, 5.008693, 5.006459, 5.002415,
  // momentumY(26,23, 0-49)
    4.983479, 4.984495, 4.985284, 4.985883, 4.986323, 4.986632, 4.986832, 
    4.98694, 4.986977, 4.986959, 4.986909, 4.98685, 4.986816, 4.986859, 
    4.987047, 0, 4.957404, 4.958957, 4.961073, 4.96328, 4.965307, 4.962757, 
    4.96076, 4.958724, 4.957712, 4.957599, 4.958509, 4.960382, 4.963464, 
    4.966908, 4.971419, 4.972058, 4.973106, 4.974591, 4.9765, 4.978821, 
    4.981529, 4.984586, 4.987936, 4.991505, 4.995192, 4.998876, 5.002409, 
    5.00561, 5.008269, 5.010154, 5.011004, 5.010548, 5.008529, 5.004719,
  // momentumY(26,24, 0-49)
    4.985459, 4.986189, 4.98672, 4.987087, 4.98732, 4.987445, 4.987481, 
    4.987444, 4.987351, 4.987216, 4.987059, 4.986901, 4.986779, 4.986742, 
    4.986866, 0, 4.954684, 4.956232, 4.958356, 4.960571, 4.962602, 4.959841, 
    4.957701, 4.955566, 4.954525, 4.954449, 4.955456, 4.957479, 4.960763, 
    4.964447, 4.969274, 4.970074, 4.971316, 4.973023, 4.975178, 4.977761, 
    4.980742, 4.984078, 4.98771, 4.991553, 4.995505, 4.999441, 5.003209, 
    5.006629, 5.009492, 5.011566, 5.012599, 5.012326, 5.010496, 5.006893,
  // momentumY(26,25, 0-49)
    4.987332, 4.987795, 4.988081, 4.988227, 4.98826, 4.988207, 4.988082, 
    4.987899, 4.987672, 4.987413, 4.98714, 4.986873, 4.986648, 4.986516, 
    4.986553, 0, 4.952617, 4.954093, 4.956138, 4.958269, 4.960216, 4.957344, 
    4.955132, 4.95296, 4.95192, 4.951881, 4.952963, 4.955096, 4.958523, 
    4.962382, 4.96742, 4.968424, 4.96989, 4.971837, 4.974241, 4.977078, 
    4.980317, 4.983906, 4.987782, 4.991862, 4.996039, 5.000186, 5.004151, 
    5.007753, 5.010787, 5.013021, 5.014207, 5.014087, 5.012415, 5.008984,
  // momentumY(26,26, 0-49)
    4.989085, 4.989303, 4.989362, 4.989299, 4.989142, 4.988912, 4.988623, 
    4.988289, 4.987917, 4.98752, 4.987116, 4.986723, 4.986379, 4.986131, 
    4.986053, 0, 4.951242, 4.952576, 4.954455, 4.95641, 4.958189, 4.955317, 
    4.953111, 4.950973, 4.949968, 4.949975, 4.951116, 4.953321, 4.956832, 
    4.960795, 4.965936, 4.967187, 4.96891, 4.971114, 4.973774, 4.976858, 
    4.980333, 4.984146, 4.988233, 4.992505, 4.996861, 5.001172, 5.005288, 
    5.009029, 5.012194, 5.014551, 5.015856, 5.015856, 5.014309, 5.011011,
  // momentumY(26,27, 0-49)
    4.990705, 4.990705, 4.990558, 4.990302, 4.989961, 4.989553, 4.989096, 
    4.988595, 4.988062, 4.987507, 4.986948, 4.986408, 4.985921, 4.985535, 
    4.985317, 0, 4.950675, 4.9518, 4.953434, 4.955128, 4.956655, 4.953875, 
    4.951737, 4.949679, 4.948724, 4.948766, 4.949928, 4.952152, 4.955673, 
    4.959657, 4.964782, 4.966302, 4.968293, 4.970756, 4.97366, 4.976973, 
    4.980659, 4.984664, 4.988923, 4.993354, 4.997853, 5.002294, 5.00653, 
    5.010384, 5.013654, 5.016113, 5.017517, 5.017615, 5.016166, 5.012967,
  // momentumY(26,28, 0-49)
    4.992178, 4.991997, 4.991673, 4.991239, 4.990721, 4.990136, 4.989495, 
    4.988809, 4.988087, 4.987344, 4.9866, 4.985881, 4.985225, 4.984678, 
    4.984301, 0, 4.951277, 4.95214, 4.953459, 4.954813, 4.956015, 4.953386, 
    4.95134, 4.949368, 4.948436, 4.948458, 4.949565, 4.951716, 4.955142, 
    4.959041, 4.964017, 4.965793, 4.968029, 4.970719, 4.973828, 4.977328, 
    4.981176, 4.985326, 4.989712, 4.994259, 4.998865, 5.003407, 5.007742, 
    5.011695, 5.015062, 5.017617, 5.019115, 5.019303, 5.017936, 5.014811,
  // momentumY(26,29, 0-49)
    4.993492, 4.993173, 4.992706, 4.992117, 4.991431, 4.990662, 4.989821, 
    4.98892, 4.987972, 4.987, 4.986029, 4.985097, 4.984242, 4.98352, 
    4.982977, 0, 4.952824, 4.953395, 4.954348, 4.955293, 4.95609, 4.953598, 
    4.951597, 4.949647, 4.948653, 4.948557, 4.949506, 4.951476, 4.95469, 
    4.958384, 4.963066, 4.965036, 4.967458, 4.970321, 4.97359, 4.977238, 
    4.981226, 4.985511, 4.990031, 4.994714, 4.999458, 5.004147, 5.00863, 
    5.012733, 5.016247, 5.018942, 5.020564, 5.020856, 5.019571, 5.016503,
  // momentumY(26,30, 0-49)
    4.99386, 4.992723, 4.991463, 4.990121, 4.988725, 4.987293, 4.985828, 
    4.984329, 4.982784, 4.98118, 4.979504, 4.977741, 4.975895, 4.973988, 
    4.972077, 4.969747, 4.956999, 4.956827, 4.957161, 4.957656, 4.958186, 
    4.95614, 4.954606, 4.953129, 4.952481, 4.952558, 4.953475, 4.955208, 
    4.957977, 4.961077, 4.964963, 4.966609, 4.968697, 4.971236, 4.974212, 
    4.977611, 4.981407, 4.985562, 4.990018, 4.994699, 4.999503, 5.004301, 
    5.008934, 5.013212, 5.016919, 5.019805, 5.021607, 5.022055, 5.020894, 
    5.017915,
  // momentumY(26,31, 0-49)
    4.994776, 4.99362, 4.992315, 4.990895, 4.989389, 4.987814, 4.986178, 
    4.984484, 4.982728, 4.980905, 4.979011, 4.977039, 4.974996, 4.972894, 
    4.97077, 4.969105, 4.957089, 4.956472, 4.956341, 4.956375, 4.956476, 
    4.954564, 4.953073, 4.951636, 4.950986, 4.951061, 4.95199, 4.953743, 
    4.956496, 4.959546, 4.963222, 4.965158, 4.96754, 4.970372, 4.973639, 
    4.977323, 4.981398, 4.985823, 4.99054, 4.995468, 5.000506, 5.005515, 
    5.010334, 5.014765, 5.01858, 5.021528, 5.023334, 5.023723, 5.022443, 
    5.01929,
  // momentumY(26,32, 0-49)
    4.995375, 4.994205, 4.99286, 4.991376, 4.989777, 4.988082, 4.986303, 
    4.984447, 4.982514, 4.980509, 4.978431, 4.976282, 4.974068, 4.971794, 
    4.969482, 4.968209, 4.95724, 4.956205, 4.955632, 4.955235, 4.954943, 
    4.953212, 4.951815, 4.950471, 4.949865, 4.949964, 4.950908, 4.952662, 
    4.955353, 4.958293, 4.961698, 4.963876, 4.966497, 4.969563, 4.973063, 
    4.976978, 4.981282, 4.985934, 4.990874, 4.996023, 5.001267, 5.006473, 
    5.011462, 5.016034, 5.019948, 5.022943, 5.024738, 5.025053, 5.023633, 
    5.020279,
  // momentumY(26,33, 0-49)
    4.995639, 4.99447, 4.9931, 4.991568, 4.989897, 4.988105, 4.98621, 
    4.984221, 4.982143, 4.979988, 4.97776, 4.975465, 4.973111, 4.970702, 
    4.968242, 4.967098, 4.957392, 4.955994, 4.955024, 4.954244, 4.95361, 
    4.952107, 4.950858, 4.949664, 4.949143, 4.949293, 4.950252, 4.951982, 
    4.954559, 4.957333, 4.960416, 4.962787, 4.965594, 4.96884, 4.972515, 
    4.976605, 4.981087, 4.985918, 4.991039, 4.996368, 5.001789, 5.007158, 
    5.012293, 5.01698, 5.020972, 5.023992, 5.025752, 5.025967, 5.02438, 
    5.020803,
  // momentumY(26,34, 0-49)
    4.995543, 4.994396, 4.993027, 4.99147, 4.98975, 4.98789, 4.985905, 
    4.983811, 4.98162, 4.979345, 4.976997, 4.97459, 4.97213, 4.969624, 
    4.967066, 4.965834, 4.957517, 4.955821, 4.954513, 4.953405, 4.952485, 
    4.951245, 4.95019, 4.9492, 4.948807, 4.949031, 4.950005, 4.951681, 
    4.954097, 4.956656, 4.959386, 4.961906, 4.964849, 4.968222, 4.972019, 
    4.97623, 4.980836, 4.985796, 4.991051, 4.996513, 5.002068, 5.007562, 
    5.012805, 5.017571, 5.021602, 5.024612, 5.026301, 5.026382, 5.024599, 
    5.020772,
  // momentumY(26,35, 0-49)
    4.995066, 4.99397, 4.992628, 4.991074, 4.989336, 4.987434, 4.985391, 
    4.983224, 4.98095, 4.978586, 4.976151, 4.97366, 4.971129, 4.968563, 
    4.965956, 4.964484, 4.957617, 4.955689, 4.954103, 4.952727, 4.951577, 
    4.950626, 4.949806, 4.949069, 4.948839, 4.949157, 4.950138, 4.951736, 
    4.953943, 4.956252, 4.958614, 4.961243, 4.964278, 4.967728, 4.971596, 
    4.975876, 4.980554, 4.985588, 4.990923, 4.996468, 5.002102, 5.007667, 
    5.012964, 5.017759, 5.02178, 5.024729, 5.026304, 5.026208, 5.024194, 
    5.02009,
  // momentumY(26,36, 0-49)
    4.99419, 4.993175, 4.991889, 4.99037, 4.988643, 4.986734, 4.984667, 
    4.98246, 4.980136, 4.977716, 4.975226, 4.972688, 4.970117, 4.967527, 
    4.964915, 4.96312, 4.957703, 4.95561, 4.953803, 4.952217, 4.950887, 
    4.950241, 4.949687, 4.949242, 4.949209, 4.949636, 4.95062, 4.952115, 
    4.954077, 4.95611, 4.958105, 4.960808, 4.963894, 4.967376, 4.971268, 
    4.975566, 4.98026, 4.985313, 4.990666, 4.996232, 5.001882, 5.007453, 
    5.012741, 5.017495, 5.021441, 5.024268, 5.025669, 5.02535, 5.023067, 
    5.018667,
  // momentumY(26,37, 0-49)
    4.992908, 4.991998, 4.9908, 4.989348, 4.987668, 4.985786, 4.983728, 
    4.981519, 4.979182, 4.976744, 4.974233, 4.971678, 4.969099, 4.966518, 
    4.963937, 4.961798, 4.957793, 4.955594, 4.953619, 4.951871, 4.950411, 
    4.950073, 4.949806, 4.949687, 4.949876, 4.950426, 4.951407, 4.952781, 
    4.954471, 4.956215, 4.957856, 4.9606, 4.963703, 4.967181, 4.971049, 
    4.975317, 4.979972, 4.984982, 4.990291, 4.995806, 5.001399, 5.006898, 
    5.012094, 5.01673, 5.020518, 5.023149, 5.024311, 5.023713, 5.021127, 
    5.016415,
  // momentumY(26,38, 0-49)
    4.991222, 4.990443, 4.98936, 4.988006, 4.986406, 4.984589, 4.98258, 
    4.980407, 4.978095, 4.975675, 4.97318, 4.970641, 4.968087, 4.965544, 
    4.963021, 4.960566, 4.957904, 4.955646, 4.953547, 4.951684, 4.950138, 
    4.950104, 4.950134, 4.950362, 4.950793, 4.951478, 4.952455, 4.953692, 
    4.955092, 4.956546, 4.957858, 4.960621, 4.96371, 4.967146, 4.970952, 
    4.975142, 4.979702, 4.98461, 4.989802, 4.995189, 5.000639, 5.005978, 
    5.010987, 5.015409, 5.01895, 5.021299, 5.022146, 5.021213, 5.018287, 
    5.013258,
  // momentumY(26,39, 0-49)
    4.989146, 4.988517, 4.987576, 4.98635, 4.984865, 4.983149, 4.981227, 
    4.979128, 4.976882, 4.974522, 4.972079, 4.969591, 4.967091, 4.96461, 
    4.962165, 4.959454, 4.95805, 4.955768, 4.953585, 4.951646, 4.950048, 
    4.950306, 4.950636, 4.951224, 4.951909, 4.952735, 4.953708, 4.954801, 
    4.955904, 4.957078, 4.958095, 4.960857, 4.963908, 4.967274, 4.970981, 
    4.975045, 4.979459, 4.984196, 4.9892, 4.994374, 4.999588, 5.004664, 
    5.009383, 5.013483, 5.016672, 5.018644, 5.019099, 5.017773, 5.014479, 
    5.009132,
  // momentumY(26,40, 0-49)
    4.986707, 4.986245, 4.985466, 4.984396, 4.983058, 4.981478, 4.979682, 
    4.977698, 4.975558, 4.973294, 4.970941, 4.968537, 4.966121, 4.963724, 
    4.961371, 4.958483, 4.95824, 4.95596, 4.953722, 4.951737, 4.950122, 
    4.950653, 4.951275, 4.952221, 4.953166, 4.954142, 4.955109, 4.956059, 
    4.956869, 4.957781, 4.958541, 4.961287, 4.964283, 4.967553, 4.97113, 
    4.975026, 4.979239, 4.983742, 4.988476, 4.993349, 4.998224, 5.002929, 
    5.007241, 5.010903, 5.013631, 5.015126, 5.015107, 5.013333, 5.009647, 
    5.004004,
  // momentumY(26,41, 0-49)
    4.983946, 4.983662, 4.983064, 4.982172, 4.981009, 4.979598, 4.977962, 
    4.976132, 4.974137, 4.972007, 4.969779, 4.967493, 4.965187, 4.962894, 
    4.960647, 4.957664, 4.958471, 4.956212, 4.953946, 4.951943, 4.950333, 
    4.951114, 4.952014, 4.953312, 4.954513, 4.955637, 4.9566, 4.957409, 
    4.957942, 4.95862, 4.959163, 4.961884, 4.964809, 4.967964, 4.97138, 
    4.97507, 4.97903, 4.983232, 4.987618, 4.992094, 4.996525, 5.000741, 
    5.004525, 5.007628, 5.009777, 5.010693, 5.010121, 5.007853, 5.003766, 
    4.997855,
  // momentumY(26,42, 0-49)
    4.980917, 4.980814, 4.98041, 4.979715, 4.978751, 4.977537, 4.976097, 
    4.974453, 4.972636, 4.970678, 4.968611, 4.966472, 4.964302, 4.962132, 
    4.959999, 4.957001, 4.958748, 4.95652, 4.954246, 4.952245, 4.950657, 
    4.95166, 4.952818, 4.954448, 4.955894, 4.957162, 4.958123, 4.958803, 
    4.95908, 4.959553, 4.959918, 4.962606, 4.965451, 4.968475, 4.971704, 
    4.97515, 4.978807, 4.982642, 4.986598, 4.990582, 4.994461, 4.998068, 
    5.0012, 5.003619, 5.005074, 5.005314, 5.004117, 5.001315, 4.996832, 
    4.990704,
  // momentumY(26,43, 0-49)
    4.977679, 4.97776, 4.977554, 4.977072, 4.976327, 4.975336, 4.974116, 
    4.972692, 4.971086, 4.969328, 4.967451, 4.965489, 4.963478, 4.961449, 
    4.959437, 4.956493, 4.959065, 4.956875, 4.954607, 4.952624, 4.951071, 
    4.952264, 4.953651, 4.955585, 4.95726, 4.958661, 4.959623, 4.960185, 
    4.960233, 4.960534, 4.960759, 4.963408, 4.966163, 4.96904, 4.97206, 
    4.975228, 4.978531, 4.981936, 4.985381, 4.988777, 4.991995, 4.994875, 
    4.99723, 4.998845, 4.999496, 4.998971, 4.997089, 4.993732, 4.988872, 
    4.982594,
  // momentumY(26,44, 0-49)
    4.974301, 4.974561, 4.974557, 4.974297, 4.973784, 4.973035, 4.972059, 
    4.970877, 4.96951, 4.967981, 4.966322, 4.964559, 4.962726, 4.960854, 
    4.958971, 4.956134, 4.959414, 4.957269, 4.955017, 4.953065, 4.951551, 
    4.952901, 4.954484, 4.956686, 4.958561, 4.960083, 4.961043, 4.961501, 
    4.961351, 4.961507, 4.961627, 4.964231, 4.966889, 4.969604, 4.972392, 
    4.975247, 4.97815, 4.981063, 4.983919, 4.986634, 4.989085, 4.991127, 
    4.992589, 4.993289, 4.99304, 4.991673, 4.989062, 4.985146, 4.979949, 
    4.973607,
  // momentumY(26,45, 0-49)
    4.970855, 4.971286, 4.971483, 4.971446, 4.971176, 4.970679, 4.969965, 
    4.969045, 4.967938, 4.96666, 4.965239, 4.963696, 4.962062, 4.960358, 
    4.958611, 4.955917, 4.95979, 4.957693, 4.955468, 4.95355, 4.952076, 
    4.95355, 4.955291, 4.957713, 4.959756, 4.961379, 4.962333, 4.9627, 
    4.962382, 4.962423, 4.96246, 4.965011, 4.967559, 4.970098, 4.972632, 
    4.97514, 4.977598, 4.979958, 4.982154, 4.984101, 4.985687, 4.986785, 
    4.987253, 4.986942, 4.985713, 4.983451, 4.980091, 4.975633, 4.970161, 
    4.963855,
  // momentumY(26,46, 0-49)
    4.967414, 4.968003, 4.968394, 4.968578, 4.968554, 4.968318, 4.967876, 
    4.967232, 4.9664, 4.96539, 4.964222, 4.962915, 4.961491, 4.959968, 
    4.958365, 4.955836, 4.960183, 4.95814, 4.955951, 4.954069, 4.952631, 
    4.954192, 4.956049, 4.95864, 4.960809, 4.962502, 4.963447, 4.963733, 
    4.963276, 4.963221, 4.963187, 4.965672, 4.968098, 4.970442, 4.972695, 
    4.974825, 4.976792, 4.978544, 4.980013, 4.981115, 4.981754, 4.981822, 
    4.98121, 4.979815, 4.977552, 4.974366, 4.970264, 4.965308, 4.959643, 
    4.953489,
  // momentumY(26,47, 0-49)
    4.964046, 4.964777, 4.965352, 4.965752, 4.96597, 4.965997, 4.965829, 
    4.96547, 4.96492, 4.964187, 4.963284, 4.962223, 4.961019, 4.959685, 
    4.958235, 4.955878, 4.960584, 4.958601, 4.956454, 4.954607, 4.953197, 
    4.954808, 4.956738, 4.959435, 4.961684, 4.963416, 4.964339, 4.964552, 
    4.96398, 4.963842, 4.963738, 4.966136, 4.968418, 4.970546, 4.972489, 
    4.974205, 4.975642, 4.976735, 4.977419, 4.977613, 4.977237, 4.976211, 
    4.974462, 4.97194, 4.968619, 4.964515, 4.959707, 4.954324, 4.948567, 
    4.942689,
  // momentumY(26,48, 0-49)
    4.96081, 4.961668, 4.962411, 4.963017, 4.963469, 4.963753, 4.96386, 
    4.963782, 4.963516, 4.963064, 4.962431, 4.961621, 4.960644, 4.959507, 
    4.958216, 4.956029, 4.960979, 4.959066, 4.956965, 4.955151, 4.953761, 
    4.955386, 4.957339, 4.960083, 4.962356, 4.964089, 4.964973, 4.965117, 
    4.964446, 4.964223, 4.964039, 4.966322, 4.968429, 4.970309, 4.971912, 
    4.973177, 4.974042, 4.974437, 4.974288, 4.973528, 4.972093, 4.969935, 
    4.967025, 4.963368, 4.959004, 4.954024, 4.948578, 4.942863, 4.937129, 
    4.93166,
  // momentumY(26,49, 0-49)
    4.957191, 4.958059, 4.958873, 4.959602, 4.960219, 4.9607, 4.961027, 
    4.961179, 4.961144, 4.960912, 4.960473, 4.959821, 4.95895, 4.957851, 
    4.956515, 4.953525, 4.964903, 4.962058, 4.958658, 4.955644, 4.953284, 
    4.956749, 4.960586, 4.965696, 4.969499, 4.971891, 4.972278, 4.970906, 
    4.967642, 4.965106, 4.962541, 4.964893, 4.966942, 4.968615, 4.969858, 
    4.970594, 4.970757, 4.97027, 4.969067, 4.967099, 4.964337, 4.960783, 
    4.956475, 4.951499, 4.945994, 4.940145, 4.934196, 4.928425, 4.923135, 
    4.918625,
  // momentumY(27,0, 0-49)
    4.952485, 4.956017, 4.95919, 4.962013, 4.964487, 4.966623, 4.968421, 
    4.969888, 4.971034, 4.971874, 4.972427, 4.972726, 4.972806, 4.972714, 
    4.972504, 4.972033, 4.971988, 4.9717, 4.971503, 4.971475, 4.971662, 
    4.97227, 4.973104, 4.974205, 4.975557, 4.977133, 4.978898, 4.980816, 
    4.982846, 4.984953, 4.987058, 4.989343, 4.991569, 4.993695, 4.995677, 
    4.997463, 4.998989, 5.00017, 5.000906, 5.001068, 5.000506, 4.999043, 
    4.996487, 4.992639, 4.987311, 4.98035, 4.971671, 4.961278, 4.9493, 
    4.936006,
  // momentumY(27,1, 0-49)
    4.953785, 4.957267, 4.960383, 4.963142, 4.965549, 4.967614, 4.969344, 
    4.970743, 4.971827, 4.97261, 4.973116, 4.973373, 4.973421, 4.973308, 
    4.973083, 4.972408, 4.972571, 4.972211, 4.971914, 4.971784, 4.971873, 
    4.97256, 4.97343, 4.974563, 4.975933, 4.977504, 4.979235, 4.981091, 
    4.983034, 4.985042, 4.987011, 4.989357, 4.991658, 4.993884, 4.995999, 
    4.997962, 4.999713, 5.001177, 5.002253, 5.002817, 5.002716, 5.001765, 
    4.999763, 4.996496, 4.991755, 4.985361, 4.977194, 4.967225, 4.955546, 
    4.942395,
  // momentumY(27,2, 0-49)
    4.9551, 4.958522, 4.961576, 4.964267, 4.96661, 4.96861, 4.970279, 
    4.971625, 4.97266, 4.973405, 4.97388, 4.974118, 4.974155, 4.974039, 
    4.97382, 4.972966, 4.973311, 4.972891, 4.972506, 4.972278, 4.972264, 
    4.973009, 4.97389, 4.975019, 4.976368, 4.9779, 4.979566, 4.981339, 
    4.983176, 4.985064, 4.98687, 4.989237, 4.991573, 4.993855, 4.996058, 
    4.998144, 5.000066, 5.00175, 5.003102, 5.003998, 5.004288, 5.003786, 
    5.002285, 4.999563, 4.995397, 4.989588, 4.981988, 4.972539, 4.961292, 
    4.948447,
  // momentumY(27,3, 0-49)
    4.956424, 4.959782, 4.962767, 4.965392, 4.967669, 4.969612, 4.971227, 
    4.972527, 4.973528, 4.974247, 4.97471, 4.974946, 4.974991, 4.974892, 
    4.974695, 4.973688, 4.974173, 4.973708, 4.973245, 4.972928, 4.972816, 
    4.973597, 4.974463, 4.975552, 4.976844, 4.978302, 4.979884, 4.981561, 
    4.983288, 4.985043, 4.986671, 4.989024, 4.991359, 4.993658, 4.995905, 
    4.99807, 5.000108, 5.001954, 5.003517, 5.004678, 5.00529, 5.005171, 
    5.004114, 5.001892, 4.998278, 4.993056, 4.986063, 4.977203, 4.966496, 
    4.9541,
  // momentumY(27,4, 0-49)
    4.957763, 4.961049, 4.963962, 4.966518, 4.968731, 4.970614, 4.97218, 
    4.973444, 4.974419, 4.975125, 4.975588, 4.975837, 4.975906, 4.975838, 
    4.975676, 4.974549, 4.975114, 4.974617, 4.974098, 4.973704, 4.973499, 
    4.974296, 4.97512, 4.976135, 4.977338, 4.978698, 4.980179, 4.981754, 
    4.983374, 4.984993, 4.986437, 4.988748, 4.991049, 4.993332, 4.995584, 
    4.997785, 4.999891, 5.001845, 5.003561, 5.004924, 5.005792, 5.005991, 
    5.00532, 5.003553, 5.000459, 4.995819, 4.98945, 4.981233, 4.971154, 
    4.959323,
  // momentumY(27,5, 0-49)
    4.959124, 4.96233, 4.965165, 4.967649, 4.969796, 4.971621, 4.973139, 
    4.974367, 4.975321, 4.976024, 4.976496, 4.976768, 4.976871, 4.976844, 
    4.976726, 4.975518, 4.976087, 4.975574, 4.975018, 4.974565, 4.97428, 
    4.975071, 4.975831, 4.976738, 4.977826, 4.979064, 4.980437, 4.981911, 
    4.983433, 4.984925, 4.986189, 4.988428, 4.990667, 4.992902, 4.995128, 
    4.997325, 4.999457, 5.001471, 5.003284, 5.004794, 5.005862, 5.006324, 
    5.005984, 5.004626, 5.002022, 4.997947, 4.992211, 4.984674, 4.975287, 
    4.964118,
  // momentumY(27,6, 0-49)
    4.960515, 4.963633, 4.966385, 4.96879, 4.970866, 4.972629, 4.974098, 
    4.975291, 4.976225, 4.976924, 4.97741, 4.977711, 4.977855, 4.977876, 
    4.977808, 4.976558, 4.977046, 4.976531, 4.97596, 4.975471, 4.975124, 
    4.975888, 4.976562, 4.977334, 4.978279, 4.979381, 4.980637, 4.982016, 
    4.983459, 4.984834, 4.985934, 4.988077, 4.990227, 4.992387, 4.994555, 
    4.996716, 4.998837, 5.000868, 5.002738, 5.004347, 5.005566, 5.006243, 
    5.006188, 5.005199, 5.003053, 4.999527, 4.994426, 4.987591, 4.978942, 
    4.968504,
  // momentumY(27,7, 0-49)
    4.961944, 4.964969, 4.96763, 4.969948, 4.971945, 4.97364, 4.975054, 
    4.976207, 4.977119, 4.977812, 4.978312, 4.978641, 4.978827, 4.978899, 
    4.97888, 4.977633, 4.977947, 4.977446, 4.976884, 4.976382, 4.975995, 
    4.976711, 4.97728, 4.977891, 4.978675, 4.97963, 4.980768, 4.982057, 
    4.98344, 4.984717, 4.985673, 4.987694, 4.989734, 4.991795, 4.99388, 
    4.995977, 4.998057, 5.000075, 5.001965, 5.003634, 5.004968, 5.005818, 
    5.006014, 5.00536, 5.003646, 5.000652, 4.996178, 4.990054, 4.982172, 
    4.972516,
  // momentumY(27,8, 0-49)
    4.96342, 4.966343, 4.968904, 4.971127, 4.973035, 4.974654, 4.976002, 
    4.977108, 4.977989, 4.978671, 4.979177, 4.979532, 4.979758, 4.979877, 
    4.979905, 4.978708, 4.978746, 4.978274, 4.97775, 4.977262, 4.976861, 
    4.977507, 4.977953, 4.978384, 4.978992, 4.979788, 4.980811, 4.982022, 
    4.983364, 4.984567, 4.985405, 4.987285, 4.989192, 4.991133, 4.993113, 
    4.995123, 4.997139, 4.999117, 5.001001, 5.002707, 5.004125, 5.005124, 
    5.005543, 5.005198, 5.003892, 5.001414, 4.997559, 4.992144, 4.985043, 
    4.976196,
  // momentumY(27,9, 0-49)
    4.964952, 4.967762, 4.970212, 4.972329, 4.974138, 4.975667, 4.976941, 
    4.977984, 4.978825, 4.979486, 4.97999, 4.980362, 4.98062, 4.980781, 
    4.980847, 4.979746, 4.979405, 4.97898, 4.978518, 4.978075, 4.977688, 
    4.978245, 4.978553, 4.978786, 4.97921, 4.979844, 4.980752, 4.981893, 
    4.983215, 4.984366, 4.985122, 4.98684, 4.988597, 4.990402, 4.992261, 
    4.994167, 4.9961, 4.998025, 4.999886, 5.001608, 5.003094, 5.004222, 
    5.004846, 5.004794, 5.003879, 5.001898, 4.998647, 4.993936, 4.987614, 
    4.979589,
  // momentumY(27,10, 0-49)
    4.966544, 4.969228, 4.971554, 4.973551, 4.975248, 4.976675, 4.977859, 
    4.97883, 4.979616, 4.980243, 4.980734, 4.981112, 4.98139, 4.981582, 
    4.981678, 4.980717, 4.979891, 4.979529, 4.979159, 4.978791, 4.978449, 
    4.978896, 4.979054, 4.97908, 4.979313, 4.979784, 4.980581, 4.981661, 
    4.982981, 4.984105, 4.984818, 4.986358, 4.987952, 4.989606, 4.991331, 
    4.993123, 4.994964, 4.996823, 4.998651, 5.000382, 5.001927, 5.003174, 
    5.003991, 5.00422, 5.003681, 5.002182, 4.999519, 4.995496, 4.989943, 
    4.982737,
  // momentumY(27,11, 0-49)
    4.968184, 4.970732, 4.972922, 4.974787, 4.976358, 4.97767, 4.978752, 
    4.979636, 4.980354, 4.980931, 4.981393, 4.981763, 4.982052, 4.982261, 
    4.982378, 4.981594, 4.980174, 4.979899, 4.979648, 4.979387, 4.979123, 
    4.979436, 4.979437, 4.979248, 4.979291, 4.979603, 4.980292, 4.981318, 
    4.98265, 4.983774, 4.984485, 4.985836, 4.987253, 4.988749, 4.990333, 
    4.992004, 4.993749, 4.995539, 4.997333, 4.99907, 5.000671, 5.002034, 
    5.00304, 5.00354, 5.003365, 5.00233, 5.000237, 4.996881, 4.992076, 
    4.985673,
  // momentumY(27,12, 0-49)
    4.969869, 4.972264, 4.974305, 4.976025, 4.977458, 4.978641, 4.979606, 
    4.98039, 4.981024, 4.981538, 4.981959, 4.982306, 4.982589, 4.982803, 
    4.982933, 4.982355, 4.980234, 4.98007, 4.979968, 4.979845, 4.979689, 
    4.97985, 4.979685, 4.979283, 4.979139, 4.979298, 4.979885, 4.980863, 
    4.982218, 4.983363, 4.984119, 4.985269, 4.986504, 4.987836, 4.989278, 
    4.990828, 4.992476, 4.9942, 4.995962, 4.997709, 4.999368, 5.000849, 
    5.002039, 5.002804, 5.002984, 5.002398, 5.00085, 4.998134, 4.99405, 
    4.988423,
  // momentumY(27,13, 0-49)
    4.971578, 4.973805, 4.975684, 4.977247, 4.978529, 4.979571, 4.980408, 
    4.98108, 4.981618, 4.982056, 4.982419, 4.982728, 4.982991, 4.983199, 
    4.983337, 4.982982, 4.980053, 4.980028, 4.980104, 4.980148, 4.980134, 
    4.980123, 4.97979, 4.979178, 4.978858, 4.978872, 4.979362, 4.980295, 
    4.981681, 4.982868, 4.983716, 4.984661, 4.98571, 4.986878, 4.988178, 
    4.989611, 4.991169, 4.992833, 4.994571, 4.996334, 4.998056, 4.999658, 
    5.001034, 5.002057, 5.002578, 5.002422, 5.001395, 4.999288, 4.995888, 
    4.991003,
  // momentumY(27,14, 0-49)
    4.973285, 4.975332, 4.977035, 4.978428, 4.979551, 4.980443, 4.981143, 
    4.981692, 4.982125, 4.982474, 4.982768, 4.983025, 4.983253, 4.983449, 
    4.983591, 4.983465, 4.979623, 4.979764, 4.980047, 4.980291, 4.980448, 
    4.980245, 4.979743, 4.978934, 4.978452, 4.978334, 4.978735, 4.979624, 
    4.981044, 4.98229, 4.983274, 4.984014, 4.98488, 4.985888, 4.987052, 
    4.988374, 4.98985, 4.991462, 4.993183, 4.994971, 4.996765, 4.998491, 
    5.000052, 5.001328, 5.002178, 5.002431, 5.001897, 5.000363, 4.99761, 
    4.993423,
  // momentumY(27,15, 0-49)
    4.974969, 4.976818, 4.97833, 4.979544, 4.980499, 4.981234, 4.981791, 
    4.982209, 4.982529, 4.98278, 4.982994, 4.983189, 4.983375, 4.983549, 
    4.983696, 4.983794, 4.978942, 4.979278, 4.979795, 4.980265, 4.98062, 
    4.980211, 4.979545, 4.978554, 4.977929, 4.977694, 4.978014, 4.978863, 
    4.980318, 4.981638, 4.982798, 4.983336, 4.984023, 4.984879, 4.985915, 
    4.987135, 4.988539, 4.990111, 4.991827, 4.993648, 4.99552, 4.997373, 
    4.999117, 5.000638, 5.001802, 5.002442, 5.002368, 5.00137, 4.999219, 
    4.995688,
  // momentumY(27,16, 0-49)
    4.9766, 4.978232, 4.979541, 4.980565, 4.981343, 4.981917, 4.982327, 
    4.982615, 4.982817, 4.982967, 4.983095, 4.98322, 4.983356, 4.983504, 
    4.983661, 4.983968, 4.978021, 4.978576, 4.979346, 4.980065, 4.980643, 
    4.980015, 4.979194, 4.97804, 4.977294, 4.976964, 4.977215, 4.978029, 
    4.979517, 4.980919, 4.982292, 4.982636, 4.983153, 4.983865, 4.984783, 
    4.985914, 4.987255, 4.988797, 4.990517, 4.992379, 4.994334, 4.996316, 
    4.99824, 4.999999, 5.001459, 5.002461, 5.002818, 5.002316, 5.000722, 
    4.997799,
  // momentumY(27,17, 0-49)
    4.97815, 4.979545, 4.980634, 4.981458, 4.982053, 4.982463, 4.982728, 
    4.982884, 4.982973, 4.983024, 4.983063, 4.983118, 4.983199, 4.983321, 
    4.983489, 4.983988, 4.976887, 4.977677, 4.978717, 4.979698, 4.980515, 
    4.97966, 4.978692, 4.977397, 4.976559, 4.976156, 4.976355, 4.977139, 
    4.97866, 4.980151, 4.981763, 4.981924, 4.982281, 4.982859, 4.983669, 
    4.98472, 4.986009, 4.987531, 4.989263, 4.991172, 4.993215, 4.995326, 
    4.997425, 4.999409, 5.001151, 5.00249, 5.003245, 5.0032, 5.002119, 
    4.999754,
  // momentumY(27,18, 0-49)
    4.979592, 4.980724, 4.981576, 4.982186, 4.982595, 4.982841, 4.982964, 
    4.983, 4.982983, 4.982941, 4.9829, 4.982886, 4.982915, 4.983007, 
    4.983186, 4.983865, 4.975588, 4.976619, 4.977927, 4.979177, 4.980241, 
    4.979152, 4.978045, 4.976635, 4.97573, 4.975284, 4.975449, 4.976212, 
    4.977769, 4.979352, 4.981221, 4.981211, 4.981418, 4.981871, 4.982583, 
    4.983562, 4.984807, 4.986314, 4.988064, 4.990025, 4.992156, 4.994394, 
    4.996664, 4.998864, 5.000867, 5.002522, 5.003644, 5.004018, 5.003407, 
    5.001557,
  // momentumY(27,19, 0-49)
    4.980903, 4.98174, 4.98233, 4.982714, 4.982932, 4.983019, 4.98301, 
    4.982938, 4.982831, 4.982711, 4.982603, 4.982526, 4.982506, 4.982572, 
    4.982763, 4.983617, 4.9742, 4.975467, 4.977031, 4.978539, 4.979841, 
    4.978513, 4.97728, 4.975773, 4.974828, 4.974364, 4.974518, 4.975278, 
    4.976873, 4.978549, 4.980679, 4.98051, 4.980577, 4.980914, 4.981531, 
    4.982439, 4.983643, 4.985138, 4.986907, 4.988921, 4.991139, 4.993503, 
    4.995936, 4.998341, 5.000593, 5.002542, 5.004004, 5.004765, 5.004586, 
    5.00321,
  // momentumY(27,20, 0-49)
    4.982862, 4.984146, 4.985185, 4.986007, 4.98664, 4.987111, 4.987448, 
    4.987677, 4.987826, 4.987921, 4.987986, 4.988048, 4.988135, 4.988278, 
    4.988526, 0, 4.972143, 4.973258, 4.97473, 4.976183, 4.977445, 4.975578, 
    4.973876, 4.971932, 4.970649, 4.969963, 4.970038, 4.970872, 4.97272, 
    4.974809, 4.977582, 4.977671, 4.978006, 4.978611, 4.979485, 4.980634, 
    4.982059, 4.983755, 4.985709, 4.987898, 4.990287, 4.992825, 4.995441, 
    4.998047, 5.000524, 5.002726, 5.004475, 5.005559, 5.005739, 5.004762,
  // momentumY(27,21, 0-49)
    4.984021, 4.985055, 4.985878, 4.986519, 4.987, 4.98735, 4.987592, 
    4.987746, 4.987836, 4.987881, 4.987903, 4.987926, 4.987977, 4.98809, 
    4.988317, 0, 4.96787, 4.969113, 4.970778, 4.972454, 4.973938, 4.971829, 
    4.970017, 4.96804, 4.966849, 4.966359, 4.966709, 4.967876, 4.970111, 
    4.97262, 4.975931, 4.976147, 4.976643, 4.977433, 4.978511, 4.979876, 
    4.981517, 4.983426, 4.985584, 4.987966, 4.990533, 4.993235, 4.996002, 
    4.998747, 5.001359, 5.003693, 5.005579, 5.006813, 5.007162, 5.006378,
  // momentumY(27,22, 0-49)
    4.9851, 4.985905, 4.986529, 4.987001, 4.987345, 4.987583, 4.987735, 
    4.987818, 4.987849, 4.987846, 4.987824, 4.987807, 4.987818, 4.987895, 
    4.988095, 0, 4.96427, 4.965615, 4.967438, 4.969296, 4.970961, 4.968601, 
    4.96665, 4.964593, 4.963428, 4.963049, 4.963583, 4.964988, 4.96751, 
    4.970334, 4.974064, 4.974349, 4.974948, 4.975873, 4.977114, 4.978661, 
    4.980502, 4.982621, 4.984995, 4.987593, 4.990371, 4.993275, 4.996236, 
    4.999167, 5.001956, 5.004463, 5.006518, 5.007926, 5.008459, 5.007876,
  // momentumY(27,23, 0-49)
    4.986108, 4.986693, 4.987132, 4.98745, 4.987665, 4.987799, 4.987868, 
    4.987884, 4.987857, 4.987806, 4.987741, 4.98768, 4.987649, 4.987686, 
    4.987846, 0, 4.961174, 4.962575, 4.964491, 4.966458, 4.968225, 4.965626, 
    4.963521, 4.961361, 4.960176, 4.959849, 4.960501, 4.962069, 4.964801, 
    4.96786, 4.971903, 4.972238, 4.972919, 4.973962, 4.97535, 4.977074, 
    4.979115, 4.981455, 4.984063, 4.986903, 4.989927, 4.993075, 4.996275, 
    4.999434, 5.00244, 5.005151, 5.007399, 5.008994, 5.009711, 5.00932,
  // momentumY(27,24, 0-49)
    4.987052, 4.987432, 4.987696, 4.987866, 4.987962, 4.987997, 4.987984, 
    4.987933, 4.987851, 4.98775, 4.987639, 4.987533, 4.987454, 4.987441, 
    4.987548, 0, 4.958886, 4.960289, 4.962229, 4.964231, 4.966028, 4.963264, 
    4.961052, 4.958817, 4.957613, 4.957313, 4.958032, 4.959703, 4.962571, 
    4.965787, 4.970043, 4.970445, 4.971216, 4.972371, 4.973891, 4.975769, 
    4.977979, 4.980506, 4.983313, 4.986362, 4.989601, 4.992966, 4.996381, 
    4.99975, 5.002959, 5.005866, 5.0083, 5.010072, 5.010966, 5.010753,
  // momentumY(27,25, 0-49)
    4.987951, 4.988135, 4.988231, 4.988259, 4.988237, 4.988174, 4.98808, 
    4.987959, 4.987818, 4.987662, 4.987497, 4.987339, 4.987206, 4.987133, 
    4.987175, 0, 4.957164, 4.958512, 4.960404, 4.962363, 4.964118, 4.961286, 
    4.959035, 4.956786, 4.955588, 4.955317, 4.956082, 4.957819, 4.960765, 
    4.964076, 4.968446, 4.968953, 4.969841, 4.971123, 4.972783, 4.974807, 
    4.977177, 4.979869, 4.98285, 4.986078, 4.989499, 4.993052, 4.996652, 
    5.000207, 5.003596, 5.006678, 5.009283, 5.011218, 5.01227, 5.012215,
  // momentumY(27,26, 0-49)
    4.988813, 4.988812, 4.98875, 4.988639, 4.9885, 4.988336, 4.988153, 
    4.987953, 4.987741, 4.987518, 4.98729, 4.987069, 4.986872, 4.986731, 
    4.986691, 0, 4.956017, 4.957257, 4.959034, 4.960871, 4.962512, 4.95972, 
    4.957509, 4.955312, 4.954154, 4.953917, 4.954714, 4.956479, 4.959447, 
    4.962788, 4.967175, 4.967828, 4.968863, 4.970294, 4.972103, 4.974275, 
    4.976792, 4.979629, 4.982756, 4.986129, 4.989699, 4.9934, 4.997152, 
    5.000857, 5.004397, 5.007628, 5.010381, 5.01246, 5.013651, 5.013734,
  // momentumY(27,27, 0-49)
    4.98965, 4.989479, 4.989264, 4.98902, 4.988759, 4.988484, 4.9882, 
    4.987906, 4.987603, 4.987295, 4.986986, 4.986688, 4.986415, 4.986197, 
    4.986067, 0, 4.955529, 4.956617, 4.958216, 4.959864, 4.961324, 4.958663, 
    4.956551, 4.954452, 4.95335, 4.953136, 4.95393, 4.955672, 4.958594, 
    4.961887, 4.966184, 4.967004, 4.968203, 4.969788, 4.971744, 4.974054, 
    4.976701, 4.979663, 4.98291, 4.986403, 4.990092, 4.993917, 4.997795, 
    5.001633, 5.005309, 5.008677, 5.011567, 5.013782, 5.015105, 5.01531,
  // momentumY(27,28, 0-49)
    4.990469, 4.990145, 4.989788, 4.989411, 4.989022, 4.988625, 4.988218, 
    4.987805, 4.987385, 4.986967, 4.986554, 4.98616, 4.985801, 4.9855, 
    4.985283, 0, 4.956028, 4.956934, 4.958307, 4.959707, 4.96093, 4.958463, 
    4.956476, 4.954484, 4.953412, 4.953169, 4.953884, 4.955516, 4.958292, 
    4.961439, 4.965523, 4.966502, 4.967848, 4.969568, 4.971642, 4.974057, 
    4.976798, 4.979848, 4.983181, 4.986762, 4.990545, 4.994473, 4.998466, 
    5.002428, 5.006239, 5.009749, 5.012783, 5.015139, 5.016596, 5.016923,
  // momentumY(27,29, 0-49)
    4.991272, 4.99082, 4.990334, 4.989828, 4.989304, 4.988763, 4.988209, 
    4.987643, 4.987072, 4.986504, 4.985958, 4.985448, 4.984994, 4.984619, 
    4.984338, 0, 4.957261, 4.957983, 4.959101, 4.960205, 4.96113, 4.958851, 
    4.956955, 4.955013, 4.953891, 4.953528, 4.954064, 4.955482, 4.958002, 
    4.960886, 4.964627, 4.965713, 4.967158, 4.968967, 4.971126, 4.973623, 
    4.976449, 4.979589, 4.983022, 4.986718, 4.990633, 4.994709, 4.998869, 
    5.003012, 5.00701, 5.010713, 5.013935, 5.016467, 5.018081, 5.018536,
  // momentumY(27,30, 0-49)
    4.991342, 4.990104, 4.98886, 4.987627, 4.986415, 4.985223, 4.984044, 
    4.982868, 4.981678, 4.980457, 4.979197, 4.977892, 4.976555, 4.975228, 
    4.973989, 4.972118, 4.961142, 4.961493, 4.962195, 4.962931, 4.963588, 
    4.961671, 4.96014, 4.958567, 4.957699, 4.957439, 4.957901, 4.95906, 
    4.961126, 4.963423, 4.966387, 4.96713, 4.968222, 4.969685, 4.971525, 
    4.973748, 4.976355, 4.979339, 4.982685, 4.986363, 4.990328, 4.994513, 
    4.998833, 5.003178, 5.007408, 5.011355, 5.014824, 5.017593, 5.019419, 
    5.020052,
  // momentumY(27,31, 0-49)
    4.992085, 4.990796, 4.989485, 4.988165, 4.986845, 4.985525, 4.9842, 
    4.982865, 4.981511, 4.980129, 4.978714, 4.977267, 4.975796, 4.974329, 
    4.972923, 4.971511, 4.96095, 4.960932, 4.961246, 4.961601, 4.961905, 
    4.960153, 4.958697, 4.957186, 4.956329, 4.956063, 4.956516, 4.957662, 
    4.959669, 4.961869, 4.964588, 4.965552, 4.966871, 4.968566, 4.970642, 
    4.973103, 4.975951, 4.979178, 4.982767, 4.986686, 4.990888, 4.995302, 
    4.99984, 5.004383, 5.008787, 5.012877, 5.016449, 5.019275, 5.021107, 
    5.021693,
  // momentumY(27,32, 0-49)
    4.992704, 4.991362, 4.989981, 4.988571, 4.987143, 4.985699, 4.984235, 
    4.982752, 4.981244, 4.979711, 4.978148, 4.976559, 4.974949, 4.97334, 
    4.971759, 4.970668, 4.96088, 4.960486, 4.96041, 4.960387, 4.96035, 
    4.958791, 4.957444, 4.956033, 4.955215, 4.954963, 4.95541, 4.956527, 
    4.958438, 4.960497, 4.962925, 4.964082, 4.965597, 4.967487, 4.969763, 
    4.972429, 4.975488, 4.97893, 4.982742, 4.986887, 4.991313, 4.995951, 
    5.000702, 5.005444, 5.010021, 5.014254, 5.017927, 5.020806, 5.022637, 
    5.023165,
  // momentumY(27,33, 0-49)
    4.993176, 4.991786, 4.990337, 4.988843, 4.987313, 4.98575, 4.984156, 
    4.982533, 4.980882, 4.979203, 4.977501, 4.975778, 4.97404, 4.972296, 
    4.97056, 4.969613, 4.960853, 4.960111, 4.959667, 4.95929, 4.95894, 
    4.957603, 4.956401, 4.955134, 4.954391, 4.954172, 4.954613, 4.955681, 
    4.957458, 4.959333, 4.961436, 4.962754, 4.964429, 4.966482, 4.968922, 
    4.971757, 4.974994, 4.978625, 4.982632, 4.986979, 4.991614, 4.996459, 
    5.001411, 5.006339, 5.011081, 5.015445, 5.019209, 5.022128, 5.023943, 
    5.024394,
  // momentumY(27,34, 0-49)
    4.993468, 4.992046, 4.990543, 4.988973, 4.98735, 4.985679, 4.983964, 
    4.982211, 4.980426, 4.978615, 4.976783, 4.974936, 4.973081, 4.971223, 
    4.96936, 4.968389, 4.960826, 4.959777, 4.958998, 4.958305, 4.957679, 
    4.956588, 4.955568, 4.954486, 4.953852, 4.953686, 4.95412, 4.955118, 
    4.956721, 4.958376, 4.960136, 4.961588, 4.963395, 4.965575, 4.968145, 
    4.971118, 4.974501, 4.978288, 4.98246, 4.986983, 4.9918, 4.996827, 
    5.001957, 5.00705, 5.011934, 5.016407, 5.020238, 5.023174, 5.024948, 
    5.025294,
  // momentumY(27,35, 0-49)
    4.993543, 4.992109, 4.990572, 4.988945, 4.987246, 4.98548, 4.983659, 
    4.98179, 4.979885, 4.977952, 4.976004, 4.97405, 4.972095, 4.970143, 
    4.968186, 4.967057, 4.960784, 4.959477, 4.958406, 4.957438, 4.956577, 
    4.955748, 4.954938, 4.954085, 4.953589, 4.953495, 4.953919, 4.954828, 
    4.956221, 4.957632, 4.959045, 4.960607, 4.962515, 4.964794, 4.967463, 
    4.970541, 4.974034, 4.977944, 4.982249, 4.986913, 4.991876, 4.997052, 
    5.002326, 5.007547, 5.012538, 5.017087, 5.020951, 5.023866, 5.025561, 
    5.025771,
  // momentumY(27,36, 0-49)
    4.993363, 4.991943, 4.990395, 4.988733, 4.986978, 4.985139, 4.983231, 
    4.981265, 4.979257, 4.977222, 4.975175, 4.973129, 4.971095, 4.969073, 
    4.967054, 4.965679, 4.960728, 4.959213, 4.957893, 4.956695, 4.95564, 
    4.955082, 4.954507, 4.953914, 4.953588, 4.953581, 4.953995, 4.954797, 
    4.955952, 4.957104, 4.958177, 4.959828, 4.961814, 4.964163, 4.966903, 
    4.970053, 4.973625, 4.977619, 4.982017, 4.986782, 4.991848, 4.997127, 
    5.002496, 5.007801, 5.012851, 5.017424, 5.021269, 5.024117, 5.025689, 
    5.025723,
  // momentumY(27,37, 0-49)
    4.992894, 4.991515, 4.989983, 4.988314, 4.986529, 4.984643, 4.982672, 
    4.980633, 4.978547, 4.97643, 4.974305, 4.972188, 4.970094, 4.968026, 
    4.965975, 4.964311, 4.960664, 4.958989, 4.957465, 4.956078, 4.95487, 
    4.954582, 4.954257, 4.953956, 4.953823, 4.953918, 4.954322, 4.955003, 
    4.955902, 4.956789, 4.957542, 4.959267, 4.961312, 4.963708, 4.96649, 
    4.969682, 4.973296, 4.977336, 4.981783, 4.986598, 4.991717, 4.997042, 
    5.00245, 5.007774, 5.01282, 5.017355, 5.021121, 5.02384, 5.025236, 
    5.025045,
  // momentumY(27,38, 0-49)
    4.992102, 4.990796, 4.989309, 4.987664, 4.985879, 4.983975, 4.981972, 
    4.979889, 4.977752, 4.97558, 4.973402, 4.971236, 4.969102, 4.967009, 
    4.964951, 4.962999, 4.960605, 4.958811, 4.957121, 4.955583, 4.954257, 
    4.954235, 4.954173, 4.954182, 4.954263, 4.954476, 4.954871, 4.955422, 
    4.956054, 4.956684, 4.957149, 4.958934, 4.961021, 4.963445, 4.966245, 
    4.969447, 4.97307, 4.977113, 4.981561, 4.986373, 4.991481, 4.996788, 
    5.002161, 5.007431, 5.012395, 5.016815, 5.020426, 5.022949, 5.024106, 
    5.023642,
  // momentumY(27,39, 0-49)
    4.990971, 4.989764, 4.988355, 4.986764, 4.985014, 4.983126, 4.981123, 
    4.97903, 4.976871, 4.974676, 4.97247, 4.970282, 4.968132, 4.966033, 
    4.963985, 4.961775, 4.960558, 4.95868, 4.956858, 4.955204, 4.953793, 
    4.954025, 4.954226, 4.954561, 4.954874, 4.955217, 4.955606, 4.956029, 
    4.956393, 4.956779, 4.956996, 4.958832, 4.960948, 4.963384, 4.966179, 
    4.969365, 4.972958, 4.976961, 4.981358, 4.986107, 4.991138, 4.99635, 
    5.001607, 5.006737, 5.011529, 5.015744, 5.019113, 5.021358, 5.022209, 
    5.021421,
  // momentumY(27,40, 0-49)
    4.989492, 4.988411, 4.987108, 4.985605, 4.983923, 4.982087, 4.980121, 
    4.978053, 4.975909, 4.973721, 4.971519, 4.969333, 4.96719, 4.965103, 
    4.963079, 4.960662, 4.960529, 4.958594, 4.956668, 4.954926, 4.953461, 
    4.953931, 4.954395, 4.955062, 4.955615, 4.956097, 4.956487, 4.956788, 
    4.956896, 4.957064, 4.957074, 4.958955, 4.961094, 4.963527, 4.966299, 
    4.96944, 4.972969, 4.976889, 4.98118, 4.9858, 4.990678, 4.995711, 
    5.000761, 5.005651, 5.010171, 5.01408, 5.017112, 5.018996, 5.019468, 
    5.018303,
  // momentumY(27,41, 0-49)
    4.98767, 4.986738, 4.98557, 4.984185, 4.982606, 4.98086, 4.978968, 
    4.97696, 4.974867, 4.972721, 4.970555, 4.9684, 4.966283, 4.964226, 
    4.962235, 4.959669, 4.96052, 4.958544, 4.956538, 4.954738, 4.95324, 
    4.953933, 4.95465, 4.955646, 4.956444, 4.957076, 4.957476, 4.957663, 
    4.957536, 4.957518, 4.957366, 4.959292, 4.961448, 4.963868, 4.9666, 
    4.969671, 4.973102, 4.976892, 4.98102, 4.985444, 4.99009, 4.994852, 
    4.999594, 5.004138, 5.008276, 5.01177, 5.014363, 5.015793, 5.015814, 
    5.014226,
  // momentumY(27,42, 0-49)
    4.985522, 4.98476, 4.983753, 4.982516, 4.981074, 4.97945, 4.977669, 
    4.975759, 4.973754, 4.971684, 4.969582, 4.967484, 4.965418, 4.963405, 
    4.961457, 4.958804, 4.960528, 4.958524, 4.956461, 4.954623, 4.953115, 
    4.954007, 4.954963, 4.956277, 4.957321, 4.958108, 4.958529, 4.958621, 
    4.958286, 4.958118, 4.957849, 4.959821, 4.961989, 4.96439, 4.967066, 
    4.970046, 4.973344, 4.976959, 4.980868, 4.985023, 4.989351, 4.993749, 
    4.998077, 5.002162, 5.005802, 5.008768, 5.010814, 5.011698, 5.011199, 
    5.009146,
  // momentumY(27,43, 0-49)
    4.983078, 4.982504, 4.981679, 4.980618, 4.979343, 4.977874, 4.976239, 
    4.974464, 4.972579, 4.970617, 4.968614, 4.966598, 4.964602, 4.962647, 
    4.96075, 4.958064, 4.960546, 4.958526, 4.956423, 4.954565, 4.953062, 
    4.954131, 4.955307, 4.956923, 4.958204, 4.959147, 4.959601, 4.959621, 
    4.959113, 4.958833, 4.958492, 4.960511, 4.962692, 4.965067, 4.967675, 
    4.97054, 4.973672, 4.977067, 4.980697, 4.984512, 4.988438, 4.992373, 
    4.996177, 4.999687, 5.00271, 5.00503, 5.006423, 5.006673, 5.005592, 
    5.003043,
  // momentumY(27,44, 0-49)
    4.980382, 4.980007, 4.979383, 4.978521, 4.97744, 4.976157, 4.974699, 
    4.973089, 4.971357, 4.969535, 4.967654, 4.965747, 4.963842, 4.961959, 
    4.960116, 4.957444, 4.96057, 4.958542, 4.956412, 4.954548, 4.953062, 
    4.954283, 4.955656, 4.957548, 4.959053, 4.960151, 4.960651, 4.960621, 
    4.959981, 4.95963, 4.959256, 4.961325, 4.963518, 4.965861, 4.968388, 
    4.971116, 4.974051, 4.97718, 4.980473, 4.983876, 4.987314, 4.990685, 
    4.993859, 4.996679, 4.998967, 5.000529, 5.001168, 5.000703, 4.998985, 
    4.995923,
  // momentumY(27,45, 0-49)
    4.977487, 4.977318, 4.976908, 4.976263, 4.975397, 4.974328, 4.973073, 
    4.971658, 4.970108, 4.968452, 4.96672, 4.964941, 4.963143, 4.961346, 
    4.959565, 4.956938, 4.960594, 4.958564, 4.956421, 4.954561, 4.953098, 
    4.954445, 4.955987, 4.958123, 4.959834, 4.961078, 4.961632, 4.961581, 
    4.960852, 4.960466, 4.960093, 4.962214, 4.964419, 4.966725, 4.969159, 
    4.971728, 4.974432, 4.977252, 4.980149, 4.983069, 4.985935, 4.988648, 
    4.991086, 4.993104, 4.994545, 4.995243, 4.995037, 4.993789, 4.991396, 
    4.987819,
  // momentumY(27,46, 0-49)
    4.974452, 4.974493, 4.974304, 4.97389, 4.973258, 4.972421, 4.971393, 
    4.970196, 4.968852, 4.967385, 4.965823, 4.964191, 4.962515, 4.960814, 
    4.959103, 4.956544, 4.960613, 4.958589, 4.956441, 4.954591, 4.953156, 
    4.954598, 4.956281, 4.95862, 4.960506, 4.961886, 4.962506, 4.96246, 
    4.961684, 4.961299, 4.960954, 4.963126, 4.965339, 4.9676, 4.969926, 
    4.972314, 4.974755, 4.97722, 4.979667, 4.982036, 4.98425, 4.986214, 
    4.987817, 4.988932, 4.989427, 4.989168, 4.988042, 4.98596, 4.982873, 
    4.9788,
  // momentumY(27,47, 0-49)
    4.971342, 4.971589, 4.971627, 4.971451, 4.971065, 4.970476, 4.969693, 
    4.968733, 4.967612, 4.966353, 4.964977, 4.963507, 4.961967, 4.960371, 
    4.958735, 4.956259, 4.960622, 4.95861, 4.956469, 4.954632, 4.953219, 
    4.954731, 4.956517, 4.959014, 4.961045, 4.962544, 4.963233, 4.963216, 
    4.962434, 4.962078, 4.961781, 4.963998, 4.966213, 4.96842, 4.970622, 
    4.972805, 4.974948, 4.977016, 4.978959, 4.98071, 4.982198, 4.983331, 
    4.98401, 4.984134, 4.9836, 4.982316, 4.980217, 4.977271, 4.973495, 
    4.968967,
  // momentumY(27,48, 0-49)
    4.968221, 4.96867, 4.968932, 4.968997, 4.968864, 4.968532, 4.968005, 
    4.967294, 4.966412, 4.965373, 4.964195, 4.962899, 4.961504, 4.960023, 
    4.958469, 4.956077, 4.960622, 4.958631, 4.9565, 4.954679, 4.953285, 
    4.954834, 4.956685, 4.959286, 4.961421, 4.963017, 4.963776, 4.963808, 
    4.963056, 4.96275, 4.962512, 4.964767, 4.96697, 4.969106, 4.971163, 
    4.973114, 4.974928, 4.976556, 4.977943, 4.97902, 4.979716, 4.979949, 
    4.979635, 4.978698, 4.977073, 4.974717, 4.971618, 4.96781, 4.963374, 
    4.958452,
  // momentumY(27,49, 0-49)
    4.964688, 4.965261, 4.965686, 4.965944, 4.966022, 4.965912, 4.965609, 
    4.96511, 4.964419, 4.963542, 4.962485, 4.96126, 4.959875, 4.958338, 
    4.95665, 4.953324, 4.963948, 4.960972, 4.957505, 4.954463, 4.952101, 
    4.95546, 4.959188, 4.964164, 4.967905, 4.970287, 4.97073, 4.969472, 
    4.966397, 4.964046, 4.961688, 4.964251, 4.966651, 4.968855, 4.970845, 
    4.972581, 4.974022, 4.975112, 4.975787, 4.975982, 4.975631, 4.974669, 
    4.973047, 4.97073, 4.967712, 4.964019, 4.959729, 4.954966, 4.949904, 
    4.944765,
  // momentumY(28,0, 0-49)
    4.963037, 4.965694, 4.96799, 4.96993, 4.971521, 4.972774, 4.973701, 
    4.974322, 4.97466, 4.974749, 4.974625, 4.974331, 4.973917, 4.973434, 
    4.972936, 4.972286, 4.972091, 4.971761, 4.971567, 4.971555, 4.971744, 
    4.972298, 4.973012, 4.97391, 4.974973, 4.97617, 4.977477, 4.978871, 
    4.980332, 4.981852, 4.983389, 4.985156, 4.986973, 4.988846, 4.990781, 
    4.992773, 4.99481, 4.99686, 4.998869, 5.000762, 5.002431, 5.003738, 
    5.00451, 5.00454, 5.003603, 5.00145, 4.997844, 4.992567, 4.985462, 
    4.976461,
  // momentumY(28,1, 0-49)
    4.964329, 4.966931, 4.969166, 4.971049, 4.972588, 4.973791, 4.974676, 
    4.975263, 4.975576, 4.975647, 4.975512, 4.975218, 4.974807, 4.97433, 
    4.973841, 4.973016, 4.97299, 4.972588, 4.972288, 4.972158, 4.972225, 
    4.97281, 4.973512, 4.974387, 4.975416, 4.976565, 4.977803, 4.979111, 
    4.980468, 4.981872, 4.983257, 4.985047, 4.986896, 4.988817, 4.990819, 
    4.992906, 4.995065, 4.997271, 4.999474, 5.001599, 5.003541, 5.005161, 
    5.006287, 5.006708, 5.006192, 5.004486, 5.001334, 4.996506, 4.989824, 
    4.981192,
  // momentumY(28,2, 0-49)
    4.965621, 4.968162, 4.970339, 4.972167, 4.973656, 4.974818, 4.975669, 
    4.976233, 4.976532, 4.976597, 4.976467, 4.976181, 4.975784, 4.975326, 
    4.974851, 4.973862, 4.973973, 4.973501, 4.973098, 4.972849, 4.972789, 
    4.973388, 4.974058, 4.974888, 4.97586, 4.976943, 4.978105, 4.979328, 
    4.98059, 4.981882, 4.983115, 4.984918, 4.986787, 4.988737, 4.990783, 
    4.992933, 4.995179, 4.997493, 4.999833, 5.002124, 5.004266, 5.00612, 
    5.007517, 5.00825, 5.008084, 5.006764, 5.004031, 4.999646, 4.993412, 
    4.985214,
  // momentumY(28,3, 0-49)
    4.966917, 4.969394, 4.971512, 4.973285, 4.974725, 4.975849, 4.976673, 
    4.977219, 4.97751, 4.977582, 4.977464, 4.977196, 4.976823, 4.976389, 
    4.975935, 4.974799, 4.974998, 4.974462, 4.973961, 4.973601, 4.973414, 
    4.97401, 4.974627, 4.975387, 4.976283, 4.977287, 4.978371, 4.979517, 
    4.980698, 4.981891, 4.98298, 4.984787, 4.986662, 4.988626, 4.990697, 
    4.992883, 4.995177, 4.997558, 4.999983, 5.002381, 5.004653, 5.00667, 
    5.008263, 5.009232, 5.009345, 5.008354, 5.006002, 5.002043, 4.996274, 
    4.988564,
  // momentumY(28,4, 0-49)
    4.968223, 4.970632, 4.972686, 4.974402, 4.975794, 4.97688, 4.977679, 
    4.97821, 4.978501, 4.97858, 4.978481, 4.97824, 4.977897, 4.977489, 
    4.97706, 4.975801, 4.976025, 4.975429, 4.974844, 4.97438, 4.974075, 
    4.974649, 4.975199, 4.975864, 4.976665, 4.977577, 4.978583, 4.979664, 
    4.980787, 4.981899, 4.982858, 4.984657, 4.986529, 4.988494, 4.99057, 
    4.992767, 4.99508, 4.997489, 4.999952, 5.002404, 5.004749, 5.006863, 
    5.008582, 5.00972, 5.010053, 5.009339, 5.007329, 5.00378, 4.998486, 
    4.991301,
  // momentumY(28,5, 0-49)
    4.969545, 4.971881, 4.973867, 4.975522, 4.976862, 4.977907, 4.978678, 
    4.979195, 4.979484, 4.979575, 4.979497, 4.979285, 4.978973, 4.978598, 
    4.978193, 4.976839, 4.977013, 4.976367, 4.975714, 4.975161, 4.97475, 
    4.975285, 4.975749, 4.976297, 4.976986, 4.977798, 4.978731, 4.979761, 
    4.980849, 4.981899, 4.982753, 4.984535, 4.986391, 4.988342, 4.990406, 
    4.992593, 4.994897, 4.997301, 4.999764, 5.002223, 5.00459, 5.006744, 
    5.008537, 5.009789, 5.010285, 5.009804, 5.008102, 5.004949, 5.000133, 
    4.993503,
  // momentumY(28,6, 0-49)
    4.970886, 4.97314, 4.975051, 4.976639, 4.977922, 4.978922, 4.979661, 
    4.98016, 4.980445, 4.980545, 4.980488, 4.980305, 4.980027, 4.979684, 
    4.979302, 4.977885, 4.977926, 4.977243, 4.97654, 4.975917, 4.975418, 
    4.975897, 4.97626, 4.976669, 4.977231, 4.977938, 4.978801, 4.979794, 
    4.980872, 4.981885, 4.982657, 4.984412, 4.986242, 4.988164, 4.990201, 
    4.992358, 4.994633, 4.997004, 4.999434, 5.001863, 5.00421, 5.006363, 
    5.008183, 5.0095, 5.010123, 5.009836, 5.008419, 5.005644, 5.001309, 
    4.995253,
  // momentumY(28,7, 0-49)
    4.97225, 4.974414, 4.976242, 4.977755, 4.978972, 4.979918, 4.980618, 
    4.981094, 4.98137, 4.981475, 4.981435, 4.981279, 4.981033, 4.980721, 
    4.98036, 4.978918, 4.978734, 4.978028, 4.977297, 4.976627, 4.976062, 
    4.976467, 4.976714, 4.976967, 4.977389, 4.977985, 4.978783, 4.979753, 
    4.980847, 4.981849, 4.982569, 4.984282, 4.986072, 4.987955, 4.989949, 
    4.992061, 4.994284, 4.996599, 4.998971, 5.001343, 5.003639, 5.005757, 
    5.007569, 5.008923, 5.00964, 5.009525, 5.00837, 5.005964, 5.002109, 
    4.996638,
  // momentumY(28,8, 0-49)
    4.973632, 4.975698, 4.977432, 4.978859, 4.980003, 4.980888, 4.981541, 
    4.981984, 4.982244, 4.982347, 4.98232, 4.982186, 4.981969, 4.981684, 
    4.98134, 4.979915, 4.979413, 4.978697, 4.977963, 4.977275, 4.97667, 
    4.976981, 4.977097, 4.97718, 4.977454, 4.977934, 4.978669, 4.97963, 
    4.980763, 4.981778, 4.982479, 4.984136, 4.985872, 4.987704, 4.989642, 
    4.991693, 4.99385, 4.996092, 4.998385, 5.00068, 5.002903, 5.004966, 
    5.006748, 5.008116, 5.00891, 5.00895, 5.008045, 5.005998, 5.00262, 
    4.997739,
  // momentumY(28,9, 0-49)
    4.975026, 4.976983, 4.978614, 4.979947, 4.981006, 4.98182, 4.982415, 
    4.982818, 4.983053, 4.983148, 4.983126, 4.983008, 4.982814, 4.982553, 
    4.982228, 4.980858, 4.979939, 4.979236, 4.978528, 4.977848, 4.977229, 
    4.97743, 4.977406, 4.977305, 4.977422, 4.977784, 4.978463, 4.979421, 
    4.980612, 4.981666, 4.98238, 4.983967, 4.985638, 4.987401, 4.989273, 
    4.991251, 4.993327, 4.995483, 4.997686, 4.999889, 5.002028, 5.004021, 
    5.005765, 5.007137, 5.007996, 5.008182, 5.00752, 5.005828, 5.002922, 
    4.998632,
  // momentumY(28,10, 0-49)
    4.976417, 4.978255, 4.979773, 4.981001, 4.981967, 4.9827, 4.98323, 
    4.983584, 4.983787, 4.983865, 4.98384, 4.983733, 4.983557, 4.983315, 
    4.983003, 4.981734, 4.980297, 4.979631, 4.978978, 4.97834, 4.977737, 
    4.977809, 4.977633, 4.977343, 4.9773, 4.977544, 4.978166, 4.979129, 
    4.980392, 4.981504, 4.982268, 4.983768, 4.985357, 4.987044, 4.988835, 
    4.990729, 4.992716, 4.994777, 4.996881, 4.998987, 5.001035, 5.002955, 
    5.004656, 5.00603, 5.006954, 5.007286, 5.006864, 5.005523, 5.003084, 
    4.999376,
  // momentumY(28,11, 0-49)
    4.977788, 4.979498, 4.980894, 4.982008, 4.982872, 4.983517, 4.983973, 
    4.984268, 4.984429, 4.984483, 4.984451, 4.984347, 4.984181, 4.983957, 
    4.983658, 4.98253, 4.980477, 4.979874, 4.979309, 4.978745, 4.978193, 
    4.978118, 4.977784, 4.977296, 4.977094, 4.977222, 4.97779, 4.978761, 
    4.980103, 4.981291, 4.982141, 4.983537, 4.985031, 4.986626, 4.988327, 
    4.990128, 4.992017, 4.993978, 4.995981, 4.997988, 4.999948, 5.001796, 
    5.00346, 5.004842, 5.005836, 5.006314, 5.006134, 5.005139, 5.003159, 
    5.000023,
  // momentumY(28,12, 0-49)
    4.979121, 4.98069, 4.981956, 4.982948, 4.983704, 4.984252, 4.984627, 
    4.984859, 4.984973, 4.984995, 4.984945, 4.984837, 4.984681, 4.984471, 
    4.984189, 4.983234, 4.980469, 4.979962, 4.979518, 4.979064, 4.978595, 
    4.978358, 4.977861, 4.977178, 4.976821, 4.976835, 4.97735, 4.978325, 
    4.979751, 4.981029, 4.981995, 4.983273, 4.984656, 4.986147, 4.987747, 
    4.989446, 4.991234, 4.993092, 4.994994, 4.996906, 4.998783, 5.000571, 
    5.002206, 5.003607, 5.004677, 5.00531, 5.005374, 5.004723, 5.003193, 
    5.000611,
  // momentumY(28,13, 0-49)
    4.980392, 4.981812, 4.982938, 4.983803, 4.984443, 4.98489, 4.985179, 
    4.985341, 4.985403, 4.985387, 4.985314, 4.985199, 4.985044, 4.984848, 
    4.984589, 4.983837, 4.980271, 4.979891, 4.979608, 4.979298, 4.978949, 
    4.978534, 4.977874, 4.977001, 4.976495, 4.976401, 4.976861, 4.977839, 
    4.979345, 4.980719, 4.981833, 4.982975, 4.984235, 4.98561, 4.987098, 
    4.988689, 4.990372, 4.992128, 4.993932, 4.995756, 4.997561, 4.999301, 
    5.00092, 5.002353, 5.003514, 5.00431, 5.004621, 5.004309, 5.003215, 
    5.001168,
  // momentumY(28,14, 0-49)
    4.981575, 4.982839, 4.983819, 4.984552, 4.985072, 4.985415, 4.985616, 
    4.985703, 4.985707, 4.98565, 4.98555, 4.985421, 4.985268, 4.985085, 
    4.984856, 4.98433, 4.97988, 4.979667, 4.979576, 4.979448, 4.979251, 
    4.97865, 4.977829, 4.976778, 4.976137, 4.975942, 4.976348, 4.97732, 
    4.978895, 4.98037, 4.981659, 4.982649, 4.98377, 4.985018, 4.986386, 
    4.987864, 4.989438, 4.991094, 4.992805, 4.99455, 4.996294, 4.998002, 
    4.999622, 5.001102, 5.002368, 5.003336, 5.003896, 5.003918, 5.003249, 
    5.001713,
  // momentumY(28,15, 0-49)
    4.982654, 4.983751, 4.984578, 4.985173, 4.985571, 4.985808, 4.985918, 
    4.98593, 4.985873, 4.985772, 4.985643, 4.985499, 4.985344, 4.985178, 
    4.984991, 4.984704, 4.979304, 4.979292, 4.979429, 4.979517, 4.979506, 
    4.978709, 4.977736, 4.976521, 4.975759, 4.975474, 4.975827, 4.976785, 
    4.978418, 4.979989, 4.981472, 4.982297, 4.983266, 4.984376, 4.985615, 
    4.986974, 4.988441, 4.989997, 4.991624, 4.993299, 4.994998, 4.996687, 
    4.998328, 4.999872, 5.001257, 5.002406, 5.003217, 5.003567, 5.003305, 
    5.002254,
  // momentumY(28,16, 0-49)
    4.983608, 4.984528, 4.985196, 4.98565, 4.985922, 4.986052, 4.98607, 
    4.986007, 4.98589, 4.985743, 4.985583, 4.985423, 4.985268, 4.985124, 
    4.984986, 4.984951, 4.978553, 4.978775, 4.979172, 4.979506, 4.979712, 
    4.978718, 4.977604, 4.976244, 4.975379, 4.975018, 4.975318, 4.976254, 
    4.977931, 4.979589, 4.981279, 4.981926, 4.98273, 4.983689, 4.984793, 
    4.986029, 4.987384, 4.988845, 4.990394, 4.992012, 4.993679, 4.995368, 
    4.997046, 4.998671, 5.000189, 5.001527, 5.002593, 5.003264, 5.003393, 
    5.002801,
  // momentumY(28,17, 0-49)
    4.984422, 4.985153, 4.985654, 4.985961, 4.986106, 4.986128, 4.986056, 
    4.985919, 4.985743, 4.985553, 4.985363, 4.985186, 4.985034, 4.984914, 
    4.984838, 4.985061, 4.977653, 4.978134, 4.978813, 4.97942, 4.979869, 
    4.978677, 4.977434, 4.975953, 4.975008, 4.974584, 4.974835, 4.975744, 
    4.977448, 4.979182, 4.981081, 4.981539, 4.982168, 4.982968, 4.983927, 
    4.985033, 4.986276, 4.987643, 4.98912, 4.990694, 4.992342, 4.994048, 
    4.995781, 4.997505, 4.999168, 5.000705, 5.002026, 5.00301, 5.003512, 
    5.003355,
  // momentumY(28,18, 0-49)
    4.985089, 4.985617, 4.985938, 4.98609, 4.986105, 4.986018, 4.985858, 
    4.985652, 4.985424, 4.985193, 4.984977, 4.984787, 4.98464, 4.984551, 
    4.984545, 4.985033, 4.976648, 4.977406, 4.978383, 4.979276, 4.979985, 
    4.978594, 4.977239, 4.975657, 4.97465, 4.974179, 4.974391, 4.975267, 
    4.976982, 4.978776, 4.980881, 4.981141, 4.981584, 4.982214, 4.98302, 
    4.983992, 4.985119, 4.986394, 4.987806, 4.989342, 4.990986, 4.992723, 
    4.994529, 4.996365, 4.998188, 4.999933, 5.00151, 5.002803, 5.003664, 
    5.003913,
  // momentumY(28,19, 0-49)
    4.985601, 4.985903, 4.986029, 4.986017, 4.985898, 4.985704, 4.985462, 
    4.985194, 4.98492, 4.984657, 4.984419, 4.984222, 4.984084, 4.984033, 
    4.984104, 4.984866, 4.975602, 4.976647, 4.977926, 4.979109, 4.980078, 
    4.978496, 4.977036, 4.975368, 4.974319, 4.973816, 4.973994, 4.974836, 
    4.976551, 4.978387, 4.980682, 4.980737, 4.980986, 4.981435, 4.982077, 
    4.982903, 4.983911, 4.985092, 4.986441, 4.987948, 4.989601, 4.991385, 
    4.993277, 4.995243, 4.997238, 4.999198, 5.001037, 5.002635, 5.003841, 
    5.004478,
  // momentumY(28,20, 0-49)
    4.986712, 4.987498, 4.98811, 4.988571, 4.988906, 4.989136, 4.989282, 
    4.98936, 4.98939, 4.989389, 4.989371, 4.989356, 4.989365, 4.989432, 
    4.989607, 0, 4.973971, 4.974906, 4.976127, 4.977295, 4.978267, 4.976232, 
    4.974376, 4.972327, 4.970971, 4.970251, 4.970322, 4.971179, 4.973058, 
    4.975195, 4.977999, 4.978202, 4.978607, 4.979215, 4.980005, 4.980972, 
    4.982105, 4.983404, 4.984862, 4.986478, 4.988243, 4.990149, 4.992177, 
    4.994302, 4.996484, 4.998657, 5.000737, 5.002606, 5.004115, 5.005083,
  // momentumY(28,21, 0-49)
    4.987054, 4.987665, 4.988129, 4.988471, 4.988711, 4.988868, 4.988958, 
    4.989, 4.989004, 4.988986, 4.988958, 4.988937, 4.988944, 4.989013, 
    4.989195, 0, 4.970282, 4.971366, 4.97281, 4.974231, 4.975453, 4.973234, 
    4.971309, 4.969253, 4.967992, 4.967446, 4.967751, 4.968876, 4.971061, 
    4.973518, 4.976734, 4.976965, 4.977419, 4.978096, 4.978973, 4.980039, 
    4.981282, 4.982694, 4.984271, 4.986003, 4.987885, 4.989907, 4.992052, 
    4.994292, 4.996589, 4.998882, 5.001087, 5.003087, 5.004737, 5.00586,
  // momentumY(28,22, 0-49)
    4.987328, 4.98778, 4.988113, 4.988348, 4.988502, 4.988594, 4.988635, 
    4.98864, 4.988618, 4.988581, 4.988539, 4.988505, 4.988502, 4.988559, 
    4.988728, 0, 4.967324, 4.968526, 4.970151, 4.971785, 4.973213, 4.970802, 
    4.968777, 4.96666, 4.965425, 4.964967, 4.965406, 4.966697, 4.969078, 
    4.97174, 4.975243, 4.975431, 4.975869, 4.976557, 4.977474, 4.978605, 
    4.979939, 4.981463, 4.98317, 4.985048, 4.987089, 4.989276, 4.991593, 
    4.994008, 4.996481, 4.99895, 5.001328, 5.003502, 5.005326, 5.006629,
  // momentumY(28,23, 0-49)
    4.987549, 4.987857, 4.98807, 4.988206, 4.988283, 4.988314, 4.98831, 
    4.988281, 4.988234, 4.988175, 4.988117, 4.988068, 4.988048, 4.988085, 
    4.988226, 0, 4.964871, 4.966145, 4.967893, 4.969668, 4.971232, 4.968641, 
    4.966502, 4.964304, 4.963049, 4.962618, 4.963121, 4.964503, 4.966997, 
    4.96978, 4.973461, 4.973578, 4.97397, 4.974645, 4.975582, 4.976766, 
    4.978186, 4.979832, 4.981688, 4.983741, 4.985978, 4.988378, 4.990917, 
    4.993559, 4.996259, 4.998947, 5.001537, 5.003915, 5.005933, 5.007423,
  // momentumY(28,24, 0-49)
    4.98774, 4.98791, 4.988009, 4.988055, 4.98806, 4.988034, 4.987987, 
    4.987925, 4.987851, 4.987772, 4.987696, 4.987629, 4.987588, 4.987599, 
    4.987702, 0, 4.963188, 4.964485, 4.966293, 4.968147, 4.969785, 4.967083, 
    4.964877, 4.962627, 4.961349, 4.960917, 4.961437, 4.962847, 4.965379, 
    4.968204, 4.971961, 4.972018, 4.972366, 4.973018, 4.973957, 4.975173, 
    4.976654, 4.97839, 4.980366, 4.982566, 4.984974, 4.987565, 4.990309, 
    4.993167, 4.996087, 4.998994, 5.001799, 5.004381, 5.006594, 5.00827,
  // momentumY(28,25, 0-49)
    4.987918, 4.987956, 4.987947, 4.987906, 4.98784, 4.98776, 4.987669, 
    4.987572, 4.98747, 4.98737, 4.987273, 4.987188, 4.987124, 4.987105, 
    4.987164, 0, 4.961998, 4.963271, 4.96508, 4.966942, 4.96859, 4.965873, 
    4.963664, 4.961417, 4.960142, 4.95971, 4.960229, 4.96163, 4.964145, 
    4.966951, 4.9707, 4.97073, 4.971062, 4.971709, 4.972658, 4.973903, 
    4.975436, 4.977246, 4.979321, 4.981645, 4.984196, 4.986951, 4.989874, 
    4.992926, 4.996044, 4.999156, 5.002161, 5.00494, 5.007341, 5.009192,
  // momentumY(28,26, 0-49)
    4.988102, 4.988014, 4.9879, 4.98777, 4.987633, 4.987494, 4.987355, 
    4.987218, 4.987085, 4.986959, 4.98684, 4.986735, 4.98665, 4.986601, 
    4.986614, 0, 4.96127, 4.962483, 4.964233, 4.96604, 4.967638, 4.965005, 
    4.962867, 4.960688, 4.95945, 4.959028, 4.95953, 4.960891, 4.963342, 
    4.966077, 4.969729, 4.969779, 4.970129, 4.970798, 4.971775, 4.973054, 
    4.974634, 4.976504, 4.978654, 4.98107, 4.983733, 4.986615, 4.989684, 
    4.992893, 4.996181, 4.99947, 5.002655, 5.005613, 5.008188, 5.010205,
  // momentumY(28,27, 0-49)
    4.988311, 4.988101, 4.987882, 4.987662, 4.987448, 4.987243, 4.987047, 
    4.986861, 4.986687, 4.986527, 4.986381, 4.986256, 4.986153, 4.986082, 
    4.986058, 0, 4.961052, 4.962173, 4.963817, 4.96551, 4.967003, 4.964544, 
    4.962538, 4.960472, 4.959287, 4.958868, 4.959324, 4.960605, 4.962934, 
    4.965534, 4.969001, 4.969101, 4.969494, 4.970201, 4.971213, 4.972528, 
    4.974146, 4.97606, 4.978265, 4.980749, 4.983495, 4.986478, 4.989666, 
    4.993008, 4.996446, 4.999894, 5.003249, 5.006377, 5.009121, 5.011301,
  // momentumY(28,28, 0-49)
    4.988558, 4.98823, 4.987906, 4.987594, 4.987296, 4.987011, 4.986745, 
    4.986495, 4.986266, 4.986061, 4.985881, 4.985734, 4.98562, 4.985543, 
    4.985505, 0, 4.961629, 4.962648, 4.964153, 4.965688, 4.967029, 4.964806, 
    4.962961, 4.961018, 4.959865, 4.959403, 4.959753, 4.960879, 4.963003, 
    4.965382, 4.968564, 4.968718, 4.969153, 4.969889, 4.97092, 4.97225, 
    4.973881, 4.975813, 4.978045, 4.980568, 4.983372, 4.986431, 4.989717, 
    4.993181, 4.996759, 5.000366, 5.003891, 5.007196, 5.010116, 5.012463,
  // momentumY(28,29, 0-49)
    4.988853, 4.988415, 4.987991, 4.98758, 4.987185, 4.986807, 4.986447, 
    4.986111, 4.985805, 4.985536, 4.985315, 4.985149, 4.985041, 4.984988, 
    4.984979, 0, 4.96272, 4.963651, 4.965005, 4.966348, 4.967486, 4.965503, 
    4.96379, 4.961924, 4.960732, 4.960146, 4.960302, 4.961183, 4.963007, 
    4.965075, 4.967861, 4.968034, 4.96848, 4.969221, 4.970254, 4.97159, 
    4.973233, 4.975191, 4.977465, 4.980054, 4.982945, 4.986122, 4.989549, 
    4.993178, 4.996941, 5.000747, 5.004481, 5.007996, 5.01112, 5.013654,
  // momentumY(28,30, 0-49)
    4.98853, 4.987349, 4.986206, 4.985108, 4.984058, 4.983053, 4.98209, 
    4.981159, 4.980254, 4.979371, 4.978508, 4.977676, 4.976903, 4.976246, 
    4.975795, 4.974938, 4.965952, 4.966966, 4.968203, 4.969349, 4.970299, 
    4.968656, 4.967254, 4.965686, 4.964678, 4.964137, 4.964175, 4.964772, 
    4.966136, 4.967617, 4.969641, 4.969453, 4.969526, 4.969896, 4.970581, 
    4.971605, 4.972989, 4.974744, 4.976882, 4.979402, 4.982292, 4.98553, 
    4.989075, 4.992872, 4.996842, 5.000887, 5.004877, 5.008653, 5.012033, 
    5.014809,
  // momentumY(28,31, 0-49)
    4.988934, 4.987695, 4.986489, 4.98532, 4.98419, 4.983098, 4.982041, 
    4.981017, 4.980021, 4.979056, 4.978122, 4.977229, 4.976397, 4.975665, 
    4.975098, 4.974432, 4.965597, 4.966311, 4.967228, 4.96806, 4.968717, 
    4.96726, 4.965956, 4.96447, 4.963483, 4.962937, 4.96296, 4.963528, 
    4.964809, 4.96617, 4.967934, 4.96792, 4.968172, 4.968722, 4.969593, 
    4.970803, 4.972375, 4.97432, 4.976649, 4.979359, 4.982438, 4.985861, 
    4.989586, 4.993555, 4.997685, 5.001874, 5.005987, 5.009863, 5.013318, 
    5.016133,
  // momentumY(28,32, 0-49)
    4.989329, 4.988023, 4.986743, 4.985494, 4.984277, 4.983092, 4.98194, 
    4.980819, 4.979729, 4.978675, 4.977658, 4.976685, 4.97577, 4.974939, 
    4.974227, 4.97373, 4.965408, 4.965789, 4.966353, 4.966842, 4.96719, 
    4.965924, 4.964731, 4.963346, 4.9624, 4.961866, 4.961875, 4.962408, 
    4.963588, 4.964805, 4.966289, 4.966444, 4.96687, 4.967595, 4.96864, 
    4.970027, 4.971777, 4.973903, 4.976413, 4.979305, 4.982565, 4.986166, 
    4.990065, 4.994201, 4.998487, 5.002816, 5.007049, 5.011023, 5.014543, 
    5.017394,
  // momentumY(28,33, 0-49)
    4.989703, 4.988327, 4.986968, 4.985633, 4.984324, 4.983045, 4.981792, 
    4.980573, 4.979386, 4.978236, 4.977127, 4.976064, 4.975055, 4.974112, 
    4.973249, 4.97283, 4.965299, 4.96534, 4.965545, 4.96569, 4.965733, 
    4.964666, 4.963603, 4.962349, 4.961465, 4.960958, 4.96096, 4.961446, 
    4.962501, 4.963549, 4.96474, 4.96506, 4.965649, 4.966537, 4.967746, 
    4.969299, 4.971216, 4.973511, 4.976191, 4.979255, 4.982684, 4.986455, 
    4.990518, 4.994809, 4.99924, 5.003698, 5.008042, 5.0121, 5.015676, 
    5.018547,
  // momentumY(28,34, 0-49)
    4.990031, 4.988589, 4.987155, 4.985735, 4.984336, 4.982958, 4.981607, 
    4.980285, 4.978996, 4.977746, 4.976541, 4.975382, 4.974274, 4.973217, 
    4.972211, 4.971758, 4.965207, 4.964923, 4.964778, 4.964593, 4.964345, 
    4.963485, 4.962573, 4.961481, 4.960687, 4.960222, 4.960217, 4.960645, 
    4.961547, 4.962411, 4.963303, 4.963782, 4.964528, 4.965569, 4.966932, 
    4.96864, 4.970713, 4.973166, 4.976003, 4.979225, 4.982812, 4.986735, 
    4.990946, 4.995378, 4.999937, 5.004506, 5.008938, 5.013061, 5.01667, 
    5.019539,
  // momentumY(28,35, 0-49)
    4.990283, 4.988789, 4.987288, 4.985792, 4.984304, 4.982832, 4.981381, 
    4.979957, 4.978567, 4.977216, 4.97591, 4.974653, 4.973446, 4.97228, 
    4.971144, 4.970554, 4.965104, 4.964519, 4.964046, 4.963553, 4.96304, 
    4.962392, 4.96165, 4.960749, 4.960071, 4.959666, 4.959654, 4.960008, 
    4.960733, 4.961397, 4.961999, 4.96263, 4.963524, 4.964712, 4.966218, 
    4.96807, 4.970286, 4.972882, 4.975864, 4.979228, 4.982954, 4.987012, 
    4.991352, 4.995899, 5.000561, 5.005215, 5.009709, 5.013865, 5.017476, 
    5.020309,
  // momentumY(28,36, 0-49)
    4.990426, 4.988896, 4.987345, 4.985782, 4.984218, 4.982658, 4.981112, 
    4.97959, 4.9781, 4.976649, 4.975245, 4.973891, 4.972588, 4.971323, 
    4.970076, 4.969267, 4.964972, 4.964121, 4.963349, 4.962579, 4.961828, 
    4.961393, 4.960837, 4.960156, 4.959619, 4.959288, 4.959268, 4.959536, 
    4.960064, 4.96052, 4.960848, 4.961624, 4.962659, 4.963984, 4.965623, 
    4.967606, 4.969953, 4.972678, 4.975785, 4.979272, 4.983116, 4.987284, 
    4.991723, 4.996358, 5.001091, 5.005792, 5.010311, 5.014461, 5.01803, 
    5.020787,
  // momentumY(28,37, 0-49)
    4.99042, 4.988878, 4.987295, 4.985683, 4.984055, 4.98242, 4.980792, 
    4.97918, 4.977595, 4.97605, 4.974551, 4.973106, 4.971712, 4.970358, 
    4.969019, 4.967945, 4.964811, 4.963729, 4.962691, 4.961675, 4.960719, 
    4.960494, 4.960138, 4.959701, 4.959327, 4.959084, 4.959058, 4.959228, 
    4.959541, 4.959791, 4.959871, 4.960784, 4.961951, 4.963401, 4.965164, 
    4.967265, 4.969728, 4.972565, 4.975777, 4.979362, 4.983298, 4.987546, 
    4.992053, 4.996737, 5.001498, 5.006205, 5.0107, 5.014793, 5.018272, 5.0209,
  // momentumY(28,38, 0-49)
    4.99023, 4.988701, 4.987109, 4.98547, 4.983797, 4.982105, 4.980407, 
    4.978717, 4.977051, 4.97542, 4.973835, 4.972305, 4.97083, 4.969398, 
    4.967984, 4.966624, 4.964621, 4.963344, 4.962071, 4.960845, 4.959713, 
    4.959695, 4.959548, 4.959376, 4.959183, 4.959043, 4.959011, 4.959078, 
    4.959167, 4.959216, 4.959079, 4.960124, 4.961415, 4.962979, 4.964853, 
    4.967059, 4.969621, 4.972549, 4.975846, 4.979504, 4.983499, 4.98779, 
    4.992322, 4.997014, 5.001755, 5.006413, 5.010828, 5.014806, 5.018132, 
    5.020571,
  // momentumY(28,39, 0-49)
    4.98982, 4.988333, 4.986758, 4.985115, 4.983422, 4.981692, 4.979945, 
    4.978195, 4.976461, 4.974759, 4.973101, 4.971496, 4.969948, 4.968448, 
    4.966973, 4.965341, 4.964407, 4.962965, 4.961492, 4.960084, 4.958814, 
    4.958994, 4.959059, 4.959167, 4.959174, 4.959148, 4.959116, 4.959077, 
    4.958942, 4.958804, 4.958484, 4.959653, 4.96106, 4.962731, 4.964701, 
    4.966998, 4.96964, 4.972637, 4.975991, 4.979691, 4.983709, 4.988005, 
    4.992517, 4.997162, 5.001826, 5.006374, 5.010642, 5.014437, 5.017542, 
    5.019726,
  // momentumY(28,40, 0-49)
    4.989163, 4.987743, 4.986215, 4.984596, 4.982908, 4.981167, 4.979392, 
    4.977604, 4.975822, 4.974064, 4.972347, 4.970681, 4.969072, 4.967516, 
    4.965992, 4.964116, 4.964172, 4.962595, 4.960951, 4.959398, 4.958017, 
    4.958385, 4.958663, 4.959061, 4.959281, 4.959382, 4.959355, 4.959212, 
    4.958863, 4.958557, 4.95809, 4.959379, 4.960891, 4.962658, 4.964714, 
    4.967083, 4.969785, 4.972829, 4.97621, 4.979917, 4.983921, 4.988175, 
    4.992615, 4.997153, 5.001677, 5.006044, 5.010092, 5.013627, 5.016435, 
    5.018291,
  // momentumY(28,41, 0-49)
    4.988236, 4.986912, 4.985459, 4.983894, 4.982239, 4.980513, 4.978737, 
    4.976935, 4.975128, 4.973335, 4.971576, 4.969865, 4.968209, 4.966607, 
    4.965042, 4.962963, 4.963916, 4.962226, 4.960443, 4.958775, 4.957313, 
    4.957856, 4.958346, 4.959037, 4.959479, 4.959718, 4.959705, 4.959471, 
    4.958921, 4.958473, 4.957899, 4.959299, 4.96091, 4.962762, 4.96489, 
    4.967316, 4.970056, 4.973118, 4.976497, 4.980174, 4.984117, 4.988278, 
    4.992589, 4.996957, 5.001267, 5.005378, 5.009124, 5.012317, 5.014746, 
    5.016197,
  // momentumY(28,42, 0-49)
    4.98703, 4.98583, 4.984478, 4.982997, 4.981404, 4.979722, 4.977974, 
    4.976183, 4.974374, 4.97257, 4.97079, 4.96905, 4.96736, 4.965723, 
    4.964126, 4.961891, 4.963639, 4.961859, 4.95996, 4.958206, 4.956691, 
    4.957398, 4.958096, 4.959077, 4.959745, 4.96013, 4.960144, 4.959831, 
    4.959105, 4.958547, 4.957901, 4.959409, 4.961112, 4.963038, 4.965222, 
    4.967688, 4.970444, 4.973498, 4.976838, 4.980443, 4.98428, 4.988293, 
    4.992411, 4.996538, 5.000558, 5.00433, 5.007689, 5.010449, 5.012415, 
    5.013385,
  // momentumY(28,43, 0-49)
    4.98554, 4.984489, 4.983268, 4.981898, 4.980398, 4.978789, 4.977099, 
    4.975349, 4.973565, 4.971771, 4.96999, 4.96824, 4.96653, 4.964868, 
    4.963245, 4.9609, 4.963339, 4.961486, 4.959499, 4.957683, 4.956139, 
    4.956997, 4.957892, 4.959154, 4.960049, 4.960588, 4.96064, 4.960272, 
    4.959402, 4.958764, 4.958083, 4.959694, 4.961483, 4.963474, 4.965702, 
    4.968185, 4.970934, 4.973947, 4.977213, 4.980706, 4.984384, 4.988188, 
    4.992046, 4.99586, 4.999508, 5.002852, 5.005733, 5.007973, 5.009391, 
    5.009803,
  // momentumY(28,44, 0-49)
    4.983782, 4.982901, 4.981836, 4.980603, 4.979224, 4.977719, 4.976113, 
    4.974431, 4.972697, 4.970939, 4.969179, 4.967435, 4.965723, 4.964047, 
    4.962406, 4.959991, 4.963014, 4.961103, 4.959048, 4.957194, 4.955643, 
    4.956639, 4.95772, 4.959247, 4.960364, 4.961061, 4.961168, 4.960768, 
    4.95979, 4.959107, 4.958425, 4.960135, 4.962002, 4.964049, 4.966306, 
    4.968788, 4.971504, 4.974445, 4.977598, 4.980931, 4.984395, 4.987931, 
    4.991458, 4.994877, 4.99807, 5.000897, 5.003209, 5.00484, 5.005627, 
    5.005414,
  // momentumY(28,45, 0-49)
    4.981774, 4.981083, 4.980196, 4.979126, 4.977894, 4.97652, 4.975028, 
    4.973438, 4.971782, 4.970082, 4.968363, 4.966645, 4.964943, 4.963265, 
    4.961613, 4.959162, 4.962658, 4.960703, 4.958603, 4.956729, 4.955187, 
    4.956307, 4.957557, 4.959331, 4.960659, 4.961514, 4.961693, 4.961289, 
    4.960246, 4.959553, 4.958898, 4.960707, 4.962646, 4.964738, 4.967009, 
    4.969471, 4.972126, 4.974962, 4.977961, 4.981081, 4.984278, 4.987478, 
    4.990602, 4.993547, 4.996198, 4.998419, 5.000072, 5.001008, 5.001089, 
    5.000189,
  // momentumY(28,46, 0-49)
    4.979548, 4.979063, 4.978371, 4.977488, 4.976427, 4.975208, 4.973854, 
    4.972385, 4.970828, 4.969208, 4.96755, 4.965873, 4.964198, 4.96253, 
    4.960874, 4.958412, 4.962271, 4.960286, 4.958158, 4.95628, 4.95476, 
    4.955986, 4.957387, 4.959378, 4.960902, 4.961915, 4.96218, 4.961805, 
    4.96074, 4.960072, 4.959472, 4.961374, 4.96338, 4.965507, 4.967777, 
    4.970197, 4.972763, 4.975461, 4.978261, 4.981122, 4.983987, 4.986786, 
    4.989431, 4.991823, 4.993845, 4.995374, 4.996282, 4.996446, 4.995755, 
    4.994122,
  // momentumY(28,47, 0-49)
    4.977147, 4.976876, 4.976397, 4.975716, 4.974848, 4.973806, 4.972611, 
    4.971286, 4.96985, 4.968332, 4.966752, 4.965134, 4.963496, 4.961848, 
    4.960196, 4.957739, 4.96185, 4.959847, 4.957707, 4.955839, 4.95435, 
    4.955663, 4.957192, 4.959366, 4.961065, 4.962229, 4.962596, 4.962281, 
    4.96124, 4.96063, 4.960107, 4.962099, 4.964166, 4.966316, 4.96857, 
    4.970924, 4.973373, 4.975894, 4.978453, 4.981, 4.983474, 4.985802, 
    4.987894, 4.98965, 4.990963, 4.991716, 4.991806, 4.991132, 4.989618, 
    4.987222,
  // momentumY(28,48, 0-49)
    4.974618, 4.974567, 4.974308, 4.973845, 4.973186, 4.972341, 4.971326, 
    4.970162, 4.968867, 4.967466, 4.965981, 4.964435, 4.962846, 4.961228, 
    4.959587, 4.957145, 4.961398, 4.959391, 4.957252, 4.9554, 4.953947, 
    4.955328, 4.956959, 4.959277, 4.961123, 4.962427, 4.962908, 4.962682, 
    4.96171, 4.961189, 4.960761, 4.962839, 4.964956, 4.967119, 4.969338, 
    4.971605, 4.973905, 4.976213, 4.978484, 4.980662, 4.982685, 4.984473, 
    4.98594, 4.986984, 4.987511, 4.987416, 4.986622, 4.985056, 4.982687, 
    4.979521,
  // momentumY(28,49, 0-49)
    4.971751, 4.97187, 4.971794, 4.971513, 4.971032, 4.970352, 4.969482, 
    4.968434, 4.96722, 4.965861, 4.964369, 4.962768, 4.961073, 4.959293, 
    4.957433, 4.953966, 4.963982, 4.960976, 4.957507, 4.954463, 4.952083, 
    4.955269, 4.95878, 4.963472, 4.966963, 4.969119, 4.969381, 4.967987, 
    4.964842, 4.962405, 4.959975, 4.962437, 4.964849, 4.967206, 4.969516, 
    4.971771, 4.973949, 4.976017, 4.977924, 4.979613, 4.981015, 4.982051, 
    4.98264, 4.982693, 4.982131, 4.980882, 4.978908, 4.976194, 4.972773, 
    4.968725,
  // momentumY(29,0, 0-49)
    4.971556, 4.973361, 4.974815, 4.975937, 4.976742, 4.97725, 4.977488, 
    4.977488, 4.977288, 4.976929, 4.976456, 4.97591, 4.975338, 4.97478, 
    4.974274, 4.973676, 4.973505, 4.973238, 4.973083, 4.97306, 4.973165, 
    4.973533, 4.973971, 4.974497, 4.975105, 4.975779, 4.976512, 4.977307, 
    4.978165, 4.979098, 4.980094, 4.981372, 4.982794, 4.984384, 4.986169, 
    4.988163, 4.99037, 4.992781, 4.995366, 4.998078, 5.000845, 5.003565, 
    5.00611, 5.008316, 5.009995, 5.010931, 5.010883, 5.009605, 5.006854, 
    5.002412,
  // momentumY(29,1, 0-49)
    4.97285, 4.9746, 4.976003, 4.977079, 4.977844, 4.97832, 4.978535, 
    4.978521, 4.978314, 4.977955, 4.977486, 4.976948, 4.976385, 4.975832, 
    4.975327, 4.974553, 4.974493, 4.974136, 4.97386, 4.973703, 4.973669, 
    4.97404, 4.974442, 4.974925, 4.975485, 4.976109, 4.976785, 4.977513, 
    4.978296, 4.979141, 4.980009, 4.981315, 4.982766, 4.984389, 4.986212, 
    4.988253, 4.990514, 4.992992, 4.995659, 4.998469, 5.001352, 5.00421, 
    5.006918, 5.009318, 5.011222, 5.012416, 5.012663, 5.011715, 5.009322, 
    5.005255,
  // momentumY(29,2, 0-49)
    4.974152, 4.975846, 4.977199, 4.978231, 4.97896, 4.979407, 4.979604, 
    4.979578, 4.979369, 4.979012, 4.978549, 4.978021, 4.977464, 4.976915, 
    4.976405, 4.97546, 4.975474, 4.975027, 4.974627, 4.974336, 4.974163, 
    4.974525, 4.97488, 4.975307, 4.975816, 4.976388, 4.977014, 4.977693, 
    4.978423, 4.979195, 4.979949, 4.981287, 4.982766, 4.984417, 4.986269, 
    4.988337, 4.990631, 4.993144, 4.995852, 4.998711, 5.001653, 5.004588, 
    5.007389, 5.009909, 5.011964, 5.013349, 5.013828, 5.013155, 5.011086, 
    5.007389,
  // momentumY(29,3, 0-49)
    4.975455, 4.977093, 4.978398, 4.979385, 4.98008, 4.980501, 4.980679, 
    4.980646, 4.980434, 4.980083, 4.979627, 4.979106, 4.978555, 4.978006, 
    4.977489, 4.976379, 4.976416, 4.975876, 4.975358, 4.974937, 4.97463, 
    4.974973, 4.975272, 4.975631, 4.976077, 4.976596, 4.977183, 4.977833, 
    4.978536, 4.979261, 4.979921, 4.981289, 4.982796, 4.98447, 4.98634, 
    4.988424, 4.990729, 4.993248, 4.995963, 4.998829, 5.001781, 5.004733, 
    5.007569, 5.010144, 5.012286, 5.013795, 5.014449, 5.014008, 5.01223, 
    5.008885,
  // momentumY(29,4, 0-49)
    4.976765, 4.978344, 4.979596, 4.980538, 4.981195, 4.981589, 4.981749, 
    4.981706, 4.981493, 4.981143, 4.980695, 4.980181, 4.979634, 4.979084, 
    4.978553, 4.977294, 4.977292, 4.976662, 4.976037, 4.975495, 4.975061, 
    4.975371, 4.975604, 4.975881, 4.976256, 4.976723, 4.97728, 4.97792, 
    4.978625, 4.979328, 4.979919, 4.98132, 4.982853, 4.984545, 4.986426, 
    4.988512, 4.990811, 4.993315, 4.996003, 4.99884, 5.00176, 5.004683, 
    5.0075, 5.010075, 5.012246, 5.013824, 5.0146, 5.014348, 5.012831, 5.009826,
  // momentumY(29,5, 0-49)
    4.978075, 4.97959, 4.980784, 4.981678, 4.982295, 4.98266, 4.9828, 
    4.982745, 4.982529, 4.982182, 4.981737, 4.981228, 4.980682, 4.980126, 
    4.979578, 4.978192, 4.978077, 4.977365, 4.976644, 4.975996, 4.975449, 
    4.975712, 4.975867, 4.976048, 4.976345, 4.976757, 4.977293, 4.977944, 
    4.978681, 4.97939, 4.979939, 4.981371, 4.982926, 4.984634, 4.986518, 
    4.988595, 4.990872, 4.99334, 4.995981, 4.998755, 5.001609, 5.004463, 
    5.007217, 5.009746, 5.0119, 5.013502, 5.014358, 5.014255, 5.012973, 
    5.010293,
  // momentumY(29,6, 0-49)
    4.979375, 4.980821, 4.981953, 4.982794, 4.983367, 4.983699, 4.983816, 
    4.983747, 4.983525, 4.983177, 4.982736, 4.982229, 4.981682, 4.981119, 
    4.980551, 4.979065, 4.978755, 4.977969, 4.97717, 4.976434, 4.975792, 
    4.975995, 4.976058, 4.976129, 4.976338, 4.976693, 4.977218, 4.977898, 
    4.978695, 4.979438, 4.979978, 4.981435, 4.98301, 4.984728, 4.986608, 
    4.988667, 4.990908, 4.993323, 4.995894, 4.998584, 5.00134, 5.004094, 
    5.006751, 5.009197, 5.011295, 5.012885, 5.013788, 5.013808, 5.012739, 
    5.010373,
  // momentumY(29,7, 0-49)
    4.980656, 4.982026, 4.983089, 4.983871, 4.984396, 4.98469, 4.984782, 
    4.984697, 4.984466, 4.984116, 4.983675, 4.98317, 4.982621, 4.982047, 
    4.981458, 4.979904, 4.979315, 4.978468, 4.977612, 4.976809, 4.976092, 
    4.976218, 4.97618, 4.976123, 4.976236, 4.976532, 4.977053, 4.977777, 
    4.978659, 4.979466, 4.980029, 4.981503, 4.983092, 4.984814, 4.986686, 
    4.988718, 4.99091, 4.993259, 4.995742, 4.998327, 5.000965, 5.003592, 
    5.006126, 5.008463, 5.010478, 5.012031, 5.012955, 5.013077, 5.012204, 
    5.010143,
  // momentumY(29,8, 0-49)
    4.981897, 4.983184, 4.984174, 4.984893, 4.985365, 4.98562, 4.985681, 
    4.985578, 4.985337, 4.984982, 4.984541, 4.984036, 4.983485, 4.982903, 
    4.982292, 4.980708, 4.979747, 4.978858, 4.977969, 4.977125, 4.976357, 
    4.976388, 4.976235, 4.976039, 4.976047, 4.976282, 4.976804, 4.977584, 
    4.978576, 4.979469, 4.980087, 4.981573, 4.983167, 4.984883, 4.986736, 
    4.988731, 4.990869, 4.993138, 4.99552, 4.997984, 5.000488, 5.002973, 
    5.005363, 5.007573, 5.009488, 5.010984, 5.011919, 5.012128, 5.011442, 
    5.009677,
  // momentumY(29,9, 0-49)
    4.983086, 4.984283, 4.985192, 4.985842, 4.986258, 4.986469, 4.986499, 
    4.986375, 4.986122, 4.985764, 4.985322, 4.984818, 4.984266, 4.983675, 
    4.983043, 4.981473, 4.980051, 4.97914, 4.978247, 4.977389, 4.976596, 
    4.976516, 4.976236, 4.97589, 4.975786, 4.975957, 4.976483, 4.977327, 
    4.978443, 4.979445, 4.980153, 4.981635, 4.983224, 4.984926, 4.986752, 
    4.988701, 4.990771, 4.992952, 4.995222, 4.997556, 4.999913, 5.002243, 
    5.004482, 5.006552, 5.008358, 5.009792, 5.010726, 5.011018, 5.010513, 
    5.009043,
  // momentumY(29,10, 0-49)
    4.984201, 4.9853, 4.986125, 4.986701, 4.987059, 4.987222, 4.987219, 
    4.987072, 4.986808, 4.986445, 4.986005, 4.985502, 4.984953, 4.984358, 
    4.983712, 4.982196, 4.980223, 4.979319, 4.978451, 4.977612, 4.976825, 
    4.976614, 4.976199, 4.975692, 4.975474, 4.975579, 4.976107, 4.977016, 
    4.978267, 4.979397, 4.980227, 4.981689, 4.983257, 4.984932, 4.986719, 
    4.988612, 4.990606, 4.992688, 4.99484, 4.997035, 4.99924, 5.001411, 
    5.003496, 5.005424, 5.007121, 5.008492, 5.009428, 5.009802, 5.009476, 
    5.008297,
  // momentumY(29,11, 0-49)
    4.985221, 4.986217, 4.986951, 4.987451, 4.987747, 4.987863, 4.987825, 
    4.987659, 4.987381, 4.987016, 4.986578, 4.986081, 4.985535, 4.984943, 
    4.984293, 4.982874, 4.980265, 4.979398, 4.978592, 4.977806, 4.977054, 
    4.9767, 4.976141, 4.975471, 4.975133, 4.975172, 4.9757, 4.976673, 
    4.978061, 4.979329, 4.980305, 4.981731, 4.983263, 4.984897, 4.98663, 
    4.988455, 4.990363, 4.992339, 4.994365, 4.996418, 4.998469, 5.000483, 
    5.002415, 5.004209, 5.005803, 5.007117, 5.008061, 5.008524, 5.008382, 
    5.00749,
  // momentumY(29,12, 0-49)
    4.986129, 4.987016, 4.987657, 4.988077, 4.98831, 4.988379, 4.988306, 
    4.988117, 4.987829, 4.987461, 4.98703, 4.986541, 4.986005, 4.985423, 
    4.984781, 4.983505, 4.980176, 4.979388, 4.978679, 4.977983, 4.977303, 
    4.976789, 4.976083, 4.975247, 4.974793, 4.974764, 4.975285, 4.976314, 
    4.977836, 4.979246, 4.980394, 4.981762, 4.983236, 4.98481, 4.986475, 
    4.98822, 4.99003, 4.991893, 4.99379, 4.9957, 4.997602, 4.999462, 5.00125, 
    5.002921, 5.004425, 5.005697, 5.00666, 5.007222, 5.007267, 5.006666,
  // momentumY(29,13, 0-49)
    4.98691, 4.987683, 4.988225, 4.988565, 4.988734, 4.988751, 4.988646, 
    4.988435, 4.988138, 4.98777, 4.987345, 4.98687, 4.986352, 4.985789, 
    4.985172, 4.984077, 4.97996, 4.979289, 4.978722, 4.978153, 4.97758, 
    4.976897, 4.976046, 4.975048, 4.974481, 4.974383, 4.974892, 4.975965, 
    4.977607, 4.979157, 4.980497, 4.98178, 4.983175, 4.984669, 4.986247, 
    4.987896, 4.989599, 4.991342, 4.993107, 4.994876, 4.996633, 4.998353, 
    5.000012, 5.001576, 5.003008, 5.004256, 5.005257, 5.005929, 5.00617, 
    5.005861,
  // momentumY(29,14, 0-49)
    4.987552, 4.988207, 4.988649, 4.988905, 4.989006, 4.988974, 4.988832, 
    4.988601, 4.988295, 4.987929, 4.987513, 4.987056, 4.986562, 4.986031, 
    4.985457, 4.984582, 4.97962, 4.979108, 4.978724, 4.978326, 4.977896, 
    4.977039, 4.976047, 4.974896, 4.974222, 4.974059, 4.974547, 4.975648, 
    4.977391, 4.979072, 4.980613, 4.981785, 4.983075, 4.984465, 4.985938, 
    4.987476, 4.989061, 4.990677, 4.992309, 4.993942, 4.995565, 4.997159, 
    4.998707, 5.000188, 5.001571, 5.002817, 5.003875, 5.004673, 5.00512, 
    5.005102,
  // momentumY(29,15, 0-49)
    4.988047, 4.988579, 4.988916, 4.989087, 4.989118, 4.989033, 4.988854, 
    4.988601, 4.988286, 4.987922, 4.98752, 4.987084, 4.986623, 4.986136, 
    4.985628, 4.985004, 4.979161, 4.978853, 4.978694, 4.978505, 4.978258, 
    4.977225, 4.976098, 4.97481, 4.974041, 4.973814, 4.974275, 4.975384, 
    4.977204, 4.978997, 4.980742, 4.981776, 4.982933, 4.984197, 4.985542, 
    4.986952, 4.988406, 4.989891, 4.991391, 4.992896, 4.994396, 4.995882, 
    4.997343, 4.998764, 5.000125, 5.001397, 5.002533, 5.003475, 5.004138, 
    5.004411,
  // momentumY(29,16, 0-49)
    4.988392, 4.988796, 4.989022, 4.989101, 4.98906, 4.98892, 4.988703, 
    4.988425, 4.988101, 4.987741, 4.987353, 4.986944, 4.986523, 4.986093, 
    4.985668, 4.985326, 4.978594, 4.978531, 4.978637, 4.978697, 4.978667, 
    4.977459, 4.976213, 4.974801, 4.973953, 4.973667, 4.974092, 4.975191, 
    4.977059, 4.978941, 4.980883, 4.98175, 4.982749, 4.983858, 4.985055, 
    4.986319, 4.987631, 4.988978, 4.990348, 4.991733, 4.993127, 4.994525, 
    4.995924, 4.997314, 4.998682, 5.000005, 5.001247, 5.002351, 5.00324, 
    5.003806,
  // momentumY(29,17, 0-49)
    4.988588, 4.988854, 4.988962, 4.988945, 4.988825, 4.988625, 4.988366, 
    4.988063, 4.987727, 4.98737, 4.986999, 4.986622, 4.986247, 4.985889, 
    4.985566, 4.98553, 4.977942, 4.97816, 4.978563, 4.978907, 4.979125, 
    4.977752, 4.9764, 4.974884, 4.973968, 4.973629, 4.97401, 4.97508, 
    4.976967, 4.978909, 4.981034, 4.981708, 4.982517, 4.983448, 4.984474, 
    4.985574, 4.986732, 4.987938, 4.98918, 4.990454, 4.991757, 4.99309, 
    4.994452, 4.995841, 4.997247, 4.998652, 5.000022, 5.001309, 5.002435, 
    5.003295,
  // momentumY(29,18, 0-49)
    4.988639, 4.988755, 4.988736, 4.98861, 4.988406, 4.988142, 4.987838, 
    4.987507, 4.987159, 4.986805, 4.986453, 4.986112, 4.985792, 4.985513, 
    4.98531, 4.985602, 4.977243, 4.977769, 4.978495, 4.979146, 4.979639, 
    4.978107, 4.976663, 4.97506, 4.974088, 4.973702, 4.974034, 4.975058, 
    4.976934, 4.978906, 4.981187, 4.981641, 4.982238, 4.982964, 4.983794, 
    4.984714, 4.985708, 4.986764, 4.987881, 4.989054, 4.990283, 4.991574, 
    4.992928, 4.994346, 4.995821, 4.997337, 4.998865, 5.000354, 5.001728, 
    5.002884,
  // momentumY(29,19, 0-49)
    4.98855, 4.988499, 4.988338, 4.988094, 4.987796, 4.987462, 4.987109, 
    4.986747, 4.986388, 4.986039, 4.985707, 4.985406, 4.985149, 4.984963, 
    4.984892, 4.98553, 4.976555, 4.977411, 4.978475, 4.979445, 4.980222, 
    4.978542, 4.977019, 4.975341, 4.974323, 4.973892, 4.974168, 4.975128, 
    4.976965, 4.978934, 4.981341, 4.981552, 4.981909, 4.982407, 4.983021, 
    4.98374, 4.984555, 4.985459, 4.98645, 4.98753, 4.988702, 4.989972, 
    4.991343, 4.99282, 4.994395, 4.996053, 4.997765, 4.999477, 5.001114, 
    5.002572,
  // momentumY(29,20, 0-49)
    4.989048, 4.989503, 4.989847, 4.990098, 4.99027, 4.990378, 4.990433, 
    4.990442, 4.990415, 4.99036, 4.990286, 4.990209, 4.990146, 4.990134, 
    4.990227, 0, 4.975359, 4.976153, 4.977207, 4.978203, 4.979018, 4.976952, 
    4.975087, 4.973069, 4.971763, 4.971109, 4.97125, 4.972173, 4.974099, 
    4.976275, 4.979077, 4.979346, 4.979769, 4.980332, 4.98101, 4.981788, 
    4.982655, 4.983606, 4.984644, 4.985774, 4.987006, 4.988348, 4.98981, 
    4.991399, 4.993111, 4.994935, 4.996837, 4.99877, 5.000656, 5.002386,
  // momentumY(29,21, 0-49)
    4.988827, 4.98916, 4.989402, 4.98957, 4.989676, 4.989734, 4.989754, 
    4.989744, 4.989711, 4.98966, 4.9896, 4.989542, 4.989507, 4.989525, 
    4.989647, 0, 4.972302, 4.973264, 4.974558, 4.975825, 4.976907, 4.974704, 
    4.972797, 4.970784, 4.969567, 4.96906, 4.969389, 4.970522, 4.972679, 
    4.975086, 4.978195, 4.978409, 4.978792, 4.979332, 4.980003, 4.980789, 
    4.981676, 4.98266, 4.983741, 4.984922, 4.986211, 4.987618, 4.989153, 
    4.990819, 4.992617, 4.994532, 4.996534, 4.998575, 5.000577, 5.002439,
  // momentumY(29,22, 0-49)
    4.988561, 4.988786, 4.988936, 4.989029, 4.989077, 4.989089, 4.989075, 
    4.989043, 4.988997, 4.988944, 4.988889, 4.988842, 4.988819, 4.988848, 
    4.988978, 0, 4.970036, 4.971129, 4.972622, 4.974118, 4.975419, 4.973063, 
    4.971076, 4.969011, 4.967807, 4.967357, 4.967772, 4.969004, 4.971275, 
    4.973795, 4.977079, 4.977161, 4.977431, 4.977885, 4.978497, 4.979252, 
    4.980139, 4.981151, 4.982288, 4.983549, 4.98494, 4.986465, 4.988132, 
    4.989944, 4.991897, 4.993972, 4.996139, 4.998345, 5.000515, 5.002546,
  // momentumY(29,23, 0-49)
    4.988266, 4.988394, 4.988463, 4.988487, 4.988479, 4.988449, 4.988403, 
    4.988348, 4.988288, 4.988229, 4.988175, 4.988132, 4.988114, 4.988146, 
    4.988268, 0, 4.968285, 4.969466, 4.971102, 4.972762, 4.974215, 4.971715, 
    4.969638, 4.967495, 4.966257, 4.9658, 4.966229, 4.967482, 4.969783, 
    4.972326, 4.975673, 4.975587, 4.97571, 4.976046, 4.976573, 4.977282, 
    4.978163, 4.979208, 4.980416, 4.981785, 4.983315, 4.985008, 4.986862, 
    4.988875, 4.991038, 4.993327, 4.995707, 4.998123, 5.000495, 5.002719,
  // momentumY(29,24, 0-49)
    4.987961, 4.987996, 4.987988, 4.98795, 4.987892, 4.987821, 4.987746, 
    4.98767, 4.987597, 4.987533, 4.987478, 4.987438, 4.987423, 4.987453, 
    4.987559, 0, 4.967278, 4.968503, 4.970228, 4.971992, 4.973543, 4.970967, 
    4.968838, 4.966646, 4.96537, 4.964878, 4.96527, 4.966482, 4.968736, 
    4.971223, 4.974539, 4.974289, 4.974264, 4.97447, 4.974896, 4.975535, 
    4.976382, 4.977432, 4.978685, 4.980134, 4.981779, 4.98362, 4.985648, 
    4.987854, 4.990224, 4.992731, 4.995331, 4.997964, 5.000548, 5.002974,
  // momentumY(29,25, 0-49)
    4.98766, 4.987607, 4.987528, 4.98743, 4.987325, 4.987216, 4.987114, 
    4.987021, 4.986938, 4.986869, 4.986818, 4.986785, 4.986776, 4.986806, 
    4.986895, 0, 4.966704, 4.967937, 4.969695, 4.971504, 4.973098, 4.970532, 
    4.968414, 4.966226, 4.964935, 4.964411, 4.964749, 4.965886, 4.968045, 
    4.970422, 4.973626, 4.973247, 4.973096, 4.973194, 4.973528, 4.974099, 
    4.974905, 4.975947, 4.977223, 4.97873, 4.980465, 4.982426, 4.984601, 
    4.986979, 4.989538, 4.992245, 4.995053, 4.997897, 5.000687, 5.003313,
  // momentumY(29,26, 0-49)
    4.987382, 4.987242, 4.987093, 4.986938, 4.986787, 4.986643, 4.986514, 
    4.986403, 4.986313, 4.986247, 4.986204, 4.986186, 4.986193, 4.986231, 
    4.986312, 0, 4.966497, 4.967708, 4.969454, 4.971251, 4.972836, 4.970378, 
    4.968344, 4.96622, 4.96495, 4.964405, 4.96468, 4.965718, 4.967741, 
    4.969964, 4.972982, 4.972522, 4.972288, 4.972305, 4.972567, 4.97308, 
    4.973845, 4.974867, 4.976147, 4.977685, 4.979478, 4.981522, 4.983808, 
    4.986319, 4.989032, 4.991911, 4.994902, 4.997937, 5.000921, 5.003737,
  // momentumY(29,27, 0-49)
    4.987139, 4.986915, 4.986696, 4.986484, 4.986285, 4.986104, 4.98595, 
    4.985823, 4.985728, 4.985668, 4.985642, 4.98565, 4.985687, 4.985753, 
    4.985845, 0, 4.966663, 4.967835, 4.969529, 4.971269, 4.972798, 4.970535, 
    4.968647, 4.966635, 4.965405, 4.964836, 4.965031, 4.96594, 4.967781, 
    4.969799, 4.972559, 4.972056, 4.971772, 4.971733, 4.971939, 4.972399, 
    4.97312, 4.974112, 4.975377, 4.97692, 4.978742, 4.980838, 4.983202, 
    4.985818, 4.98866, 4.991688, 4.994846, 4.998058, 5.001228, 5.00423,
  // momentumY(29,28, 0-49)
    4.986944, 4.986639, 4.986349, 4.986075, 4.985826, 4.985606, 4.985421, 
    4.985277, 4.985176, 4.985127, 4.985129, 4.985179, 4.985272, 4.985394, 
    4.985533, 0, 4.967456, 4.968589, 4.970207, 4.971852, 4.973289, 4.971285, 
    4.969576, 4.967695, 4.966493, 4.965866, 4.965929, 4.966646, 4.968236, 
    4.969983, 4.972405, 4.971874, 4.97155, 4.971457, 4.971603, 4.971999, 
    4.97266, 4.973596, 4.97482, 4.976341, 4.978161, 4.980283, 4.982701, 
    4.985398, 4.98835, 4.991515, 4.994833, 4.998222, 5.001579, 5.004774,
  // momentumY(29,29, 0-49)
    4.986812, 4.986425, 4.986062, 4.985725, 4.98542, 4.985151, 4.984928, 
    4.984759, 4.984652, 4.984617, 4.984658, 4.984773, 4.984951, 4.985173, 
    4.985413, 0, 4.968573, 4.969682, 4.971219, 4.972744, 4.974048, 4.972317, 
    4.970768, 4.968982, 4.967752, 4.967, 4.966858, 4.967312, 4.968576, 
    4.969975, 4.971971, 4.971394, 4.971013, 4.970857, 4.970938, 4.971271, 
    4.971876, 4.97277, 4.97397, 4.975489, 4.977334, 4.979512, 4.982013, 
    4.984826, 4.987921, 4.991253, 4.994759, 4.998352, 5.001921, 5.005327,
  // momentumY(29,30, 0-49)
    4.986113, 4.985028, 4.983992, 4.98301, 4.982088, 4.981229, 4.980436, 
    4.979713, 4.979061, 4.978491, 4.978013, 4.977649, 4.977439, 4.977439, 
    4.97774, 4.978108, 4.970986, 4.972597, 4.974332, 4.975877, 4.977121, 
    4.975759, 4.974507, 4.972983, 4.97189, 4.971142, 4.970854, 4.971008, 
    4.971807, 4.972627, 4.973881, 4.972935, 4.972168, 4.971625, 4.971332, 
    4.971322, 4.971624, 4.972265, 4.973269, 4.974652, 4.976425, 4.978588, 
    4.981136, 4.984048, 4.987289, 4.990808, 4.994532, 4.998365, 5.002188, 
    5.005852,
  // momentumY(29,31, 0-49)
    4.986139, 4.985011, 4.983933, 4.982914, 4.981956, 4.981061, 4.980238, 
    4.979491, 4.978826, 4.978252, 4.977779, 4.977426, 4.97722, 4.9772, 
    4.977429, 4.977726, 4.970573, 4.971944, 4.973413, 4.974692, 4.97569, 
    4.974526, 4.973392, 4.971966, 4.970906, 4.970163, 4.969861, 4.969983, 
    4.970693, 4.971382, 4.972375, 4.971571, 4.970947, 4.970544, 4.970392, 
    4.970518, 4.970953, 4.971724, 4.972854, 4.974358, 4.976247, 4.978524, 
    4.98118, 4.984198, 4.987542, 4.991161, 4.99498, 4.998902, 5.002809, 
    5.006545,
  // momentumY(29,32, 0-49)
    4.98621, 4.985024, 4.983895, 4.982825, 4.981821, 4.980885, 4.980024, 
    4.979245, 4.978554, 4.977959, 4.97747, 4.977098, 4.97686, 4.97678, 
    4.976899, 4.977179, 4.970335, 4.971414, 4.972563, 4.973532, 4.974247, 
    4.973269, 4.972249, 4.970926, 4.969913, 4.969187, 4.968878, 4.968968, 
    4.969584, 4.97014, 4.970872, 4.970227, 4.969762, 4.969515, 4.969513, 
    4.969784, 4.970358, 4.971261, 4.972516, 4.974138, 4.976139, 4.978522, 
    4.98128, 4.984394, 4.98783, 4.991536, 4.99544, 4.999442, 5.00342, 5.007222,
  // momentumY(29,33, 0-49)
    4.986322, 4.985071, 4.98388, 4.982752, 4.981695, 4.980709, 4.979803, 
    4.978983, 4.978255, 4.977623, 4.977099, 4.976686, 4.976392, 4.976228, 
    4.976206, 4.976455, 4.97019, 4.970946, 4.971748, 4.972381, 4.972796, 
    4.971999, 4.971097, 4.969897, 4.968946, 4.968251, 4.967942, 4.968001, 
    4.96851, 4.968925, 4.969399, 4.968927, 4.968636, 4.968554, 4.968711, 
    4.969135, 4.969853, 4.970891, 4.972271, 4.97401, 4.976117, 4.978599, 
    4.981448, 4.984647, 4.988163, 4.991945, 4.995917, 4.999985, 5.00402, 
    5.007871,
  // momentumY(29,34, 0-49)
    4.986467, 4.98515, 4.983893, 4.982704, 4.981585, 4.980543, 4.979585, 
    4.978714, 4.977937, 4.977258, 4.976682, 4.976209, 4.97584, 4.975573, 
    4.9754, 4.975558, 4.97007, 4.970491, 4.970932, 4.971223, 4.971337, 
    4.970714, 4.969939, 4.968884, 4.968016, 4.967366, 4.967063, 4.967083, 
    4.967473, 4.967741, 4.967969, 4.967685, 4.967576, 4.96767, 4.967996, 
    4.96858, 4.969448, 4.970625, 4.972131, 4.973985, 4.976196, 4.978769, 
    4.981701, 4.984973, 4.988553, 4.992392, 4.996415, 5.000526, 5.0046, 
    5.008479,
  // momentumY(29,35, 0-49)
    4.986632, 4.985251, 4.98393, 4.982677, 4.981496, 4.980392, 4.979373, 
    4.978443, 4.977607, 4.976867, 4.976226, 4.97568, 4.975222, 4.97484, 
    4.974514, 4.974512, 4.969934, 4.970024, 4.970108, 4.97006, 4.969883, 
    4.969428, 4.968791, 4.967904, 4.967138, 4.966548, 4.966253, 4.966227, 
    4.96648, 4.966601, 4.966601, 4.96651, 4.966591, 4.96687, 4.967371, 
    4.968122, 4.969146, 4.970466, 4.972102, 4.974071, 4.976381, 4.979041, 
    4.982045, 4.985377, 4.989005, 4.99288, 4.996932, 5.001062, 5.005144, 
    5.009022,
  // momentumY(29,36, 0-49)
    4.986797, 4.985363, 4.983984, 4.98267, 4.981424, 4.980255, 4.97917, 
    4.978174, 4.977268, 4.976458, 4.97574, 4.97511, 4.974553, 4.974052, 
    4.973577, 4.973351, 4.969756, 4.969531, 4.96927, 4.968902, 4.968448, 
    4.968158, 4.967667, 4.966969, 4.966328, 4.965811, 4.965522, 4.965443, 
    4.965545, 4.965516, 4.965311, 4.965418, 4.965693, 4.96616, 4.966842, 
    4.967765, 4.968948, 4.970416, 4.972183, 4.974266, 4.976675, 4.979414, 
    4.98248, 4.985857, 4.989515, 4.993406, 4.99746, 5.001577, 5.005634, 
    5.009474,
  // momentumY(29,37, 0-49)
    4.986938, 4.985464, 4.984036, 4.982665, 4.981359, 4.980126, 4.978973, 
    4.977904, 4.976924, 4.976033, 4.97523, 4.974505, 4.973844, 4.973222, 
    4.972605, 4.972109, 4.969525, 4.969004, 4.968421, 4.967756, 4.967048, 
    4.966916, 4.966578, 4.966092, 4.965594, 4.965162, 4.964882, 4.964739, 
    4.964676, 4.9645, 4.964114, 4.96442, 4.964892, 4.965548, 4.966413, 
    4.96751, 4.968857, 4.970472, 4.972372, 4.974567, 4.97707, 4.979882, 
    4.983001, 4.986409, 4.990077, 4.993959, 4.997983, 5.002053, 5.006046, 
    5.009804,
  // momentumY(29,38, 0-49)
    4.987028, 4.985529, 4.984065, 4.982647, 4.981288, 4.979993, 4.978771, 
    4.977629, 4.976569, 4.975593, 4.974696, 4.973871, 4.973101, 4.972361, 
    4.971611, 4.970821, 4.969233, 4.968444, 4.967564, 4.96663, 4.965697, 
    4.965714, 4.965539, 4.96528, 4.964942, 4.964607, 4.964337, 4.964119, 
    4.963884, 4.963566, 4.96303, 4.963531, 4.964195, 4.965038, 4.966087, 
    4.967357, 4.968866, 4.970628, 4.972659, 4.974966, 4.977559, 4.980438, 
    4.983595, 4.98702, 4.990678, 4.994521, 4.998483, 5.002466, 5.006349, 
    5.009973,
  // momentumY(29,39, 0-49)
    4.98703, 4.985528, 4.984045, 4.982595, 4.981189, 4.97984, 4.978554, 
    4.977337, 4.976196, 4.975132, 4.974139, 4.97321, 4.972332, 4.971474, 
    4.970599, 4.969515, 4.96888, 4.967854, 4.966705, 4.965531, 4.964404, 
    4.964564, 4.964558, 4.964538, 4.964377, 4.964149, 4.963889, 4.963593, 
    4.96318, 4.96273, 4.962073, 4.962762, 4.963613, 4.964639, 4.965863, 
    4.967302, 4.96897, 4.970879, 4.973037, 4.975451, 4.978129, 4.981064, 
    4.984251, 4.987672, 4.991296, 4.995074, 4.998935, 5.002787, 5.006506, 
    5.009941,
  // momentumY(29,40, 0-49)
    4.986917, 4.985433, 4.98395, 4.982483, 4.981046, 4.979649, 4.978304, 
    4.977018, 4.975799, 4.974646, 4.973557, 4.972527, 4.971539, 4.970568, 
    4.969579, 4.968217, 4.968469, 4.967233, 4.965849, 4.964469, 4.963177, 
    4.963475, 4.963636, 4.963868, 4.963894, 4.963784, 4.963535, 4.963162, 
    4.962571, 4.962003, 4.961255, 4.962122, 4.963151, 4.964351, 4.965744, 
    4.967346, 4.969165, 4.971212, 4.973492, 4.976008, 4.978761, 4.981743, 
    4.984945, 4.988344, 4.991908, 4.995585, 4.999307, 5.002978, 5.006479, 
    5.00966,
  // momentumY(29,41, 0-49)
    4.986656, 4.985214, 4.983752, 4.982286, 4.980833, 4.979402, 4.978008, 
    4.976662, 4.975368, 4.97413, 4.97295, 4.971819, 4.970726, 4.969647, 
    4.968551, 4.96694, 4.968, 4.966581, 4.964995, 4.963443, 4.96202, 
    4.962448, 4.962779, 4.963267, 4.963491, 4.963505, 4.963273, 4.962823, 
    4.962065, 4.961395, 4.960584, 4.96162, 4.962814, 4.964176, 4.965727, 
    4.967481, 4.969442, 4.971618, 4.974011, 4.976619, 4.979436, 4.98245, 
    4.98565, 4.989006, 4.992481, 4.996022, 4.99956, 5.002998, 5.00622, 5.00908,
  // momentumY(29,42, 0-49)
    4.986219, 4.984845, 4.983426, 4.981982, 4.980528, 4.979081, 4.977652, 
    4.976253, 4.974894, 4.973581, 4.972313, 4.971088, 4.969896, 4.968716, 
    4.96752, 4.965698, 4.967477, 4.965904, 4.964147, 4.962456, 4.960933, 
    4.961483, 4.961984, 4.962727, 4.963152, 4.963299, 4.96309, 4.962575, 
    4.961663, 4.96091, 4.960064, 4.961257, 4.962603, 4.964114, 4.96581, 
    4.967701, 4.969793, 4.972085, 4.974578, 4.977262, 4.980129, 4.98316, 
    4.986334, 4.989621, 4.992977, 4.996344, 4.99965, 5.0028, 5.00568, 5.00815,
  // momentumY(29,43, 0-49)
    4.985586, 4.984303, 4.982952, 4.981551, 4.980116, 4.978669, 4.977219, 
    4.975782, 4.97437, 4.97299, 4.971644, 4.970334, 4.969049, 4.967778, 
    4.966492, 4.964496, 4.966899, 4.965197, 4.963301, 4.961505, 4.959913, 
    4.960582, 4.961247, 4.96224, 4.962868, 4.963152, 4.962977, 4.962408, 
    4.961366, 4.960551, 4.959695, 4.961031, 4.962516, 4.964162, 4.965988, 
    4.968001, 4.970206, 4.972599, 4.975173, 4.977917, 4.980814, 4.983839, 
    4.986966, 4.990153, 4.993352, 4.996504, 4.999529, 5.002333, 5.004804, 
    5.006812,
  // momentumY(29,44, 0-49)
    4.984741, 4.983572, 4.98231, 4.980974, 4.979583, 4.978152, 4.9767, 
    4.975242, 4.973791, 4.972355, 4.970943, 4.969557, 4.968193, 4.966837, 
    4.96547, 4.96334, 4.966269, 4.964459, 4.962457, 4.960586, 4.958953, 
    4.959734, 4.960559, 4.961791, 4.962621, 4.963047, 4.962915, 4.962311, 
    4.961167, 4.960318, 4.959472, 4.96094, 4.96255, 4.964314, 4.966252, 
    4.968369, 4.970668, 4.973141, 4.975777, 4.978558, 4.981461, 4.984454, 
    4.987502, 4.990557, 4.993561, 4.996449, 4.999139, 5.001537, 5.003535, 
    5.00501,
  // momentumY(29,45, 0-49)
    4.983676, 4.982643, 4.981495, 4.980247, 4.978919, 4.977528, 4.976092, 
    4.974628, 4.973153, 4.971678, 4.970212, 4.968764, 4.967327, 4.965899, 
    4.964459, 4.962228, 4.965582, 4.963693, 4.96161, 4.959693, 4.958048, 
    4.958934, 4.95991, 4.961367, 4.962389, 4.962958, 4.962886, 4.962271, 
    4.961058, 4.960199, 4.959386, 4.960973, 4.962695, 4.964563, 4.966595, 
    4.968796, 4.971167, 4.973697, 4.976369, 4.979159, 4.982038, 4.984967, 
    4.987901, 4.990783, 4.99355, 4.996124, 4.998423, 5.000354, 5.001812, 
    5.002688,
  // momentumY(29,46, 0-49)
    4.982392, 4.981516, 4.980502, 4.979363, 4.978121, 4.976789, 4.97539, 
    4.973942, 4.972459, 4.970959, 4.969454, 4.967954, 4.96646, 4.964968, 
    4.963467, 4.961162, 4.96484, 4.962892, 4.96076, 4.958823, 4.957186, 
    4.958171, 4.959288, 4.960949, 4.962153, 4.962865, 4.962866, 4.962266, 
    4.961024, 4.960183, 4.959423, 4.961119, 4.962938, 4.964893, 4.967002, 
    4.969267, 4.971686, 4.974245, 4.976924, 4.979692, 4.982513, 4.985339, 
    4.988117, 4.990781, 4.993258, 4.995465, 4.997318, 4.998721, 4.999578, 
    4.999793,
  // momentumY(29,47, 0-49)
    4.980901, 4.9802, 4.979339, 4.97833, 4.977193, 4.975943, 4.9746, 
    4.973184, 4.971713, 4.970206, 4.968677, 4.967138, 4.965598, 4.964054, 
    4.962501, 4.960147, 4.964045, 4.96206, 4.959902, 4.957967, 4.956358, 
    4.957434, 4.958677, 4.960518, 4.961888, 4.96274, 4.962831, 4.962277, 
    4.961047, 4.960255, 4.959564, 4.961359, 4.963265, 4.965293, 4.967459, 
    4.969764, 4.972204, 4.974763, 4.977415, 4.980123, 4.982846, 4.985526, 
    4.988099, 4.990493, 4.992628, 4.994412, 4.995758, 4.996574, 4.996771, 
    4.996272,
  // momentumY(29,48, 0-49)
    4.979223, 4.978709, 4.978018, 4.977159, 4.976146, 4.974998, 4.973732, 
    4.972368, 4.970926, 4.969428, 4.967888, 4.966326, 4.96475, 4.963166, 
    4.961571, 4.959184, 4.963201, 4.961198, 4.959035, 4.957121, 4.955557, 
    4.956709, 4.958065, 4.960053, 4.961572, 4.96256, 4.962756, 4.96228, 
    4.961107, 4.960392, 4.959789, 4.961674, 4.963654, 4.965738, 4.967942, 
    4.970265, 4.972701, 4.975228, 4.977816, 4.980423, 4.983, 4.985481, 
    4.987796, 4.989864, 4.991597, 4.992898, 4.993679, 4.993851, 4.993337, 
    4.992082,
  // momentumY(29,49, 0-49)
    4.977364, 4.976999, 4.976442, 4.975697, 4.974771, 4.973678, 4.972433, 
    4.97105, 4.96955, 4.967954, 4.966277, 4.964537, 4.96275, 4.960918, 
    4.959042, 4.955583, 4.965085, 4.962095, 4.958641, 4.955575, 4.95313, 
    4.956073, 4.959288, 4.963607, 4.966753, 4.968592, 4.96859, 4.966987, 
    4.963706, 4.96112, 4.958558, 4.960826, 4.963123, 4.965455, 4.967843, 
    4.970289, 4.972789, 4.975318, 4.977843, 4.980316, 4.982681, 4.984867, 
    4.986794, 4.988374, 4.989514, 4.990113, 4.990091, 4.989372, 4.987904, 
    4.98567 ;
}
