netcdf netCdfTest {
dimensions:
	x = 10 ;
	y = 10 ;
variables:
	float height(x, y) ;
	float momentumX(x, y) ;
	float momentumY(x, y) ;
	float bathymetry(x, y) ;
	float time ;
	float timeStep ;
	float writingStepsCount ;
	float simulationSizeX ;
	float simulationSizeY ;
	float offsetX ;
	float offsetY ;
data:

 height =
  // height(0, 0-9)
    100, 1100, 2100, 3100, 4100, 5100, 6100, 7100, 8100, 9100,
  // height(1, 0-9)
    200, 1200, 2200, 3200, 4200, 5200, 6200, 7200, 8200, 9200,
  // height(2, 0-9)
    300, 1300, 2300, 3300, 4300, 5300, 6300, 7300, 8300, 9300,
  // height(3, 0-9)
    400, 1400, 2400, 3400, 4400, 5400, 6400, 7400, 8400, 9400,
  // height(4, 0-9)
    500, 1500, 2500, 3500, 4500, 5500, 6500, 7500, 8500, 9500,
  // height(5, 0-9)
    600, 1600, 2600, 3600, 4600, 5600, 6600, 7600, 8600, 9600,
  // height(6, 0-9)
    700, 1700, 2700, 3700, 4700, 5700, 6700, 7700, 8700, 9700,
  // height(7, 0-9)
    800, 1800, 2800, 3800, 4800, 5800, 6800, 7800, 8800, 9800,
  // height(8, 0-9)
    900, 1900, 2900, 3900, 4900, 5900, 6900, 7900, 8900, 9900,
  // height(9, 0-9)
    1000, 2000, 3000, 4000, 5000, 6000, 7000, 8000, 9000, 10000 ;

 momentumX =
  // momentumX(0, 0-9)
    13, 143, 273, 403, 533, 663, 793, 923, 1053, 1183,
  // momentumX(1, 0-9)
    26, 156, 286, 416, 546, 676, 806, 936, 1066, 1196,
  // momentumX(2, 0-9)
    39, 169, 299, 429, 559, 689, 819, 949, 1079, 1209,
  // momentumX(3, 0-9)
    52, 182, 312, 442, 572, 702, 832, 962, 1092, 1222,
  // momentumX(4, 0-9)
    65, 195, 325, 455, 585, 715, 845, 975, 1105, 1235,
  // momentumX(5, 0-9)
    78, 208, 338, 468, 598, 728, 858, 988, 1118, 1248,
  // momentumX(6, 0-9)
    91, 221, 351, 481, 611, 741, 871, 1001, 1131, 1261,
  // momentumX(7, 0-9)
    104, 234, 364, 494, 624, 754, 884, 1014, 1144, 1274,
  // momentumX(8, 0-9)
    117, 247, 377, 507, 637, 767, 897, 1027, 1157, 1287,
  // momentumX(9, 0-9)
    130, 260, 390, 520, 650, 780, 910, 1040, 1170, 1300 ;

 momentumY =
  // momentumY(0, 0-9)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  // momentumY(1, 0-9)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  // momentumY(2, 0-9)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  // momentumY(3, 0-9)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  // momentumY(4, 0-9)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  // momentumY(5, 0-9)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  // momentumY(6, 0-9)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  // momentumY(7, 0-9)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  // momentumY(8, 0-9)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  // momentumY(9, 0-9)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 bathymetry =
  // bathymetry(0, 0-9)
    1.844674e+19, 1.844674e+19, 1.844674e+19, 1.844674e+19, 1.844674e+19, 
    1.844674e+19, 1.844674e+19, 1.844674e+19, 1.844674e+19, 1.844674e+19,
  // bathymetry(1, 0-9)
    1.844674e+19, 1.844674e+19, 1.844674e+19, 1.844674e+19, 1.844674e+19, 
    1.844674e+19, 1.844674e+19, 1.844674e+19, 1.844674e+19, 1.844674e+19,
  // bathymetry(2, 0-9)
    1.844674e+19, 1.844674e+19, 1.844674e+19, 1.844674e+19, 1.844674e+19, 
    1.844674e+19, 1.844674e+19, 1.844674e+19, 1.844674e+19, 1.844674e+19,
  // bathymetry(3, 0-9)
    1.844674e+19, 1.844674e+19, 1.844674e+19, 1.844674e+19, 1.844674e+19, 
    1.844674e+19, 1.844674e+19, 1.844674e+19, 1.844674e+19, 1.844674e+19,
  // bathymetry(4, 0-9)
    1.844674e+19, 1.844674e+19, 1.844674e+19, 1.844674e+19, 1.844674e+19, 
    1.844674e+19, 1.844674e+19, 1.844674e+19, 1.844674e+19, 1.844674e+19,
  // bathymetry(5, 0-9)
    1.844674e+19, 1.844674e+19, 1.844674e+19, 1.844674e+19, 1.844674e+19, 
    1.844674e+19, 1.844674e+19, 1.844674e+19, 1.844674e+19, 1.844674e+19,
  // bathymetry(6, 0-9)
    1.844674e+19, 1.844674e+19, 1.844674e+19, 1.844674e+19, 1.844674e+19, 
    1.844674e+19, 1.844674e+19, 1.844674e+19, 1.844674e+19, 1.844674e+19,
  // bathymetry(7, 0-9)
    1.844674e+19, 1.844674e+19, 1.844674e+19, 1.844674e+19, 1.844674e+19, 
    1.844674e+19, 1.844674e+19, 1.844674e+19, 1.844674e+19, 1.844674e+19,
  // bathymetry(8, 0-9)
    1.844674e+19, 1.844674e+19, 1.844674e+19, 1.844674e+19, 1.844674e+19, 
    1.844674e+19, 1.844674e+19, 1.844674e+19, 1.844674e+19, 1.844674e+19,
  // bathymetry(9, 0-9)
    1.844674e+19, 1.844674e+19, 1.844674e+19, 1.844674e+19, 1.844674e+19, 
    1.844674e+19, 1.844674e+19, 1.844674e+19, 1.844674e+19, 1.844674e+19 ;

 time = 7.826369e-05 ;

 timeStep = 131 ;

 writingStepsCount = 0 ;

 simulationSizeX = 10 ;

 simulationSizeY = 10 ;

 offsetX = -5 ;

 offsetY = -5 ;
}
