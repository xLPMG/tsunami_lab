netcdf artificialtsunami_displ_1000 {
dimensions:
	x = 100 ;
	y = 100 ;
variables:
	float x(x) ;
	float y(y) ;
	float z(y, x) ;

// global attributes:
		:Conventions = "COARDS" ;
data:

 x = -495, -485, -475, -465, -455, -445, -435, -425, -415, -405, -395, -385, 
    -375, -365, -355, -345, -335, -325, -315, -305, -295, -285, -275, -265, 
    -255, -245, -235, -225, -215, -205, -195, -185, -175, -165, -155, -145, 
    -135, -125, -115, -105, -95, -85, -75, -65, -55, -45, -35, -25, -15, -5, 
    5, 15, 25, 35, 45, 55, 65, 75, 85, 95, 105, 115, 125, 135, 145, 155, 165, 
    175, 185, 195, 205, 215, 225, 235, 245, 255, 265, 275, 285, 295, 305, 
    315, 325, 335, 345, 355, 365, 375, 385, 395, 405, 415, 425, 435, 445, 
    455, 465, 475, 485, 495 ;

 y = -495, -485, -475, -465, -455, -445, -435, -425, -415, -405, -395, -385, 
    -375, -365, -355, -345, -335, -325, -315, -305, -295, -285, -275, -265, 
    -255, -245, -235, -225, -215, -205, -195, -185, -175, -165, -155, -145, 
    -135, -125, -115, -105, -95, -85, -75, -65, -55, -45, -35, -25, -15, -5, 
    5, 15, 25, 35, 45, 55, 65, 75, 85, 95, 105, 115, 125, 135, 145, 155, 165, 
    175, 185, 195, 205, 215, 225, 235, 245, 255, 265, 275, 285, 295, 305, 
    315, 325, 335, 345, 355, 365, 375, 385, 395, 405, 415, 425, 435, 445, 
    455, 465, 475, 485, 495 ;

 z =
  // z(0, 0-99)
    0.00312537, 0.009363777, 0.01556523, 0.02170525, 0.02775962, 0.03370442, 
    0.03951621, 0.04517205, 0.05064962, 0.0559273, 0.06098425, 0.06580053, 
    0.07035712, 0.07463605, 0.07862043, 0.08229452, 0.08564384, 0.08865515, 
    0.09131659, 0.09361763, 0.09554922, 0.09710371, 0.09827499, 0.09905841, 
    0.0994509, 0.0994509, 0.09905841, 0.09827499, 0.09710371, 0.09554922, 
    0.09361763, 0.09131659, 0.08865515, 0.08564384, 0.08229452, 0.07862043, 
    0.07463605, 0.07035712, 0.06580053, 0.06098425, 0.0559273, 0.05064962, 
    0.04517205, 0.03951621, 0.03370442, 0.02775962, 0.02170525, 0.01556523, 
    0.009363777, 0.00312537, -0.00312537, -0.009363777, -0.01556523, 
    -0.02170525, -0.02775962, -0.03370442, -0.03951621, -0.04517205, 
    -0.05064962, -0.0559273, -0.06098425, -0.06580053, -0.07035712, 
    -0.07463605, -0.07862043, -0.08229452, -0.08564384, -0.08865515, 
    -0.09131659, -0.09361763, -0.09554922, -0.09710371, -0.09827499, 
    -0.09905841, -0.0994509, -0.0994509, -0.09905841, -0.09827499, 
    -0.09710371, -0.09554922, -0.09361763, -0.09131659, -0.08865515, 
    -0.08564384, -0.08229452, -0.07862043, -0.07463605, -0.07035712, 
    -0.06580053, -0.06098425, -0.0559273, -0.05064962, -0.04517205, 
    -0.03951621, -0.03370442, -0.02775962, -0.02170525, -0.01556523, 
    -0.009363777, -0.00312537,
  // z(1, 0-99)
    0.009281879, 0.02780901, 0.04622639, 0.06446133, 0.08244187, 0.1000971, 
    0.1173572, 0.1341542, 0.1504217, 0.1660956, 0.181114, 0.1954177, 
    0.2089501, 0.2216578, 0.2334908, 0.2444023, 0.2543493, 0.2632924, 
    0.2711965, 0.2780303, 0.2837668, 0.2883834, 0.2918619, 0.2941886, 
    0.2953542, 0.2953542, 0.2941886, 0.2918619, 0.2883834, 0.2837668, 
    0.2780303, 0.2711965, 0.2632924, 0.2543493, 0.2444023, 0.2334908, 
    0.2216578, 0.2089501, 0.1954177, 0.181114, 0.1660956, 0.1504217, 
    0.1341542, 0.1173572, 0.1000971, 0.08244187, 0.06446133, 0.04622639, 
    0.02780901, 0.009281879, -0.009281879, -0.02780901, -0.04622639, 
    -0.06446133, -0.08244187, -0.1000971, -0.1173572, -0.1341542, -0.1504217, 
    -0.1660956, -0.181114, -0.1954177, -0.2089501, -0.2216578, -0.2334908, 
    -0.2444023, -0.2543493, -0.2632924, -0.2711965, -0.2780303, -0.2837668, 
    -0.2883834, -0.2918619, -0.2941886, -0.2953542, -0.2953542, -0.2941886, 
    -0.2918619, -0.2883834, -0.2837668, -0.2780303, -0.2711965, -0.2632924, 
    -0.2543493, -0.2444023, -0.2334908, -0.2216578, -0.2089501, -0.1954177, 
    -0.181114, -0.1660956, -0.1504217, -0.1341542, -0.1173572, -0.1000971, 
    -0.08244187, -0.06446133, -0.04622639, -0.02780901, -0.009281879,
  // z(2, 0-99)
    0.01531275, 0.0458778, 0.0762618, 0.1063448, 0.1360082, 0.1651347, 
    0.1936096, 0.2213204, 0.2481577, 0.2740156, 0.2987922, 0.3223895, 
    0.3447146, 0.3656791, 0.3852006, 0.4032018, 0.4196118, 0.4343657, 
    0.4474054, 0.4586794, 0.4681432, 0.4757594, 0.4814981, 0.4853365, 
    0.4872594, 0.4872594, 0.4853365, 0.4814981, 0.4757594, 0.4681432, 
    0.4586794, 0.4474054, 0.4343657, 0.4196118, 0.4032018, 0.3852006, 
    0.3656791, 0.3447146, 0.3223895, 0.2987922, 0.2740156, 0.2481577, 
    0.2213204, 0.1936096, 0.1651347, 0.1360082, 0.1063448, 0.0762618, 
    0.0458778, 0.01531275, -0.01531275, -0.0458778, -0.0762618, -0.1063448, 
    -0.1360082, -0.1651347, -0.1936096, -0.2213204, -0.2481577, -0.2740156, 
    -0.2987922, -0.3223895, -0.3447146, -0.3656791, -0.3852006, -0.4032018, 
    -0.4196118, -0.4343657, -0.4474054, -0.4586794, -0.4681432, -0.4757594, 
    -0.4814981, -0.4853365, -0.4872594, -0.4872594, -0.4853365, -0.4814981, 
    -0.4757594, -0.4681432, -0.4586794, -0.4474054, -0.4343657, -0.4196118, 
    -0.4032018, -0.3852006, -0.3656791, -0.3447146, -0.3223895, -0.2987922, 
    -0.2740156, -0.2481577, -0.2213204, -0.1936096, -0.1651347, -0.1360082, 
    -0.1063448, -0.0762618, -0.0458778, -0.01531275,
  // z(3, 0-99)
    0.02121797, 0.06357016, 0.1056715, 0.1473558, 0.1884585, 0.2288175, 
    0.2682734, 0.3066706, 0.3438575, 0.3796873, 0.4140187, 0.4467162, 
    0.4776506, 0.5067, 0.5337497, 0.5586929, 0.5814312, 0.6018749, 0.6199433, 
    0.635565, 0.6486784, 0.6592318, 0.6671835, 0.6725021, 0.6751667, 
    0.6751667, 0.6725021, 0.6671835, 0.6592318, 0.6486784, 0.635565, 
    0.6199433, 0.6018749, 0.5814312, 0.5586929, 0.5337497, 0.5067, 0.4776506, 
    0.4467162, 0.4140187, 0.3796873, 0.3438575, 0.3066706, 0.2682734, 
    0.2288175, 0.1884585, 0.1473558, 0.1056715, 0.06357016, 0.02121797, 
    -0.02121797, -0.06357016, -0.1056715, -0.1473558, -0.1884585, -0.2288175, 
    -0.2682734, -0.3066706, -0.3438575, -0.3796873, -0.4140187, -0.4467162, 
    -0.4776506, -0.5067, -0.5337497, -0.5586929, -0.5814312, -0.6018749, 
    -0.6199433, -0.635565, -0.6486784, -0.6592318, -0.6671835, -0.6725021, 
    -0.6751667, -0.6751667, -0.6725021, -0.6671835, -0.6592318, -0.6486784, 
    -0.635565, -0.6199433, -0.6018749, -0.5814312, -0.5586929, -0.5337497, 
    -0.5067, -0.4776506, -0.4467162, -0.4140187, -0.3796873, -0.3438575, 
    -0.3066706, -0.2682734, -0.2288175, -0.1884585, -0.1473558, -0.1056715, 
    -0.06357016, -0.02121797,
  // z(4, 0-99)
    0.02699755, 0.0808861, 0.1344554, 0.1874941, 0.2397929, 0.2911452, 
    0.3413486, 0.3902048, 0.4375211, 0.4831107, 0.5267936, 0.5683975, 
    0.6077583, 0.6447204, 0.6791382, 0.7108757, 0.7398078, 0.7658201, 
    0.7888101, 0.808687, 0.8253724, 0.8388004, 0.8489181, 0.8556855, 
    0.8590759, 0.8590759, 0.8556855, 0.8489181, 0.8388004, 0.8253724, 
    0.808687, 0.7888101, 0.7658201, 0.7398078, 0.7108757, 0.6791382, 
    0.6447204, 0.6077583, 0.5683975, 0.5267936, 0.4831107, 0.4375211, 
    0.3902048, 0.3413486, 0.2911452, 0.2397929, 0.1874941, 0.1344554, 
    0.0808861, 0.02699755, -0.02699755, -0.0808861, -0.1344554, -0.1874941, 
    -0.2397929, -0.2911452, -0.3413486, -0.3902048, -0.4375211, -0.4831107, 
    -0.5267936, -0.5683975, -0.6077583, -0.6447204, -0.6791382, -0.7108757, 
    -0.7398078, -0.7658201, -0.7888101, -0.808687, -0.8253724, -0.8388004, 
    -0.8489181, -0.8556855, -0.8590759, -0.8590759, -0.8556855, -0.8489181, 
    -0.8388004, -0.8253724, -0.808687, -0.7888101, -0.7658201, -0.7398078, 
    -0.7108757, -0.6791382, -0.6447204, -0.6077583, -0.5683975, -0.5267936, 
    -0.4831107, -0.4375211, -0.3902048, -0.3413486, -0.2911452, -0.2397929, 
    -0.1874941, -0.1344554, -0.0808861, -0.02699755,
  // z(5, 0-99)
    0.03265148, 0.09782559, 0.1626136, 0.2267599, 0.2900113, 0.3521181, 
    0.4128352, 0.4719231, 0.5291486, 0.5842857, 0.6371169, 0.6874337, 
    0.7350375, 0.7797405, 0.8213661, 0.8597503, 0.8947414, 0.9262013, 
    0.954006, 0.9780456, 0.9982253, 1.014465, 1.026702, 1.034887, 1.038987, 
    1.038987, 1.034887, 1.026702, 1.014465, 0.9982253, 0.9780456, 0.954006, 
    0.9262013, 0.8947414, 0.8597503, 0.8213661, 0.7797405, 0.7350375, 
    0.6874337, 0.6371169, 0.5842857, 0.5291486, 0.4719231, 0.4128352, 
    0.3521181, 0.2900113, 0.2267599, 0.1626136, 0.09782559, 0.03265148, 
    -0.03265148, -0.09782559, -0.1626136, -0.2267599, -0.2900113, -0.3521181, 
    -0.4128352, -0.4719231, -0.5291486, -0.5842857, -0.6371169, -0.6874337, 
    -0.7350375, -0.7797405, -0.8213661, -0.8597503, -0.8947414, -0.9262013, 
    -0.954006, -0.9780456, -0.9982253, -1.014465, -1.026702, -1.034887, 
    -1.038987, -1.038987, -1.034887, -1.026702, -1.014465, -0.9982253, 
    -0.9780456, -0.954006, -0.9262013, -0.8947414, -0.8597503, -0.8213661, 
    -0.7797405, -0.7350375, -0.6874337, -0.6371169, -0.5842857, -0.5291486, 
    -0.4719231, -0.4128352, -0.3521181, -0.2900113, -0.2267599, -0.1626136, 
    -0.09782559, -0.03265148,
  // z(6, 0-99)
    0.03817978, 0.1143887, 0.1901461, 0.2651531, 0.3391137, 0.411736, 
    0.4827332, 0.5518255, 0.6187398, 0.6832123, 0.7449885, 0.8038245, 
    0.8594883, 0.91176, 0.9604334, 1.005316, 1.046232, 1.083018, 1.115531, 
    1.143641, 1.167237, 1.186227, 1.200535, 1.210106, 1.2149, 1.2149, 
    1.210106, 1.200535, 1.186227, 1.167237, 1.143641, 1.115531, 1.083018, 
    1.046232, 1.005316, 0.9604334, 0.91176, 0.8594883, 0.8038245, 0.7449885, 
    0.6832123, 0.6187398, 0.5518255, 0.4827332, 0.411736, 0.3391137, 
    0.2651531, 0.1901461, 0.1143887, 0.03817978, -0.03817978, -0.1143887, 
    -0.1901461, -0.2651531, -0.3391137, -0.411736, -0.4827332, -0.5518255, 
    -0.6187398, -0.6832123, -0.7449885, -0.8038245, -0.8594883, -0.91176, 
    -0.9604334, -1.005316, -1.046232, -1.083018, -1.115531, -1.143641, 
    -1.167237, -1.186227, -1.200535, -1.210106, -1.2149, -1.2149, -1.210106, 
    -1.200535, -1.186227, -1.167237, -1.143641, -1.115531, -1.083018, 
    -1.046232, -1.005316, -0.9604334, -0.91176, -0.8594883, -0.8038245, 
    -0.7449885, -0.6832123, -0.6187398, -0.5518255, -0.4827332, -0.411736, 
    -0.3391137, -0.2651531, -0.1901461, -0.1143887, -0.03817978,
  // z(7, 0-99)
    0.04358243, 0.1305753, 0.2170528, 0.3026738, 0.3871002, 0.4699989, 
    0.5510427, 0.6299118, 0.706295, 0.7798907, 0.8504086, 0.9175702, 
    0.9811106, 1.040779, 1.09634, 1.147574, 1.19428, 1.236272, 1.273385, 
    1.305472, 1.332407, 1.354084, 1.370418, 1.381342, 1.386815, 1.386815, 
    1.381342, 1.370418, 1.354084, 1.332407, 1.305472, 1.273385, 1.236272, 
    1.19428, 1.147574, 1.09634, 1.040779, 0.9811106, 0.9175702, 0.8504086, 
    0.7798907, 0.706295, 0.6299118, 0.5510427, 0.4699989, 0.3871002, 
    0.3026738, 0.2170528, 0.1305753, 0.04358243, -0.04358243, -0.1305753, 
    -0.2170528, -0.3026738, -0.3871002, -0.4699989, -0.5510427, -0.6299118, 
    -0.706295, -0.7798907, -0.8504086, -0.9175702, -0.9811106, -1.040779, 
    -1.09634, -1.147574, -1.19428, -1.236272, -1.273385, -1.305472, 
    -1.332407, -1.354084, -1.370418, -1.381342, -1.386815, -1.386815, 
    -1.381342, -1.370418, -1.354084, -1.332407, -1.305472, -1.273385, 
    -1.236272, -1.19428, -1.147574, -1.09634, -1.040779, -0.9811106, 
    -0.9175702, -0.8504086, -0.7798907, -0.706295, -0.6299118, -0.5510427, 
    -0.4699989, -0.3871002, -0.3026738, -0.2170528, -0.1305753, -0.04358243,
  // z(8, 0-99)
    0.04885944, 0.1463855, 0.2433338, 0.3393218, 0.4339707, 0.5269068, 
    0.6177635, 0.7061822, 0.7918139, 0.8743207, 0.9533769, 1.028671, 
    1.099905, 1.166798, 1.229086, 1.286524, 1.338884, 1.385961, 1.427567, 
    1.46354, 1.493737, 1.518039, 1.536349, 1.548597, 1.554732, 1.554732, 
    1.548597, 1.536349, 1.518039, 1.493737, 1.46354, 1.427567, 1.385961, 
    1.338884, 1.286524, 1.229086, 1.166798, 1.099905, 1.028671, 0.9533769, 
    0.8743207, 0.7918139, 0.7061822, 0.6177635, 0.5269068, 0.4339707, 
    0.3393218, 0.2433338, 0.1463855, 0.04885944, -0.04885944, -0.1463855, 
    -0.2433338, -0.3393218, -0.4339707, -0.5269068, -0.6177635, -0.7061822, 
    -0.7918139, -0.8743207, -0.9533769, -1.028671, -1.099905, -1.166798, 
    -1.229086, -1.286524, -1.338884, -1.385961, -1.427567, -1.46354, 
    -1.493737, -1.518039, -1.536349, -1.548597, -1.554732, -1.554732, 
    -1.548597, -1.536349, -1.518039, -1.493737, -1.46354, -1.427567, 
    -1.385961, -1.338884, -1.286524, -1.229086, -1.166798, -1.099905, 
    -1.028671, -0.9533769, -0.8743207, -0.7918139, -0.7061822, -0.6177635, 
    -0.5269068, -0.4339707, -0.3393218, -0.2433338, -0.1463855, -0.04885944,
  // z(9, 0-99)
    0.0540108, 0.1618192, 0.2689891, 0.3750973, 0.4797252, 0.5824599, 
    0.6828958, 0.7806367, 0.8752967, 0.9665024, 1.053894, 1.137126, 1.21587, 
    1.289816, 1.358672, 1.422165, 1.480046, 1.532086, 1.578079, 1.617844, 
    1.651225, 1.678089, 1.69833, 1.711869, 1.718652, 1.718652, 1.711869, 
    1.69833, 1.678089, 1.651225, 1.617844, 1.578079, 1.532086, 1.480046, 
    1.422165, 1.358672, 1.289816, 1.21587, 1.137126, 1.053894, 0.9665024, 
    0.8752967, 0.7806367, 0.6828958, 0.5824599, 0.4797252, 0.3750973, 
    0.2689891, 0.1618192, 0.0540108, -0.0540108, -0.1618192, -0.2689891, 
    -0.3750973, -0.4797252, -0.5824599, -0.6828958, -0.7806367, -0.8752967, 
    -0.9665024, -1.053894, -1.137126, -1.21587, -1.289816, -1.358672, 
    -1.422165, -1.480046, -1.532086, -1.578079, -1.617844, -1.651225, 
    -1.678089, -1.69833, -1.711869, -1.718652, -1.718652, -1.711869, 
    -1.69833, -1.678089, -1.651225, -1.617844, -1.578079, -1.532086, 
    -1.480046, -1.422165, -1.358672, -1.289816, -1.21587, -1.137126, 
    -1.053894, -0.9665024, -0.8752967, -0.7806367, -0.6828958, -0.5824599, 
    -0.4797252, -0.3750973, -0.2689891, -0.1618192, -0.0540108,
  // z(10, 0-99)
    0.05903652, 0.1768766, 0.2940186, 0.4100002, 0.5243638, 0.6366579, 
    0.7464395, 0.8532751, 0.9567434, 1.056436, 1.151959, 1.242936, 1.329007, 
    1.409834, 1.485096, 1.554498, 1.617765, 1.674647, 1.72492, 1.768385, 
    1.804872, 1.834236, 1.85636, 1.871159, 1.878573, 1.878573, 1.871159, 
    1.85636, 1.834236, 1.804872, 1.768385, 1.72492, 1.674647, 1.617765, 
    1.554498, 1.485096, 1.409834, 1.329007, 1.242936, 1.151959, 1.056436, 
    0.9567434, 0.8532751, 0.7464395, 0.6366579, 0.5243638, 0.4100002, 
    0.2940186, 0.1768766, 0.05903652, -0.05903652, -0.1768766, -0.2940186, 
    -0.4100002, -0.5243638, -0.6366579, -0.7464395, -0.8532751, -0.9567434, 
    -1.056436, -1.151959, -1.242936, -1.329007, -1.409834, -1.485096, 
    -1.554498, -1.617765, -1.674647, -1.72492, -1.768385, -1.804872, 
    -1.834236, -1.85636, -1.871159, -1.878573, -1.878573, -1.871159, 
    -1.85636, -1.834236, -1.804872, -1.768385, -1.72492, -1.674647, 
    -1.617765, -1.554498, -1.485096, -1.409834, -1.329007, -1.242936, 
    -1.151959, -1.056436, -0.9567434, -0.8532751, -0.7464395, -0.6366579, 
    -0.5243638, -0.4100002, -0.2940186, -0.1768766, -0.05903652,
  // z(11, 0-99)
    0.0639366, 0.1915575, 0.3184223, 0.4440306, 0.5678864, 0.689501, 
    0.8083946, 0.9240977, 1.036154, 1.144121, 1.247572, 1.3461, 1.439316, 
    1.526851, 1.608361, 1.683522, 1.75204, 1.813644, 1.86809, 1.915163, 
    1.954678, 1.986479, 2.01044, 2.026466, 2.034496, 2.034496, 2.026466, 
    2.01044, 1.986479, 1.954678, 1.915163, 1.86809, 1.813644, 1.75204, 
    1.683522, 1.608361, 1.526851, 1.439316, 1.3461, 1.247572, 1.144121, 
    1.036154, 0.9240977, 0.8083946, 0.689501, 0.5678864, 0.4440306, 
    0.3184223, 0.1915575, 0.0639366, -0.0639366, -0.1915575, -0.3184223, 
    -0.4440306, -0.5678864, -0.689501, -0.8083946, -0.9240977, -1.036154, 
    -1.144121, -1.247572, -1.3461, -1.439316, -1.526851, -1.608361, 
    -1.683522, -1.75204, -1.813644, -1.86809, -1.915163, -1.954678, 
    -1.986479, -2.01044, -2.026466, -2.034496, -2.034496, -2.026466, 
    -2.01044, -1.986479, -1.954678, -1.915163, -1.86809, -1.813644, -1.75204, 
    -1.683522, -1.608361, -1.526851, -1.439316, -1.3461, -1.247572, 
    -1.144121, -1.036154, -0.9240977, -0.8083946, -0.689501, -0.5678864, 
    -0.4440306, -0.3184223, -0.1915575, -0.0639366,
  // z(12, 0-99)
    0.06871103, 0.2058619, 0.3422004, 0.4771883, 0.610293, 0.7409892, 
    0.868761, 0.9931042, 1.113528, 1.229557, 1.340734, 1.44662, 1.546796, 
    1.640868, 1.728464, 1.809239, 1.882873, 1.949077, 2.007588, 2.058177, 
    2.100642, 2.134818, 2.160568, 2.177792, 2.186421, 2.186421, 2.177792, 
    2.160568, 2.134818, 2.100642, 2.058177, 2.007588, 1.949077, 1.882873, 
    1.809239, 1.728464, 1.640868, 1.546796, 1.44662, 1.340734, 1.229557, 
    1.113528, 0.9931042, 0.868761, 0.7409892, 0.610293, 0.4771883, 0.3422004, 
    0.2058619, 0.06871103, -0.06871103, -0.2058619, -0.3422004, -0.4771883, 
    -0.610293, -0.7409892, -0.868761, -0.9931042, -1.113528, -1.229557, 
    -1.340734, -1.44662, -1.546796, -1.640868, -1.728464, -1.809239, 
    -1.882873, -1.949077, -2.007588, -2.058177, -2.100642, -2.134818, 
    -2.160568, -2.177792, -2.186421, -2.186421, -2.177792, -2.160568, 
    -2.134818, -2.100642, -2.058177, -2.007588, -1.949077, -1.882873, 
    -1.809239, -1.728464, -1.640868, -1.546796, -1.44662, -1.340734, 
    -1.229557, -1.113528, -0.9931042, -0.868761, -0.7409892, -0.610293, 
    -0.4771883, -0.3422004, -0.2058619, -0.06871103,
  // z(13, 0-99)
    0.07335982, 0.21979, 0.3653527, 0.5094736, 0.6515837, 0.7911224, 
    0.9275389, 1.060295, 1.188866, 1.312746, 1.431444, 1.544494, 1.651448, 
    1.751884, 1.845407, 1.931647, 2.010263, 2.080946, 2.143416, 2.197427, 
    2.242766, 2.279253, 2.306746, 2.325135, 2.334347, 2.334347, 2.325135, 
    2.306746, 2.279253, 2.242766, 2.197427, 2.143416, 2.080946, 2.010263, 
    1.931647, 1.845407, 1.751884, 1.651448, 1.544494, 1.431444, 1.312746, 
    1.188866, 1.060295, 0.9275389, 0.7911224, 0.6515837, 0.5094736, 
    0.3653527, 0.21979, 0.07335982, -0.07335982, -0.21979, -0.3653527, 
    -0.5094736, -0.6515837, -0.7911224, -0.9275389, -1.060295, -1.188866, 
    -1.312746, -1.431444, -1.544494, -1.651448, -1.751884, -1.845407, 
    -1.931647, -2.010263, -2.080946, -2.143416, -2.197427, -2.242766, 
    -2.279253, -2.306746, -2.325135, -2.334347, -2.334347, -2.325135, 
    -2.306746, -2.279253, -2.242766, -2.197427, -2.143416, -2.080946, 
    -2.010263, -1.931647, -1.845407, -1.751884, -1.651448, -1.544494, 
    -1.431444, -1.312746, -1.188866, -1.060295, -0.9275389, -0.7911224, 
    -0.6515837, -0.5094736, -0.3653527, -0.21979, -0.07335982,
  // z(14, 0-99)
    0.07788298, 0.2333416, 0.3878793, 0.5408862, 0.6917585, 0.8399007, 
    0.9847282, 1.125669, 1.262168, 1.393686, 1.519703, 1.639723, 1.753271, 
    1.8599, 1.959189, 2.050746, 2.13421, 2.209251, 2.275573, 2.332914, 
    2.381048, 2.419785, 2.448973, 2.468496, 2.478276, 2.478276, 2.468496, 
    2.448973, 2.419785, 2.381048, 2.332914, 2.275573, 2.209251, 2.13421, 
    2.050746, 1.959189, 1.8599, 1.753271, 1.639723, 1.519703, 1.393686, 
    1.262168, 1.125669, 0.9847282, 0.8399007, 0.6917585, 0.5408862, 
    0.3878793, 0.2333416, 0.07788298, -0.07788298, -0.2333416, -0.3878793, 
    -0.5408862, -0.6917585, -0.8399007, -0.9847282, -1.125669, -1.262168, 
    -1.393686, -1.519703, -1.639723, -1.753271, -1.8599, -1.959189, 
    -2.050746, -2.13421, -2.209251, -2.275573, -2.332914, -2.381048, 
    -2.419785, -2.448973, -2.468496, -2.478276, -2.478276, -2.468496, 
    -2.448973, -2.419785, -2.381048, -2.332914, -2.275573, -2.209251, 
    -2.13421, -2.050746, -1.959189, -1.8599, -1.753271, -1.639723, -1.519703, 
    -1.393686, -1.262168, -1.125669, -0.9847282, -0.8399007, -0.6917585, 
    -0.5408862, -0.3878793, -0.2333416, -0.07788298,
  // z(15, 0-99)
    0.08228049, 0.2465167, 0.4097801, 0.5714262, 0.7308172, 0.887324, 
    1.040329, 1.189228, 1.333434, 1.472377, 1.60551, 1.732306, 1.852266, 
    1.964916, 2.069811, 2.166538, 2.254714, 2.333992, 2.404058, 2.464637, 
    2.515489, 2.556414, 2.58725, 2.607875, 2.618207, 2.618207, 2.607875, 
    2.58725, 2.556414, 2.515489, 2.464637, 2.404058, 2.333992, 2.254714, 
    2.166538, 2.069811, 1.964916, 1.852266, 1.732306, 1.60551, 1.472377, 
    1.333434, 1.189228, 1.040329, 0.887324, 0.7308172, 0.5714262, 0.4097801, 
    0.2465167, 0.08228049, -0.08228049, -0.2465167, -0.4097801, -0.5714262, 
    -0.7308172, -0.887324, -1.040329, -1.189228, -1.333434, -1.472377, 
    -1.60551, -1.732306, -1.852266, -1.964916, -2.069811, -2.166538, 
    -2.254714, -2.333992, -2.404058, -2.464637, -2.515489, -2.556414, 
    -2.58725, -2.607875, -2.618207, -2.618207, -2.607875, -2.58725, 
    -2.556414, -2.515489, -2.464637, -2.404058, -2.333992, -2.254714, 
    -2.166538, -2.069811, -1.964916, -1.852266, -1.732306, -1.60551, 
    -1.472377, -1.333434, -1.189228, -1.040329, -0.887324, -0.7308172, 
    -0.5714262, -0.4097801, -0.2465167, -0.08228049,
  // z(16, 0-99)
    0.08655234, 0.2593155, 0.4310552, 0.6010937, 0.76876, 0.9333923, 
    1.094341, 1.250971, 1.402664, 1.548821, 1.688865, 1.822245, 1.948433, 
    2.066931, 2.177272, 2.279021, 2.371775, 2.455168, 2.528873, 2.592597, 
    2.646089, 2.689139, 2.721575, 2.743271, 2.75414, 2.75414, 2.743271, 
    2.721575, 2.689139, 2.646089, 2.592597, 2.528873, 2.455168, 2.371775, 
    2.279021, 2.177272, 2.066931, 1.948433, 1.822245, 1.688865, 1.548821, 
    1.402664, 1.250971, 1.094341, 0.9333923, 0.76876, 0.6010937, 0.4310552, 
    0.2593155, 0.08655234, -0.08655234, -0.2593155, -0.4310552, -0.6010937, 
    -0.76876, -0.9333923, -1.094341, -1.250971, -1.402664, -1.548821, 
    -1.688865, -1.822245, -1.948433, -2.066931, -2.177272, -2.279021, 
    -2.371775, -2.455168, -2.528873, -2.592597, -2.646089, -2.689139, 
    -2.721575, -2.743271, -2.75414, -2.75414, -2.743271, -2.721575, 
    -2.689139, -2.646089, -2.592597, -2.528873, -2.455168, -2.371775, 
    -2.279021, -2.177272, -2.066931, -1.948433, -1.822245, -1.688865, 
    -1.548821, -1.402664, -1.250971, -1.094341, -0.9333923, -0.76876, 
    -0.6010937, -0.4310552, -0.2593155, -0.08655234,
  // z(17, 0-99)
    0.09069857, 0.2717378, 0.4517045, 0.6298886, 0.8055868, 0.9781057, 
    1.146765, 1.310898, 1.469857, 1.623016, 1.769769, 1.909538, 2.041771, 
    2.165946, 2.281573, 2.388195, 2.485393, 2.572781, 2.650017, 2.716793, 
    2.772848, 2.81796, 2.85195, 2.874685, 2.886075, 2.886075, 2.874685, 
    2.85195, 2.81796, 2.772848, 2.716793, 2.650017, 2.572781, 2.485393, 
    2.388195, 2.281573, 2.165946, 2.041771, 1.909538, 1.769769, 1.623016, 
    1.469857, 1.310898, 1.146765, 0.9781057, 0.8055868, 0.6298886, 0.4517045, 
    0.2717378, 0.09069857, -0.09069857, -0.2717378, -0.4517045, -0.6298886, 
    -0.8055868, -0.9781057, -1.146765, -1.310898, -1.469857, -1.623016, 
    -1.769769, -1.909538, -2.041771, -2.165946, -2.281573, -2.388195, 
    -2.485393, -2.572781, -2.650017, -2.716793, -2.772848, -2.81796, 
    -2.85195, -2.874685, -2.886075, -2.886075, -2.874685, -2.85195, -2.81796, 
    -2.772848, -2.716793, -2.650017, -2.572781, -2.485393, -2.388195, 
    -2.281573, -2.165946, -2.041771, -1.909538, -1.769769, -1.623016, 
    -1.469857, -1.310898, -1.146765, -0.9781057, -0.8055868, -0.6298886, 
    -0.4517045, -0.2717378, -0.09069857,
  // z(18, 0-99)
    0.09471914, 0.2837836, 0.4717281, 0.6578109, 0.8412977, 1.021464, 
    1.197599, 1.369008, 1.535014, 1.694962, 1.848221, 1.994186, 2.132281, 
    2.26196, 2.382712, 2.494061, 2.595567, 2.68683, 2.767489, 2.837226, 
    2.895766, 2.942877, 2.978374, 3.002117, 3.014012, 3.014012, 3.002117, 
    2.978374, 2.942877, 2.895766, 2.837226, 2.767489, 2.68683, 2.595567, 
    2.494061, 2.382712, 2.26196, 2.132281, 1.994186, 1.848221, 1.694962, 
    1.535014, 1.369008, 1.197599, 1.021464, 0.8412977, 0.6578109, 0.4717281, 
    0.2837836, 0.09471914, -0.09471914, -0.2837836, -0.4717281, -0.6578109, 
    -0.8412977, -1.021464, -1.197599, -1.369008, -1.535014, -1.694962, 
    -1.848221, -1.994186, -2.132281, -2.26196, -2.382712, -2.494061, 
    -2.595567, -2.68683, -2.767489, -2.837226, -2.895766, -2.942877, 
    -2.978374, -3.002117, -3.014012, -3.014012, -3.002117, -2.978374, 
    -2.942877, -2.895766, -2.837226, -2.767489, -2.68683, -2.595567, 
    -2.494061, -2.382712, -2.26196, -2.132281, -1.994186, -1.848221, 
    -1.694962, -1.535014, -1.369008, -1.197599, -1.021464, -0.8412977, 
    -0.6578109, -0.4717281, -0.2837836, -0.09471914,
  // z(19, 0-99)
    0.09861408, 0.295453, 0.491126, 0.6848607, 0.8758926, 1.063468, 1.246846, 
    1.425303, 1.598135, 1.764661, 1.924222, 2.076189, 2.219962, 2.354974, 
    2.480692, 2.596619, 2.7023, 2.797315, 2.881291, 2.953895, 3.014842, 
    3.063891, 3.100847, 3.125567, 3.137951, 3.137951, 3.125567, 3.100847, 
    3.063891, 3.014842, 2.953895, 2.881291, 2.797315, 2.7023, 2.596619, 
    2.480692, 2.354974, 2.219962, 2.076189, 1.924222, 1.764661, 1.598135, 
    1.425303, 1.246846, 1.063468, 0.8758926, 0.6848607, 0.491126, 0.295453, 
    0.09861408, -0.09861408, -0.295453, -0.491126, -0.6848607, -0.8758926, 
    -1.063468, -1.246846, -1.425303, -1.598135, -1.764661, -1.924222, 
    -2.076189, -2.219962, -2.354974, -2.480692, -2.596619, -2.7023, 
    -2.797315, -2.881291, -2.953895, -3.014842, -3.063891, -3.100847, 
    -3.125567, -3.137951, -3.137951, -3.125567, -3.100847, -3.063891, 
    -3.014842, -2.953895, -2.881291, -2.797315, -2.7023, -2.596619, 
    -2.480692, -2.354974, -2.219962, -2.076189, -1.924222, -1.764661, 
    -1.598135, -1.425303, -1.246846, -1.063468, -0.8758926, -0.6848607, 
    -0.491126, -0.295453, -0.09861408,
  // z(20, 0-99)
    0.1023834, 0.306746, 0.5098981, 0.7110379, 0.9093715, 1.104116, 1.294504, 
    1.479782, 1.65922, 1.832111, 1.997771, 2.155546, 2.304815, 2.444987, 
    2.57551, 2.695869, 2.805589, 2.904236, 2.991421, 3.066801, 3.130077, 
    3.181001, 3.21937, 3.245034, 3.257892, 3.257892, 3.245034, 3.21937, 
    3.181001, 3.130077, 3.066801, 2.991421, 2.904236, 2.805589, 2.695869, 
    2.57551, 2.444987, 2.304815, 2.155546, 1.997771, 1.832111, 1.65922, 
    1.479782, 1.294504, 1.104116, 0.9093715, 0.7110379, 0.5098981, 0.306746, 
    0.1023834, -0.1023834, -0.306746, -0.5098981, -0.7110379, -0.9093715, 
    -1.104116, -1.294504, -1.479782, -1.65922, -1.832111, -1.997771, 
    -2.155546, -2.304815, -2.444987, -2.57551, -2.695869, -2.805589, 
    -2.904236, -2.991421, -3.066801, -3.130077, -3.181001, -3.21937, 
    -3.245034, -3.257892, -3.257892, -3.245034, -3.21937, -3.181001, 
    -3.130077, -3.066801, -2.991421, -2.904236, -2.805589, -2.695869, 
    -2.57551, -2.444987, -2.304815, -2.155546, -1.997771, -1.832111, 
    -1.65922, -1.479782, -1.294504, -1.104116, -0.9093715, -0.7110379, 
    -0.5098981, -0.306746, -0.1023834,
  // z(21, 0-99)
    0.106027, 0.3176626, 0.5280445, 0.7363425, 0.9417345, 1.14341, 1.340573, 
    1.532445, 1.718269, 1.897312, 2.068868, 2.232258, 2.386839, 2.532, 
    2.667168, 2.791811, 2.905435, 3.007592, 3.097881, 3.175943, 3.241471, 
    3.294207, 3.333942, 3.360519, 3.373834, 3.373834, 3.360519, 3.333942, 
    3.294207, 3.241471, 3.175943, 3.097881, 3.007592, 2.905435, 2.791811, 
    2.667168, 2.532, 2.386839, 2.232258, 2.068868, 1.897312, 1.718269, 
    1.532445, 1.340573, 1.14341, 0.9417345, 0.7363425, 0.5280445, 0.3176626, 
    0.106027, -0.106027, -0.3176626, -0.5280445, -0.7363425, -0.9417345, 
    -1.14341, -1.340573, -1.532445, -1.718269, -1.897312, -2.068868, 
    -2.232258, -2.386839, -2.532, -2.667168, -2.791811, -2.905435, -3.007592, 
    -3.097881, -3.175943, -3.241471, -3.294207, -3.333942, -3.360519, 
    -3.373834, -3.373834, -3.360519, -3.333942, -3.294207, -3.241471, 
    -3.175943, -3.097881, -3.007592, -2.905435, -2.791811, -2.667168, -2.532, 
    -2.386839, -2.232258, -2.068868, -1.897312, -1.718269, -1.532445, 
    -1.340573, -1.14341, -0.9417345, -0.7363425, -0.5280445, -0.3176626, 
    -0.106027,
  // z(22, 0-99)
    0.109545, 0.3282028, 0.5455652, 0.7607746, 0.9729815, 1.181348, 1.385053, 
    1.583292, 1.775282, 1.960266, 2.137513, 2.306325, 2.466035, 2.616012, 
    2.755666, 2.884444, 3.001838, 3.107385, 3.200669, 3.281322, 3.349024, 
    3.40351, 3.444563, 3.472022, 3.485779, 3.485779, 3.472022, 3.444563, 
    3.40351, 3.349024, 3.281322, 3.200669, 3.107385, 3.001838, 2.884444, 
    2.755666, 2.616012, 2.466035, 2.306325, 2.137513, 1.960266, 1.775282, 
    1.583292, 1.385053, 1.181348, 0.9729815, 0.7607746, 0.5455652, 0.3282028, 
    0.109545, -0.109545, -0.3282028, -0.5455652, -0.7607746, -0.9729815, 
    -1.181348, -1.385053, -1.583292, -1.775282, -1.960266, -2.137513, 
    -2.306325, -2.466035, -2.616012, -2.755666, -2.884444, -3.001838, 
    -3.107385, -3.200669, -3.281322, -3.349024, -3.40351, -3.444563, 
    -3.472022, -3.485779, -3.485779, -3.472022, -3.444563, -3.40351, 
    -3.349024, -3.281322, -3.200669, -3.107385, -3.001838, -2.884444, 
    -2.755666, -2.616012, -2.466035, -2.306325, -2.137513, -1.960266, 
    -1.775282, -1.583292, -1.385053, -1.181348, -0.9729815, -0.7607746, 
    -0.5455652, -0.3282028, -0.109545,
  // z(23, 0-99)
    0.1129374, 0.3383664, 0.5624601, 0.784334, 1.003113, 1.217932, 1.427945, 
    1.632323, 1.830258, 2.020971, 2.203707, 2.377747, 2.542403, 2.697024, 
    2.841002, 2.973768, 3.094798, 3.203614, 3.299787, 3.382937, 3.452736, 
    3.508909, 3.551234, 3.579543, 3.593726, 3.593726, 3.579543, 3.551234, 
    3.508909, 3.452736, 3.382937, 3.299787, 3.203614, 3.094798, 2.973768, 
    2.841002, 2.697024, 2.542403, 2.377747, 2.203707, 2.020971, 1.830258, 
    1.632323, 1.427945, 1.217932, 1.003113, 0.784334, 0.5624601, 0.3383664, 
    0.1129374, -0.1129374, -0.3383664, -0.5624601, -0.784334, -1.003113, 
    -1.217932, -1.427945, -1.632323, -1.830258, -2.020971, -2.203707, 
    -2.377747, -2.542403, -2.697024, -2.841002, -2.973768, -3.094798, 
    -3.203614, -3.299787, -3.382937, -3.452736, -3.508909, -3.551234, 
    -3.579543, -3.593726, -3.593726, -3.579543, -3.551234, -3.508909, 
    -3.452736, -3.382937, -3.299787, -3.203614, -3.094798, -2.973768, 
    -2.841002, -2.697024, -2.542403, -2.377747, -2.203707, -2.020971, 
    -1.830258, -1.632323, -1.427945, -1.217932, -1.003113, -0.784334, 
    -0.5624601, -0.3383664, -0.1129374,
  // z(24, 0-99)
    0.1162041, 0.3481537, 0.5787293, 0.8070209, 1.032128, 1.253161, 1.469249, 
    1.679538, 1.883199, 2.079427, 2.26745, 2.446523, 2.615942, 2.775036, 
    2.923178, 3.059785, 3.184315, 3.296279, 3.395233, 3.480788, 3.552607, 
    3.610404, 3.653953, 3.683081, 3.697675, 3.697675, 3.683081, 3.653953, 
    3.610404, 3.552607, 3.480788, 3.395233, 3.296279, 3.184315, 3.059785, 
    2.923178, 2.775036, 2.615942, 2.446523, 2.26745, 2.079427, 1.883199, 
    1.679538, 1.469249, 1.253161, 1.032128, 0.8070209, 0.5787293, 0.3481537, 
    0.1162041, -0.1162041, -0.3481537, -0.5787293, -0.8070209, -1.032128, 
    -1.253161, -1.469249, -1.679538, -1.883199, -2.079427, -2.26745, 
    -2.446523, -2.615942, -2.775036, -2.923178, -3.059785, -3.184315, 
    -3.296279, -3.395233, -3.480788, -3.552607, -3.610404, -3.653953, 
    -3.683081, -3.697675, -3.697675, -3.683081, -3.653953, -3.610404, 
    -3.552607, -3.480788, -3.395233, -3.296279, -3.184315, -3.059785, 
    -2.923178, -2.775036, -2.615942, -2.446523, -2.26745, -2.079427, 
    -1.883199, -1.679538, -1.469249, -1.253161, -1.032128, -0.8070209, 
    -0.5787293, -0.3481537, -0.1162041,
  // z(25, 0-99)
    0.1193452, 0.3575645, 0.5943727, 0.8288352, 1.060027, 1.287035, 1.508963, 
    1.724937, 1.934103, 2.135636, 2.32874, 2.512655, 2.686652, 2.850047, 
    3.002194, 3.142493, 3.270389, 3.385379, 3.487009, 3.574877, 3.648636, 
    3.707996, 3.752722, 3.782638, 3.797625, 3.797625, 3.782638, 3.752722, 
    3.707996, 3.648636, 3.574877, 3.487009, 3.385379, 3.270389, 3.142493, 
    3.002194, 2.850047, 2.686652, 2.512655, 2.32874, 2.135636, 1.934103, 
    1.724937, 1.508963, 1.287035, 1.060027, 0.8288352, 0.5943727, 0.3575645, 
    0.1193452, -0.1193452, -0.3575645, -0.5943727, -0.8288352, -1.060027, 
    -1.287035, -1.508963, -1.724937, -1.934103, -2.135636, -2.32874, 
    -2.512655, -2.686652, -2.850047, -3.002194, -3.142493, -3.270389, 
    -3.385379, -3.487009, -3.574877, -3.648636, -3.707996, -3.752722, 
    -3.782638, -3.797625, -3.797625, -3.782638, -3.752722, -3.707996, 
    -3.648636, -3.574877, -3.487009, -3.385379, -3.270389, -3.142493, 
    -3.002194, -2.850047, -2.686652, -2.512655, -2.32874, -2.135636, 
    -1.934103, -1.724937, -1.508963, -1.287035, -1.060027, -0.8288352, 
    -0.5943727, -0.3575645, -0.1193452,
  // z(26, 0-99)
    0.1223606, 0.3665989, 0.6093904, 0.849777, 1.08681, 1.319554, 1.54709, 
    1.76852, 1.982971, 2.189596, 2.387579, 2.57614, 2.754534, 2.922058, 
    3.078049, 3.221892, 3.353021, 3.470916, 3.575113, 3.665201, 3.740824, 
    3.801684, 3.84754, 3.878212, 3.893578, 3.893578, 3.878212, 3.84754, 
    3.801684, 3.740824, 3.665201, 3.575113, 3.470916, 3.353021, 3.221892, 
    3.078049, 2.922058, 2.754534, 2.57614, 2.387579, 2.189596, 1.982971, 
    1.76852, 1.54709, 1.319554, 1.08681, 0.849777, 0.6093904, 0.3665989, 
    0.1223606, -0.1223606, -0.3665989, -0.6093904, -0.849777, -1.08681, 
    -1.319554, -1.54709, -1.76852, -1.982971, -2.189596, -2.387579, -2.57614, 
    -2.754534, -2.922058, -3.078049, -3.221892, -3.353021, -3.470916, 
    -3.575113, -3.665201, -3.740824, -3.801684, -3.84754, -3.878212, 
    -3.893578, -3.893578, -3.878212, -3.84754, -3.801684, -3.740824, 
    -3.665201, -3.575113, -3.470916, -3.353021, -3.221892, -3.078049, 
    -2.922058, -2.754534, -2.57614, -2.387579, -2.189596, -1.982971, 
    -1.76852, -1.54709, -1.319554, -1.08681, -0.849777, -0.6093904, 
    -0.3665989, -0.1223606,
  // z(27, 0-99)
    0.1252504, 0.3752569, 0.6237825, 0.8698462, 1.112477, 1.350717, 1.583627, 
    1.810287, 2.029803, 2.241307, 2.443967, 2.636981, 2.819588, 2.991068, 
    3.150743, 3.297984, 3.432209, 3.552889, 3.659547, 3.751762, 3.829171, 
    3.891468, 3.938407, 3.969803, 3.985533, 3.985533, 3.969803, 3.938407, 
    3.891468, 3.829171, 3.751762, 3.659547, 3.552889, 3.432209, 3.297984, 
    3.150743, 2.991068, 2.819588, 2.636981, 2.443967, 2.241307, 2.029803, 
    1.810287, 1.583627, 1.350717, 1.112477, 0.8698462, 0.6237825, 0.3752569, 
    0.1252504, -0.1252504, -0.3752569, -0.6237825, -0.8698462, -1.112477, 
    -1.350717, -1.583627, -1.810287, -2.029803, -2.241307, -2.443967, 
    -2.636981, -2.819588, -2.991068, -3.150743, -3.297984, -3.432209, 
    -3.552889, -3.659547, -3.751762, -3.829171, -3.891468, -3.938407, 
    -3.969803, -3.985533, -3.985533, -3.969803, -3.938407, -3.891468, 
    -3.829171, -3.751762, -3.659547, -3.552889, -3.432209, -3.297984, 
    -3.150743, -2.991068, -2.819588, -2.636981, -2.443967, -2.241307, 
    -2.029803, -1.810287, -1.583627, -1.350717, -1.112477, -0.8698462, 
    -0.6237825, -0.3752569, -0.1252504,
  // z(28, 0-99)
    0.1280145, 0.3835384, 0.6375487, 0.8890428, 1.137028, 1.380526, 1.618576, 
    1.850238, 2.074598, 2.290771, 2.497903, 2.695177, 2.881814, 3.057078, 
    3.220277, 3.370767, 3.507954, 3.631297, 3.740309, 3.83456, 3.913677, 
    3.977349, 4.025324, 4.057413, 4.073489, 4.073489, 4.057413, 4.025324, 
    3.977349, 3.913677, 3.83456, 3.740309, 3.631297, 3.507954, 3.370767, 
    3.220277, 3.057078, 2.881814, 2.695177, 2.497903, 2.290771, 2.074598, 
    1.850238, 1.618576, 1.380526, 1.137028, 0.8890428, 0.6375487, 0.3835384, 
    0.1280145, -0.1280145, -0.3835384, -0.6375487, -0.8890428, -1.137028, 
    -1.380526, -1.618576, -1.850238, -2.074598, -2.290771, -2.497903, 
    -2.695177, -2.881814, -3.057078, -3.220277, -3.370767, -3.507954, 
    -3.631297, -3.740309, -3.83456, -3.913677, -3.977349, -4.025324, 
    -4.057413, -4.073489, -4.073489, -4.057413, -4.025324, -3.977349, 
    -3.913677, -3.83456, -3.740309, -3.631297, -3.507954, -3.370767, 
    -3.220277, -3.057078, -2.881814, -2.695177, -2.497903, -2.290771, 
    -2.074598, -1.850238, -1.618576, -1.380526, -1.137028, -0.8890428, 
    -0.6375487, -0.3835384, -0.1280145,
  // z(29, 0-99)
    0.1306531, 0.3914435, 0.6506892, 0.9073668, 1.160463, 1.40898, 1.651937, 
    1.888373, 2.117358, 2.337986, 2.549387, 2.750727, 2.941211, 3.120087, 
    3.28665, 3.440242, 3.580256, 3.706142, 3.8174, 3.913594, 3.994342, 
    4.059326, 4.10829, 4.14104, 4.157447, 4.157447, 4.14104, 4.10829, 
    4.059326, 3.994342, 3.913594, 3.8174, 3.706142, 3.580256, 3.440242, 
    3.28665, 3.120087, 2.941211, 2.750727, 2.549387, 2.337986, 2.117358, 
    1.888373, 1.651937, 1.40898, 1.160463, 0.9073668, 0.6506892, 0.3914435, 
    0.1306531, -0.1306531, -0.3914435, -0.6506892, -0.9073668, -1.160463, 
    -1.40898, -1.651937, -1.888373, -2.117358, -2.337986, -2.549387, 
    -2.750727, -2.941211, -3.120087, -3.28665, -3.440242, -3.580256, 
    -3.706142, -3.8174, -3.913594, -3.994342, -4.059326, -4.10829, -4.14104, 
    -4.157447, -4.157447, -4.14104, -4.10829, -4.059326, -3.994342, 
    -3.913594, -3.8174, -3.706142, -3.580256, -3.440242, -3.28665, -3.120087, 
    -2.941211, -2.750727, -2.549387, -2.337986, -2.117358, -1.888373, 
    -1.651937, -1.40898, -1.160463, -0.9073668, -0.6506892, -0.3914435, 
    -0.1306531,
  // z(30, 0-99)
    0.1331659, 0.3989722, 0.6632039, 0.9248183, 1.182783, 1.436079, 1.683708, 
    1.924693, 2.158081, 2.382952, 2.598419, 2.803632, 2.997779, 3.180096, 
    3.349862, 3.506408, 3.649116, 3.777422, 3.890821, 3.988864, 4.071165, 
    4.137399, 4.187304, 4.220685, 4.237408, 4.237408, 4.220685, 4.187304, 
    4.137399, 4.071165, 3.988864, 3.890821, 3.777422, 3.649116, 3.506408, 
    3.349862, 3.180096, 2.997779, 2.803632, 2.598419, 2.382952, 2.158081, 
    1.924693, 1.683708, 1.436079, 1.182783, 0.9248183, 0.6632039, 0.3989722, 
    0.1331659, -0.1331659, -0.3989722, -0.6632039, -0.9248183, -1.182783, 
    -1.436079, -1.683708, -1.924693, -2.158081, -2.382952, -2.598419, 
    -2.803632, -2.997779, -3.180096, -3.349862, -3.506408, -3.649116, 
    -3.777422, -3.890821, -3.988864, -4.071165, -4.137399, -4.187304, 
    -4.220685, -4.237408, -4.237408, -4.220685, -4.187304, -4.137399, 
    -4.071165, -3.988864, -3.890821, -3.777422, -3.649116, -3.506408, 
    -3.349862, -3.180096, -2.997779, -2.803632, -2.598419, -2.382952, 
    -2.158081, -1.924693, -1.683708, -1.436079, -1.182783, -0.9248183, 
    -0.6632039, -0.3989722, -0.1331659,
  // z(31, 0-99)
    0.1355531, 0.4061244, 0.6750929, 0.9413971, 1.203986, 1.461823, 1.713892, 
    1.959196, 2.196768, 2.425671, 2.645, 2.853891, 3.051519, 3.237104, 
    3.409914, 3.569266, 3.714532, 3.845139, 3.96057, 4.060371, 4.144147, 
    4.211569, 4.262369, 4.296348, 4.313371, 4.313371, 4.296348, 4.262369, 
    4.211569, 4.144147, 4.060371, 3.96057, 3.845139, 3.714532, 3.569266, 
    3.409914, 3.237104, 3.051519, 2.853891, 2.645, 2.425671, 2.196768, 
    1.959196, 1.713892, 1.461823, 1.203986, 0.9413971, 0.6750929, 0.4061244, 
    0.1355531, -0.1355531, -0.4061244, -0.6750929, -0.9413971, -1.203986, 
    -1.461823, -1.713892, -1.959196, -2.196768, -2.425671, -2.645, -2.853891, 
    -3.051519, -3.237104, -3.409914, -3.569266, -3.714532, -3.845139, 
    -3.96057, -4.060371, -4.144147, -4.211569, -4.262369, -4.296348, 
    -4.313371, -4.313371, -4.296348, -4.262369, -4.211569, -4.144147, 
    -4.060371, -3.96057, -3.845139, -3.714532, -3.569266, -3.409914, 
    -3.237104, -3.051519, -2.853891, -2.645, -2.425671, -2.196768, -1.959196, 
    -1.713892, -1.461823, -1.203986, -0.9413971, -0.6750929, -0.4061244, 
    -0.1355531,
  // z(32, 0-99)
    0.1378147, 0.4129002, 0.6863562, 0.9571035, 1.224074, 1.486213, 1.742486, 
    1.991883, 2.233419, 2.466141, 2.68913, 2.901506, 3.102431, 3.291112, 
    3.466805, 3.628816, 3.776506, 3.909291, 4.026649, 4.128114, 4.213289, 
    4.281835, 4.333483, 4.368028, 4.385335, 4.385335, 4.368028, 4.333483, 
    4.281835, 4.213289, 4.128114, 4.026649, 3.909291, 3.776506, 3.628816, 
    3.466805, 3.291112, 3.102431, 2.901506, 2.68913, 2.466141, 2.233419, 
    1.991883, 1.742486, 1.486213, 1.224074, 0.9571035, 0.6863562, 0.4129002, 
    0.1378147, -0.1378147, -0.4129002, -0.6863562, -0.9571035, -1.224074, 
    -1.486213, -1.742486, -1.991883, -2.233419, -2.466141, -2.68913, 
    -2.901506, -3.102431, -3.291112, -3.466805, -3.628816, -3.776506, 
    -3.909291, -4.026649, -4.128114, -4.213289, -4.281835, -4.333483, 
    -4.368028, -4.385335, -4.385335, -4.368028, -4.333483, -4.281835, 
    -4.213289, -4.128114, -4.026649, -3.909291, -3.776506, -3.628816, 
    -3.466805, -3.291112, -3.102431, -2.901506, -2.68913, -2.466141, 
    -2.233419, -1.991883, -1.742486, -1.486213, -1.224074, -0.9571035, 
    -0.6863562, -0.4129002, -0.1378147,
  // z(33, 0-99)
    0.1399506, 0.4192996, 0.6969938, 0.9719372, 1.243045, 1.509247, 1.769492, 
    2.022755, 2.268034, 2.504363, 2.730807, 2.946475, 3.150514, 3.34212, 
    3.520536, 3.685057, 3.835036, 3.96988, 4.089056, 4.192094, 4.278588, 
    4.348197, 4.400645, 4.435726, 4.453301, 4.453301, 4.435726, 4.400645, 
    4.348197, 4.278588, 4.192094, 4.089056, 3.96988, 3.835036, 3.685057, 
    3.520536, 3.34212, 3.150514, 2.946475, 2.730807, 2.504363, 2.268034, 
    2.022755, 1.769492, 1.509247, 1.243045, 0.9719372, 0.6969938, 0.4192996, 
    0.1399506, -0.1399506, -0.4192996, -0.6969938, -0.9719372, -1.243045, 
    -1.509247, -1.769492, -2.022755, -2.268034, -2.504363, -2.730807, 
    -2.946475, -3.150514, -3.34212, -3.520536, -3.685057, -3.835036, 
    -3.96988, -4.089056, -4.192094, -4.278588, -4.348197, -4.400645, 
    -4.435726, -4.453301, -4.453301, -4.435726, -4.400645, -4.348197, 
    -4.278588, -4.192094, -4.089056, -3.96988, -3.835036, -3.685057, 
    -3.520536, -3.34212, -3.150514, -2.946475, -2.730807, -2.504363, 
    -2.268034, -2.022755, -1.769492, -1.509247, -1.243045, -0.9719372, 
    -0.6969938, -0.4192996, -0.1399506,
  // z(34, 0-99)
    0.1419609, 0.4253225, 0.7070056, 0.9858984, 1.2609, 1.530926, 1.79491, 
    2.05181, 2.300613, 2.540336, 2.770033, 2.988799, 3.195769, 3.390127, 
    3.571105, 3.737991, 3.890124, 4.026904, 4.147792, 4.252311, 4.340047, 
    4.410656, 4.463858, 4.499442, 4.51727, 4.51727, 4.499442, 4.463858, 
    4.410656, 4.340047, 4.252311, 4.147792, 4.026904, 3.890124, 3.737991, 
    3.571105, 3.390127, 3.195769, 2.988799, 2.770033, 2.540336, 2.300613, 
    2.05181, 1.79491, 1.530926, 1.2609, 0.9858984, 0.7070056, 0.4253225, 
    0.1419609, -0.1419609, -0.4253225, -0.7070056, -0.9858984, -1.2609, 
    -1.530926, -1.79491, -2.05181, -2.300613, -2.540336, -2.770033, 
    -2.988799, -3.195769, -3.390127, -3.571105, -3.737991, -3.890124, 
    -4.026904, -4.147792, -4.252311, -4.340047, -4.410656, -4.463858, 
    -4.499442, -4.51727, -4.51727, -4.499442, -4.463858, -4.410656, 
    -4.340047, -4.252311, -4.147792, -4.026904, -3.890124, -3.737991, 
    -3.571105, -3.390127, -3.195769, -2.988799, -2.770033, -2.540336, 
    -2.300613, -2.05181, -1.79491, -1.530926, -1.2609, -0.9858984, 
    -0.7070056, -0.4253225, -0.1419609,
  // z(35, 0-99)
    0.1438456, 0.430969, 0.7163916, 0.998987, 1.27764, 1.55125, 1.818739, 
    2.07905, 2.331155, 2.574061, 2.806808, 3.028478, 3.238195, 3.435134, 
    3.618515, 3.787616, 3.941768, 4.080364, 4.202857, 4.308764, 4.397665, 
    4.469211, 4.523119, 4.559176, 4.57724, 4.57724, 4.559176, 4.523119, 
    4.469211, 4.397665, 4.308764, 4.202857, 4.080364, 3.941768, 3.787616, 
    3.618515, 3.435134, 3.238195, 3.028478, 2.806808, 2.574061, 2.331155, 
    2.07905, 1.818739, 1.55125, 1.27764, 0.998987, 0.7163916, 0.430969, 
    0.1438456, -0.1438456, -0.430969, -0.7163916, -0.998987, -1.27764, 
    -1.55125, -1.818739, -2.07905, -2.331155, -2.574061, -2.806808, 
    -3.028478, -3.238195, -3.435134, -3.618515, -3.787616, -3.941768, 
    -4.080364, -4.202857, -4.308764, -4.397665, -4.469211, -4.523119, 
    -4.559176, -4.57724, -4.57724, -4.559176, -4.523119, -4.469211, 
    -4.397665, -4.308764, -4.202857, -4.080364, -3.941768, -3.787616, 
    -3.618515, -3.435134, -3.238195, -3.028478, -2.806808, -2.574061, 
    -2.331155, -2.07905, -1.818739, -1.55125, -1.27764, -0.998987, 
    -0.7163916, -0.430969, -0.1438456,
  // z(36, 0-99)
    0.1456046, 0.4362391, 0.725152, 1.011203, 1.293263, 1.57022, 1.840979, 
    2.104473, 2.359662, 2.605537, 2.841131, 3.065511, 3.277793, 3.47714, 
    3.662764, 3.833932, 3.98997, 4.130261, 4.254251, 4.361453, 4.451441, 
    4.523862, 4.578429, 4.614927, 4.633213, 4.633213, 4.614927, 4.578429, 
    4.523862, 4.451441, 4.361453, 4.254251, 4.130261, 3.98997, 3.833932, 
    3.662764, 3.47714, 3.277793, 3.065511, 2.841131, 2.605537, 2.359662, 
    2.104473, 1.840979, 1.57022, 1.293263, 1.011203, 0.725152, 0.4362391, 
    0.1456046, -0.1456046, -0.4362391, -0.725152, -1.011203, -1.293263, 
    -1.57022, -1.840979, -2.104473, -2.359662, -2.605537, -2.841131, 
    -3.065511, -3.277793, -3.47714, -3.662764, -3.833932, -3.98997, 
    -4.130261, -4.254251, -4.361453, -4.451441, -4.523862, -4.578429, 
    -4.614927, -4.633213, -4.633213, -4.614927, -4.578429, -4.523862, 
    -4.451441, -4.361453, -4.254251, -4.130261, -3.98997, -3.833932, 
    -3.662764, -3.47714, -3.277793, -3.065511, -2.841131, -2.605537, 
    -2.359662, -2.104473, -1.840979, -1.57022, -1.293263, -1.011203, 
    -0.725152, -0.4362391, -0.1456046,
  // z(37, 0-99)
    0.1472379, 0.4411327, 0.7332866, 1.022546, 1.307771, 1.587834, 1.861631, 
    2.12808, 2.386132, 2.634766, 2.873002, 3.099899, 3.314563, 3.516146, 
    3.703852, 3.87694, 4.034728, 4.176593, 4.301975, 4.410378, 4.501377, 
    4.57461, 4.629789, 4.666697, 4.685187, 4.685187, 4.666697, 4.629789, 
    4.57461, 4.501377, 4.410378, 4.301975, 4.176593, 4.034728, 3.87694, 
    3.703852, 3.516146, 3.314563, 3.099899, 2.873002, 2.634766, 2.386132, 
    2.12808, 1.861631, 1.587834, 1.307771, 1.022546, 0.7332866, 0.4411327, 
    0.1472379, -0.1472379, -0.4411327, -0.7332866, -1.022546, -1.307771, 
    -1.587834, -1.861631, -2.12808, -2.386132, -2.634766, -2.873002, 
    -3.099899, -3.314563, -3.516146, -3.703852, -3.87694, -4.034728, 
    -4.176593, -4.301975, -4.410378, -4.501377, -4.57461, -4.629789, 
    -4.666697, -4.685187, -4.685187, -4.666697, -4.629789, -4.57461, 
    -4.501377, -4.410378, -4.301975, -4.176593, -4.034728, -3.87694, 
    -3.703852, -3.516146, -3.314563, -3.099899, -2.873002, -2.634766, 
    -2.386132, -2.12808, -1.861631, -1.587834, -1.307771, -1.022546, 
    -0.7332866, -0.4411327, -0.1472379,
  // z(38, 0-99)
    0.1487457, 0.4456499, 0.7407954, 1.033017, 1.321162, 1.604093, 1.880694, 
    2.149872, 2.410566, 2.661746, 2.902421, 3.131642, 3.348504, 3.552151, 
    3.741779, 3.91664, 4.076044, 4.219361, 4.346027, 4.455541, 4.547471, 
    4.621454, 4.677198, 4.714484, 4.733163, 4.733163, 4.714484, 4.677198, 
    4.621454, 4.547471, 4.455541, 4.346027, 4.219361, 4.076044, 3.91664, 
    3.741779, 3.552151, 3.348504, 3.131642, 2.902421, 2.661746, 2.410566, 
    2.149872, 1.880694, 1.604093, 1.321162, 1.033017, 0.7407954, 0.4456499, 
    0.1487457, -0.1487457, -0.4456499, -0.7407954, -1.033017, -1.321162, 
    -1.604093, -1.880694, -2.149872, -2.410566, -2.661746, -2.902421, 
    -3.131642, -3.348504, -3.552151, -3.741779, -3.91664, -4.076044, 
    -4.219361, -4.346027, -4.455541, -4.547471, -4.621454, -4.677198, 
    -4.714484, -4.733163, -4.733163, -4.714484, -4.677198, -4.621454, 
    -4.547471, -4.455541, -4.346027, -4.219361, -4.076044, -3.91664, 
    -3.741779, -3.552151, -3.348504, -3.131642, -2.902421, -2.661746, 
    -2.410566, -2.149872, -1.880694, -1.604093, -1.321162, -1.033017, 
    -0.7407954, -0.4456499, -0.1487457,
  // z(39, 0-99)
    0.1501277, 0.4497907, 0.7476785, 1.042616, 1.333438, 1.618998, 1.898168, 
    2.169847, 2.432963, 2.686477, 2.929389, 3.16074, 3.379617, 3.585156, 
    3.776546, 3.953032, 4.113916, 4.258566, 4.386408, 4.49694, 4.589724, 
    4.664394, 4.720656, 4.758288, 4.777142, 4.777142, 4.758288, 4.720656, 
    4.664394, 4.589724, 4.49694, 4.386408, 4.258566, 4.113916, 3.953032, 
    3.776546, 3.585156, 3.379617, 3.16074, 2.929389, 2.686477, 2.432963, 
    2.169847, 1.898168, 1.618998, 1.333438, 1.042616, 0.7476785, 0.4497907, 
    0.1501277, -0.1501277, -0.4497907, -0.7476785, -1.042616, -1.333438, 
    -1.618998, -1.898168, -2.169847, -2.432963, -2.686477, -2.929389, 
    -3.16074, -3.379617, -3.585156, -3.776546, -3.953032, -4.113916, 
    -4.258566, -4.386408, -4.49694, -4.589724, -4.664394, -4.720656, 
    -4.758288, -4.777142, -4.777142, -4.758288, -4.720656, -4.664394, 
    -4.589724, -4.49694, -4.386408, -4.258566, -4.113916, -3.953032, 
    -3.776546, -3.585156, -3.379617, -3.16074, -2.929389, -2.686477, 
    -2.432963, -2.169847, -1.898168, -1.618998, -1.333438, -1.042616, 
    -0.7476785, -0.4497907, -0.1501277,
  // z(40, 0-99)
    0.1513842, 0.453555, 0.7539359, 1.051341, 1.344598, 1.632547, 1.914054, 
    2.188007, 2.453325, 2.708961, 2.953906, 3.187192, 3.407901, 3.61516, 
    3.808152, 3.986115, 4.148346, 4.294206, 4.423119, 4.534575, 4.628135, 
    4.703431, 4.760164, 4.798111, 4.817122, 4.817122, 4.798111, 4.760164, 
    4.703431, 4.628135, 4.534575, 4.423119, 4.294206, 4.148346, 3.986115, 
    3.808152, 3.61516, 3.407901, 3.187192, 2.953906, 2.708961, 2.453325, 
    2.188007, 1.914054, 1.632547, 1.344598, 1.051341, 0.7539359, 0.453555, 
    0.1513842, -0.1513842, -0.453555, -0.7539359, -1.051341, -1.344598, 
    -1.632547, -1.914054, -2.188007, -2.453325, -2.708961, -2.953906, 
    -3.187192, -3.407901, -3.61516, -3.808152, -3.986115, -4.148346, 
    -4.294206, -4.423119, -4.534575, -4.628135, -4.703431, -4.760164, 
    -4.798111, -4.817122, -4.817122, -4.798111, -4.760164, -4.703431, 
    -4.628135, -4.534575, -4.423119, -4.294206, -4.148346, -3.986115, 
    -3.808152, -3.61516, -3.407901, -3.187192, -2.953906, -2.708961, 
    -2.453325, -2.188007, -1.914054, -1.632547, -1.344598, -1.051341, 
    -0.7539359, -0.453555, -0.1513842,
  // z(41, 0-99)
    0.1525149, 0.4569429, 0.7595676, 1.059195, 1.354641, 1.644742, 1.928352, 
    2.204351, 2.471651, 2.729196, 2.97597, 3.211, 3.433357, 3.642164, 
    3.836598, 4.01589, 4.179333, 4.326282, 4.456158, 4.568447, 4.662706, 
    4.738564, 4.795721, 4.833951, 4.853104, 4.853104, 4.833951, 4.795721, 
    4.738564, 4.662706, 4.568447, 4.456158, 4.326282, 4.179333, 4.01589, 
    3.836598, 3.642164, 3.433357, 3.211, 2.97597, 2.729196, 2.471651, 
    2.204351, 1.928352, 1.644742, 1.354641, 1.059195, 0.7595676, 0.4569429, 
    0.1525149, -0.1525149, -0.4569429, -0.7595676, -1.059195, -1.354641, 
    -1.644742, -1.928352, -2.204351, -2.471651, -2.729196, -2.97597, -3.211, 
    -3.433357, -3.642164, -3.836598, -4.01589, -4.179333, -4.326282, 
    -4.456158, -4.568447, -4.662706, -4.738564, -4.795721, -4.833951, 
    -4.853104, -4.853104, -4.833951, -4.795721, -4.738564, -4.662706, 
    -4.568447, -4.456158, -4.326282, -4.179333, -4.01589, -3.836598, 
    -3.642164, -3.433357, -3.211, -2.97597, -2.729196, -2.471651, -2.204351, 
    -1.928352, -1.644742, -1.354641, -1.059195, -0.7595676, -0.4569429, 
    -0.1525149,
  // z(42, 0-99)
    0.1535201, 0.4599544, 0.7645735, 1.066175, 1.363569, 1.655582, 1.94106, 
    2.218879, 2.48794, 2.747183, 2.995583, 3.232162, 3.455984, 3.666168, 
    3.861883, 4.042356, 4.206877, 4.354795, 4.485526, 4.598555, 4.693435, 
    4.769793, 4.827327, 4.865809, 4.885088, 4.885088, 4.865809, 4.827327, 
    4.769793, 4.693435, 4.598555, 4.485526, 4.354795, 4.206877, 4.042356, 
    3.861883, 3.666168, 3.455984, 3.232162, 2.995583, 2.747183, 2.48794, 
    2.218879, 1.94106, 1.655582, 1.363569, 1.066175, 0.7645735, 0.4599544, 
    0.1535201, -0.1535201, -0.4599544, -0.7645735, -1.066175, -1.363569, 
    -1.655582, -1.94106, -2.218879, -2.48794, -2.747183, -2.995583, 
    -3.232162, -3.455984, -3.666168, -3.861883, -4.042356, -4.206877, 
    -4.354795, -4.485526, -4.598555, -4.693435, -4.769793, -4.827327, 
    -4.865809, -4.885088, -4.885088, -4.865809, -4.827327, -4.769793, 
    -4.693435, -4.598555, -4.485526, -4.354795, -4.206877, -4.042356, 
    -3.861883, -3.666168, -3.455984, -3.232162, -2.995583, -2.747183, 
    -2.48794, -2.218879, -1.94106, -1.655582, -1.363569, -1.066175, 
    -0.7645735, -0.4599544, -0.1535201,
  // z(43, 0-99)
    0.1543996, 0.4625894, 0.7689536, 1.072283, 1.371381, 1.665066, 1.952181, 
    2.23159, 2.502193, 2.762921, 3.012745, 3.250679, 3.475783, 3.687171, 
    3.884007, 4.065515, 4.230978, 4.379743, 4.511223, 4.624899, 4.720324, 
    4.797119, 4.854982, 4.893685, 4.913074, 4.913074, 4.893685, 4.854982, 
    4.797119, 4.720324, 4.624899, 4.511223, 4.379743, 4.230978, 4.065515, 
    3.884007, 3.687171, 3.475783, 3.250679, 3.012745, 2.762921, 2.502193, 
    2.23159, 1.952181, 1.665066, 1.371381, 1.072283, 0.7689536, 0.4625894, 
    0.1543996, -0.1543996, -0.4625894, -0.7689536, -1.072283, -1.371381, 
    -1.665066, -1.952181, -2.23159, -2.502193, -2.762921, -3.012745, 
    -3.250679, -3.475783, -3.687171, -3.884007, -4.065515, -4.230978, 
    -4.379743, -4.511223, -4.624899, -4.720324, -4.797119, -4.854982, 
    -4.893685, -4.913074, -4.913074, -4.893685, -4.854982, -4.797119, 
    -4.720324, -4.624899, -4.511223, -4.379743, -4.230978, -4.065515, 
    -3.884007, -3.687171, -3.475783, -3.250679, -3.012745, -2.762921, 
    -2.502193, -2.23159, -1.952181, -1.665066, -1.371381, -1.072283, 
    -0.7689536, -0.4625894, -0.1543996,
  // z(44, 0-99)
    0.1551534, 0.464848, 0.7727081, 1.077519, 1.378077, 1.673196, 1.961712, 
    2.242486, 2.51441, 2.776411, 3.027454, 3.26655, 3.492754, 3.705174, 
    3.902971, 4.085364, 4.251635, 4.401127, 4.533249, 4.64748, 4.743371, 
    4.820541, 4.878686, 4.917578, 4.937063, 4.937063, 4.917578, 4.878686, 
    4.820541, 4.743371, 4.64748, 4.533249, 4.401127, 4.251635, 4.085364, 
    3.902971, 3.705174, 3.492754, 3.26655, 3.027454, 2.776411, 2.51441, 
    2.242486, 1.961712, 1.673196, 1.378077, 1.077519, 0.7727081, 0.464848, 
    0.1551534, -0.1551534, -0.464848, -0.7727081, -1.077519, -1.378077, 
    -1.673196, -1.961712, -2.242486, -2.51441, -2.776411, -3.027454, 
    -3.26655, -3.492754, -3.705174, -3.902971, -4.085364, -4.251635, 
    -4.401127, -4.533249, -4.64748, -4.743371, -4.820541, -4.878686, 
    -4.917578, -4.937063, -4.937063, -4.917578, -4.878686, -4.820541, 
    -4.743371, -4.64748, -4.533249, -4.401127, -4.251635, -4.085364, 
    -3.902971, -3.705174, -3.492754, -3.26655, -3.027454, -2.776411, 
    -2.51441, -2.242486, -1.961712, -1.673196, -1.378077, -1.077519, 
    -0.7727081, -0.464848, -0.1551534,
  // z(45, 0-99)
    0.1557817, 0.4667302, 0.7758367, 1.081881, 1.383656, 1.679971, 1.969655, 
    2.251566, 2.524591, 2.787652, 3.039712, 3.279776, 3.506896, 3.720176, 
    3.918774, 4.101906, 4.26885, 4.418947, 4.551604, 4.666298, 4.762577, 
    4.840059, 4.89844, 4.93749, 4.957053, 4.957053, 4.93749, 4.89844, 
    4.840059, 4.762577, 4.666298, 4.551604, 4.418947, 4.26885, 4.101906, 
    3.918774, 3.720176, 3.506896, 3.279776, 3.039712, 2.787652, 2.524591, 
    2.251566, 1.969655, 1.679971, 1.383656, 1.081881, 0.7758367, 0.4667302, 
    0.1557817, -0.1557817, -0.4667302, -0.7758367, -1.081881, -1.383656, 
    -1.679971, -1.969655, -2.251566, -2.524591, -2.787652, -3.039712, 
    -3.279776, -3.506896, -3.720176, -3.918774, -4.101906, -4.26885, 
    -4.418947, -4.551604, -4.666298, -4.762577, -4.840059, -4.89844, 
    -4.93749, -4.957053, -4.957053, -4.93749, -4.89844, -4.840059, -4.762577, 
    -4.666298, -4.551604, -4.418947, -4.26885, -4.101906, -3.918774, 
    -3.720176, -3.506896, -3.279776, -3.039712, -2.787652, -2.524591, 
    -2.251566, -1.969655, -1.679971, -1.383656, -1.081881, -0.7758367, 
    -0.4667302, -0.1557817,
  // z(46, 0-99)
    0.1562842, 0.4682359, 0.7783397, 1.085372, 1.38812, 1.68539, 1.976009, 
    2.25883, 2.532736, 2.796646, 3.049519, 3.290357, 3.51821, 3.732178, 
    3.931416, 4.115139, 4.282622, 4.433203, 4.566288, 4.681352, 4.777941, 
    4.855674, 4.914243, 4.953419, 4.973045, 4.973045, 4.953419, 4.914243, 
    4.855674, 4.777941, 4.681352, 4.566288, 4.433203, 4.282622, 4.115139, 
    3.931416, 3.732178, 3.51821, 3.290357, 3.049519, 2.796646, 2.532736, 
    2.25883, 1.976009, 1.68539, 1.38812, 1.085372, 0.7783397, 0.4682359, 
    0.1562842, -0.1562842, -0.4682359, -0.7783397, -1.085372, -1.38812, 
    -1.68539, -1.976009, -2.25883, -2.532736, -2.796646, -3.049519, 
    -3.290357, -3.51821, -3.732178, -3.931416, -4.115139, -4.282622, 
    -4.433203, -4.566288, -4.681352, -4.777941, -4.855674, -4.914243, 
    -4.953419, -4.973045, -4.973045, -4.953419, -4.914243, -4.855674, 
    -4.777941, -4.681352, -4.566288, -4.433203, -4.282622, -4.115139, 
    -3.931416, -3.732178, -3.51821, -3.290357, -3.049519, -2.796646, 
    -2.532736, -2.25883, -1.976009, -1.68539, -1.38812, -1.085372, 
    -0.7783397, -0.4682359, -0.1562842,
  // z(47, 0-99)
    0.1566612, 0.4693652, 0.7802169, 1.087989, 1.391468, 1.689455, 1.980775, 
    2.264278, 2.538844, 2.803391, 3.056874, 3.298293, 3.526695, 3.741179, 
    3.940898, 4.125064, 4.292951, 4.443895, 4.577301, 4.692643, 4.789465, 
    4.867385, 4.926095, 4.965365, 4.985039, 4.985039, 4.965365, 4.926095, 
    4.867385, 4.789465, 4.692643, 4.577301, 4.443895, 4.292951, 4.125064, 
    3.940898, 3.741179, 3.526695, 3.298293, 3.056874, 2.803391, 2.538844, 
    2.264278, 1.980775, 1.689455, 1.391468, 1.087989, 0.7802169, 0.4693652, 
    0.1566612, -0.1566612, -0.4693652, -0.7802169, -1.087989, -1.391468, 
    -1.689455, -1.980775, -2.264278, -2.538844, -2.803391, -3.056874, 
    -3.298293, -3.526695, -3.741179, -3.940898, -4.125064, -4.292951, 
    -4.443895, -4.577301, -4.692643, -4.789465, -4.867385, -4.926095, 
    -4.965365, -4.985039, -4.985039, -4.965365, -4.926095, -4.867385, 
    -4.789465, -4.692643, -4.577301, -4.443895, -4.292951, -4.125064, 
    -3.940898, -3.741179, -3.526695, -3.298293, -3.056874, -2.803391, 
    -2.538844, -2.264278, -1.980775, -1.689455, -1.391468, -1.087989, 
    -0.7802169, -0.4693652, -0.1566612,
  // z(48, 0-99)
    0.1569124, 0.4701181, 0.7814684, 1.089735, 1.3937, 1.692165, 1.983952, 
    2.26791, 2.542916, 2.807888, 3.061777, 3.303583, 3.532352, 3.74718, 
    3.947219, 4.131681, 4.299837, 4.451023, 4.584643, 4.70017, 4.797147, 
    4.875192, 4.933997, 4.97333, 4.993035, 4.993035, 4.97333, 4.933997, 
    4.875192, 4.797147, 4.70017, 4.584643, 4.451023, 4.299837, 4.131681, 
    3.947219, 3.74718, 3.532352, 3.303583, 3.061777, 2.807888, 2.542916, 
    2.26791, 1.983952, 1.692165, 1.3937, 1.089735, 0.7814684, 0.4701181, 
    0.1569124, -0.1569124, -0.4701181, -0.7814684, -1.089735, -1.3937, 
    -1.692165, -1.983952, -2.26791, -2.542916, -2.807888, -3.061777, 
    -3.303583, -3.532352, -3.74718, -3.947219, -4.131681, -4.299837, 
    -4.451023, -4.584643, -4.70017, -4.797147, -4.875192, -4.933997, 
    -4.97333, -4.993035, -4.993035, -4.97333, -4.933997, -4.875192, 
    -4.797147, -4.70017, -4.584643, -4.451023, -4.299837, -4.131681, 
    -3.947219, -3.74718, -3.532352, -3.303583, -3.061777, -2.807888, 
    -2.542916, -2.26791, -1.983952, -1.692165, -1.3937, -1.089735, 
    -0.7814684, -0.4701181, -0.1569124,
  // z(49, 0-99)
    0.1570381, 0.4704945, 0.7820941, 1.090607, 1.394816, 1.69352, 1.985541, 
    2.269726, 2.544953, 2.810136, 3.064229, 3.306229, 3.53518, 3.75018, 
    3.95038, 4.134989, 4.30328, 4.454587, 4.588314, 4.703933, 4.800988, 
    4.879096, 4.937948, 4.977312, 4.997033, 4.997033, 4.977312, 4.937948, 
    4.879096, 4.800988, 4.703933, 4.588314, 4.454587, 4.30328, 4.134989, 
    3.95038, 3.75018, 3.53518, 3.306229, 3.064229, 2.810136, 2.544953, 
    2.269726, 1.985541, 1.69352, 1.394816, 1.090607, 0.7820941, 0.4704945, 
    0.1570381, -0.1570381, -0.4704945, -0.7820941, -1.090607, -1.394816, 
    -1.69352, -1.985541, -2.269726, -2.544953, -2.810136, -3.064229, 
    -3.306229, -3.53518, -3.75018, -3.95038, -4.134989, -4.30328, -4.454587, 
    -4.588314, -4.703933, -4.800988, -4.879096, -4.937948, -4.977312, 
    -4.997033, -4.997033, -4.977312, -4.937948, -4.879096, -4.800988, 
    -4.703933, -4.588314, -4.454587, -4.30328, -4.134989, -3.95038, -3.75018, 
    -3.53518, -3.306229, -3.064229, -2.810136, -2.544953, -2.269726, 
    -1.985541, -1.69352, -1.394816, -1.090607, -0.7820941, -0.4704945, 
    -0.1570381,
  // z(50, 0-99)
    0.1570381, 0.4704945, 0.7820941, 1.090607, 1.394816, 1.69352, 1.985541, 
    2.269726, 2.544953, 2.810136, 3.064229, 3.306229, 3.53518, 3.75018, 
    3.95038, 4.134989, 4.30328, 4.454587, 4.588314, 4.703933, 4.800988, 
    4.879096, 4.937948, 4.977312, 4.997033, 4.997033, 4.977312, 4.937948, 
    4.879096, 4.800988, 4.703933, 4.588314, 4.454587, 4.30328, 4.134989, 
    3.95038, 3.75018, 3.53518, 3.306229, 3.064229, 2.810136, 2.544953, 
    2.269726, 1.985541, 1.69352, 1.394816, 1.090607, 0.7820941, 0.4704945, 
    0.1570381, -0.1570381, -0.4704945, -0.7820941, -1.090607, -1.394816, 
    -1.69352, -1.985541, -2.269726, -2.544953, -2.810136, -3.064229, 
    -3.306229, -3.53518, -3.75018, -3.95038, -4.134989, -4.30328, -4.454587, 
    -4.588314, -4.703933, -4.800988, -4.879096, -4.937948, -4.977312, 
    -4.997033, -4.997033, -4.977312, -4.937948, -4.879096, -4.800988, 
    -4.703933, -4.588314, -4.454587, -4.30328, -4.134989, -3.95038, -3.75018, 
    -3.53518, -3.306229, -3.064229, -2.810136, -2.544953, -2.269726, 
    -1.985541, -1.69352, -1.394816, -1.090607, -0.7820941, -0.4704945, 
    -0.1570381,
  // z(51, 0-99)
    0.1569124, 0.4701181, 0.7814684, 1.089735, 1.3937, 1.692165, 1.983952, 
    2.26791, 2.542916, 2.807888, 3.061777, 3.303583, 3.532352, 3.74718, 
    3.947219, 4.131681, 4.299837, 4.451023, 4.584643, 4.70017, 4.797147, 
    4.875192, 4.933997, 4.97333, 4.993035, 4.993035, 4.97333, 4.933997, 
    4.875192, 4.797147, 4.70017, 4.584643, 4.451023, 4.299837, 4.131681, 
    3.947219, 3.74718, 3.532352, 3.303583, 3.061777, 2.807888, 2.542916, 
    2.26791, 1.983952, 1.692165, 1.3937, 1.089735, 0.7814684, 0.4701181, 
    0.1569124, -0.1569124, -0.4701181, -0.7814684, -1.089735, -1.3937, 
    -1.692165, -1.983952, -2.26791, -2.542916, -2.807888, -3.061777, 
    -3.303583, -3.532352, -3.74718, -3.947219, -4.131681, -4.299837, 
    -4.451023, -4.584643, -4.70017, -4.797147, -4.875192, -4.933997, 
    -4.97333, -4.993035, -4.993035, -4.97333, -4.933997, -4.875192, 
    -4.797147, -4.70017, -4.584643, -4.451023, -4.299837, -4.131681, 
    -3.947219, -3.74718, -3.532352, -3.303583, -3.061777, -2.807888, 
    -2.542916, -2.26791, -1.983952, -1.692165, -1.3937, -1.089735, 
    -0.7814684, -0.4701181, -0.1569124,
  // z(52, 0-99)
    0.1566612, 0.4693652, 0.7802169, 1.087989, 1.391468, 1.689455, 1.980775, 
    2.264278, 2.538844, 2.803391, 3.056874, 3.298293, 3.526695, 3.741179, 
    3.940898, 4.125064, 4.292951, 4.443895, 4.577301, 4.692643, 4.789465, 
    4.867385, 4.926095, 4.965365, 4.985039, 4.985039, 4.965365, 4.926095, 
    4.867385, 4.789465, 4.692643, 4.577301, 4.443895, 4.292951, 4.125064, 
    3.940898, 3.741179, 3.526695, 3.298293, 3.056874, 2.803391, 2.538844, 
    2.264278, 1.980775, 1.689455, 1.391468, 1.087989, 0.7802169, 0.4693652, 
    0.1566612, -0.1566612, -0.4693652, -0.7802169, -1.087989, -1.391468, 
    -1.689455, -1.980775, -2.264278, -2.538844, -2.803391, -3.056874, 
    -3.298293, -3.526695, -3.741179, -3.940898, -4.125064, -4.292951, 
    -4.443895, -4.577301, -4.692643, -4.789465, -4.867385, -4.926095, 
    -4.965365, -4.985039, -4.985039, -4.965365, -4.926095, -4.867385, 
    -4.789465, -4.692643, -4.577301, -4.443895, -4.292951, -4.125064, 
    -3.940898, -3.741179, -3.526695, -3.298293, -3.056874, -2.803391, 
    -2.538844, -2.264278, -1.980775, -1.689455, -1.391468, -1.087989, 
    -0.7802169, -0.4693652, -0.1566612,
  // z(53, 0-99)
    0.1562842, 0.4682359, 0.7783397, 1.085372, 1.38812, 1.68539, 1.976009, 
    2.25883, 2.532736, 2.796646, 3.049519, 3.290357, 3.51821, 3.732178, 
    3.931416, 4.115139, 4.282622, 4.433203, 4.566288, 4.681352, 4.777941, 
    4.855674, 4.914243, 4.953419, 4.973045, 4.973045, 4.953419, 4.914243, 
    4.855674, 4.777941, 4.681352, 4.566288, 4.433203, 4.282622, 4.115139, 
    3.931416, 3.732178, 3.51821, 3.290357, 3.049519, 2.796646, 2.532736, 
    2.25883, 1.976009, 1.68539, 1.38812, 1.085372, 0.7783397, 0.4682359, 
    0.1562842, -0.1562842, -0.4682359, -0.7783397, -1.085372, -1.38812, 
    -1.68539, -1.976009, -2.25883, -2.532736, -2.796646, -3.049519, 
    -3.290357, -3.51821, -3.732178, -3.931416, -4.115139, -4.282622, 
    -4.433203, -4.566288, -4.681352, -4.777941, -4.855674, -4.914243, 
    -4.953419, -4.973045, -4.973045, -4.953419, -4.914243, -4.855674, 
    -4.777941, -4.681352, -4.566288, -4.433203, -4.282622, -4.115139, 
    -3.931416, -3.732178, -3.51821, -3.290357, -3.049519, -2.796646, 
    -2.532736, -2.25883, -1.976009, -1.68539, -1.38812, -1.085372, 
    -0.7783397, -0.4682359, -0.1562842,
  // z(54, 0-99)
    0.1557817, 0.4667302, 0.7758367, 1.081881, 1.383656, 1.679971, 1.969655, 
    2.251566, 2.524591, 2.787652, 3.039712, 3.279776, 3.506896, 3.720176, 
    3.918774, 4.101906, 4.26885, 4.418947, 4.551604, 4.666298, 4.762577, 
    4.840059, 4.89844, 4.93749, 4.957053, 4.957053, 4.93749, 4.89844, 
    4.840059, 4.762577, 4.666298, 4.551604, 4.418947, 4.26885, 4.101906, 
    3.918774, 3.720176, 3.506896, 3.279776, 3.039712, 2.787652, 2.524591, 
    2.251566, 1.969655, 1.679971, 1.383656, 1.081881, 0.7758367, 0.4667302, 
    0.1557817, -0.1557817, -0.4667302, -0.7758367, -1.081881, -1.383656, 
    -1.679971, -1.969655, -2.251566, -2.524591, -2.787652, -3.039712, 
    -3.279776, -3.506896, -3.720176, -3.918774, -4.101906, -4.26885, 
    -4.418947, -4.551604, -4.666298, -4.762577, -4.840059, -4.89844, 
    -4.93749, -4.957053, -4.957053, -4.93749, -4.89844, -4.840059, -4.762577, 
    -4.666298, -4.551604, -4.418947, -4.26885, -4.101906, -3.918774, 
    -3.720176, -3.506896, -3.279776, -3.039712, -2.787652, -2.524591, 
    -2.251566, -1.969655, -1.679971, -1.383656, -1.081881, -0.7758367, 
    -0.4667302, -0.1557817,
  // z(55, 0-99)
    0.1551534, 0.464848, 0.7727081, 1.077519, 1.378077, 1.673196, 1.961712, 
    2.242486, 2.51441, 2.776411, 3.027454, 3.26655, 3.492754, 3.705174, 
    3.902971, 4.085364, 4.251635, 4.401127, 4.533249, 4.64748, 4.743371, 
    4.820541, 4.878686, 4.917578, 4.937063, 4.937063, 4.917578, 4.878686, 
    4.820541, 4.743371, 4.64748, 4.533249, 4.401127, 4.251635, 4.085364, 
    3.902971, 3.705174, 3.492754, 3.26655, 3.027454, 2.776411, 2.51441, 
    2.242486, 1.961712, 1.673196, 1.378077, 1.077519, 0.7727081, 0.464848, 
    0.1551534, -0.1551534, -0.464848, -0.7727081, -1.077519, -1.378077, 
    -1.673196, -1.961712, -2.242486, -2.51441, -2.776411, -3.027454, 
    -3.26655, -3.492754, -3.705174, -3.902971, -4.085364, -4.251635, 
    -4.401127, -4.533249, -4.64748, -4.743371, -4.820541, -4.878686, 
    -4.917578, -4.937063, -4.937063, -4.917578, -4.878686, -4.820541, 
    -4.743371, -4.64748, -4.533249, -4.401127, -4.251635, -4.085364, 
    -3.902971, -3.705174, -3.492754, -3.26655, -3.027454, -2.776411, 
    -2.51441, -2.242486, -1.961712, -1.673196, -1.378077, -1.077519, 
    -0.7727081, -0.464848, -0.1551534,
  // z(56, 0-99)
    0.1543996, 0.4625894, 0.7689536, 1.072283, 1.371381, 1.665066, 1.952181, 
    2.23159, 2.502193, 2.762921, 3.012745, 3.250679, 3.475783, 3.687171, 
    3.884007, 4.065515, 4.230978, 4.379743, 4.511223, 4.624899, 4.720324, 
    4.797119, 4.854982, 4.893685, 4.913074, 4.913074, 4.893685, 4.854982, 
    4.797119, 4.720324, 4.624899, 4.511223, 4.379743, 4.230978, 4.065515, 
    3.884007, 3.687171, 3.475783, 3.250679, 3.012745, 2.762921, 2.502193, 
    2.23159, 1.952181, 1.665066, 1.371381, 1.072283, 0.7689536, 0.4625894, 
    0.1543996, -0.1543996, -0.4625894, -0.7689536, -1.072283, -1.371381, 
    -1.665066, -1.952181, -2.23159, -2.502193, -2.762921, -3.012745, 
    -3.250679, -3.475783, -3.687171, -3.884007, -4.065515, -4.230978, 
    -4.379743, -4.511223, -4.624899, -4.720324, -4.797119, -4.854982, 
    -4.893685, -4.913074, -4.913074, -4.893685, -4.854982, -4.797119, 
    -4.720324, -4.624899, -4.511223, -4.379743, -4.230978, -4.065515, 
    -3.884007, -3.687171, -3.475783, -3.250679, -3.012745, -2.762921, 
    -2.502193, -2.23159, -1.952181, -1.665066, -1.371381, -1.072283, 
    -0.7689536, -0.4625894, -0.1543996,
  // z(57, 0-99)
    0.1535201, 0.4599544, 0.7645735, 1.066175, 1.363569, 1.655582, 1.94106, 
    2.218879, 2.48794, 2.747183, 2.995583, 3.232162, 3.455984, 3.666168, 
    3.861883, 4.042356, 4.206877, 4.354795, 4.485526, 4.598555, 4.693435, 
    4.769793, 4.827327, 4.865809, 4.885088, 4.885088, 4.865809, 4.827327, 
    4.769793, 4.693435, 4.598555, 4.485526, 4.354795, 4.206877, 4.042356, 
    3.861883, 3.666168, 3.455984, 3.232162, 2.995583, 2.747183, 2.48794, 
    2.218879, 1.94106, 1.655582, 1.363569, 1.066175, 0.7645735, 0.4599544, 
    0.1535201, -0.1535201, -0.4599544, -0.7645735, -1.066175, -1.363569, 
    -1.655582, -1.94106, -2.218879, -2.48794, -2.747183, -2.995583, 
    -3.232162, -3.455984, -3.666168, -3.861883, -4.042356, -4.206877, 
    -4.354795, -4.485526, -4.598555, -4.693435, -4.769793, -4.827327, 
    -4.865809, -4.885088, -4.885088, -4.865809, -4.827327, -4.769793, 
    -4.693435, -4.598555, -4.485526, -4.354795, -4.206877, -4.042356, 
    -3.861883, -3.666168, -3.455984, -3.232162, -2.995583, -2.747183, 
    -2.48794, -2.218879, -1.94106, -1.655582, -1.363569, -1.066175, 
    -0.7645735, -0.4599544, -0.1535201,
  // z(58, 0-99)
    0.1525149, 0.4569429, 0.7595676, 1.059195, 1.354641, 1.644742, 1.928352, 
    2.204351, 2.471651, 2.729196, 2.97597, 3.211, 3.433357, 3.642164, 
    3.836598, 4.01589, 4.179333, 4.326282, 4.456158, 4.568447, 4.662706, 
    4.738564, 4.795721, 4.833951, 4.853104, 4.853104, 4.833951, 4.795721, 
    4.738564, 4.662706, 4.568447, 4.456158, 4.326282, 4.179333, 4.01589, 
    3.836598, 3.642164, 3.433357, 3.211, 2.97597, 2.729196, 2.471651, 
    2.204351, 1.928352, 1.644742, 1.354641, 1.059195, 0.7595676, 0.4569429, 
    0.1525149, -0.1525149, -0.4569429, -0.7595676, -1.059195, -1.354641, 
    -1.644742, -1.928352, -2.204351, -2.471651, -2.729196, -2.97597, -3.211, 
    -3.433357, -3.642164, -3.836598, -4.01589, -4.179333, -4.326282, 
    -4.456158, -4.568447, -4.662706, -4.738564, -4.795721, -4.833951, 
    -4.853104, -4.853104, -4.833951, -4.795721, -4.738564, -4.662706, 
    -4.568447, -4.456158, -4.326282, -4.179333, -4.01589, -3.836598, 
    -3.642164, -3.433357, -3.211, -2.97597, -2.729196, -2.471651, -2.204351, 
    -1.928352, -1.644742, -1.354641, -1.059195, -0.7595676, -0.4569429, 
    -0.1525149,
  // z(59, 0-99)
    0.1513842, 0.453555, 0.7539359, 1.051341, 1.344598, 1.632547, 1.914054, 
    2.188007, 2.453325, 2.708961, 2.953906, 3.187192, 3.407901, 3.61516, 
    3.808152, 3.986115, 4.148346, 4.294206, 4.423119, 4.534575, 4.628135, 
    4.703431, 4.760164, 4.798111, 4.817122, 4.817122, 4.798111, 4.760164, 
    4.703431, 4.628135, 4.534575, 4.423119, 4.294206, 4.148346, 3.986115, 
    3.808152, 3.61516, 3.407901, 3.187192, 2.953906, 2.708961, 2.453325, 
    2.188007, 1.914054, 1.632547, 1.344598, 1.051341, 0.7539359, 0.453555, 
    0.1513842, -0.1513842, -0.453555, -0.7539359, -1.051341, -1.344598, 
    -1.632547, -1.914054, -2.188007, -2.453325, -2.708961, -2.953906, 
    -3.187192, -3.407901, -3.61516, -3.808152, -3.986115, -4.148346, 
    -4.294206, -4.423119, -4.534575, -4.628135, -4.703431, -4.760164, 
    -4.798111, -4.817122, -4.817122, -4.798111, -4.760164, -4.703431, 
    -4.628135, -4.534575, -4.423119, -4.294206, -4.148346, -3.986115, 
    -3.808152, -3.61516, -3.407901, -3.187192, -2.953906, -2.708961, 
    -2.453325, -2.188007, -1.914054, -1.632547, -1.344598, -1.051341, 
    -0.7539359, -0.453555, -0.1513842,
  // z(60, 0-99)
    0.1501277, 0.4497907, 0.7476785, 1.042616, 1.333438, 1.618998, 1.898168, 
    2.169847, 2.432963, 2.686477, 2.929389, 3.16074, 3.379617, 3.585156, 
    3.776546, 3.953032, 4.113916, 4.258566, 4.386408, 4.49694, 4.589724, 
    4.664394, 4.720656, 4.758288, 4.777142, 4.777142, 4.758288, 4.720656, 
    4.664394, 4.589724, 4.49694, 4.386408, 4.258566, 4.113916, 3.953032, 
    3.776546, 3.585156, 3.379617, 3.16074, 2.929389, 2.686477, 2.432963, 
    2.169847, 1.898168, 1.618998, 1.333438, 1.042616, 0.7476785, 0.4497907, 
    0.1501277, -0.1501277, -0.4497907, -0.7476785, -1.042616, -1.333438, 
    -1.618998, -1.898168, -2.169847, -2.432963, -2.686477, -2.929389, 
    -3.16074, -3.379617, -3.585156, -3.776546, -3.953032, -4.113916, 
    -4.258566, -4.386408, -4.49694, -4.589724, -4.664394, -4.720656, 
    -4.758288, -4.777142, -4.777142, -4.758288, -4.720656, -4.664394, 
    -4.589724, -4.49694, -4.386408, -4.258566, -4.113916, -3.953032, 
    -3.776546, -3.585156, -3.379617, -3.16074, -2.929389, -2.686477, 
    -2.432963, -2.169847, -1.898168, -1.618998, -1.333438, -1.042616, 
    -0.7476785, -0.4497907, -0.1501277,
  // z(61, 0-99)
    0.1487457, 0.4456499, 0.7407954, 1.033017, 1.321162, 1.604093, 1.880694, 
    2.149872, 2.410566, 2.661746, 2.902421, 3.131642, 3.348504, 3.552151, 
    3.741779, 3.91664, 4.076044, 4.219361, 4.346027, 4.455541, 4.547471, 
    4.621454, 4.677198, 4.714484, 4.733163, 4.733163, 4.714484, 4.677198, 
    4.621454, 4.547471, 4.455541, 4.346027, 4.219361, 4.076044, 3.91664, 
    3.741779, 3.552151, 3.348504, 3.131642, 2.902421, 2.661746, 2.410566, 
    2.149872, 1.880694, 1.604093, 1.321162, 1.033017, 0.7407954, 0.4456499, 
    0.1487457, -0.1487457, -0.4456499, -0.7407954, -1.033017, -1.321162, 
    -1.604093, -1.880694, -2.149872, -2.410566, -2.661746, -2.902421, 
    -3.131642, -3.348504, -3.552151, -3.741779, -3.91664, -4.076044, 
    -4.219361, -4.346027, -4.455541, -4.547471, -4.621454, -4.677198, 
    -4.714484, -4.733163, -4.733163, -4.714484, -4.677198, -4.621454, 
    -4.547471, -4.455541, -4.346027, -4.219361, -4.076044, -3.91664, 
    -3.741779, -3.552151, -3.348504, -3.131642, -2.902421, -2.661746, 
    -2.410566, -2.149872, -1.880694, -1.604093, -1.321162, -1.033017, 
    -0.7407954, -0.4456499, -0.1487457,
  // z(62, 0-99)
    0.1472379, 0.4411327, 0.7332866, 1.022546, 1.307771, 1.587834, 1.861631, 
    2.12808, 2.386132, 2.634766, 2.873002, 3.099899, 3.314563, 3.516146, 
    3.703852, 3.87694, 4.034728, 4.176593, 4.301975, 4.410378, 4.501377, 
    4.57461, 4.629789, 4.666697, 4.685187, 4.685187, 4.666697, 4.629789, 
    4.57461, 4.501377, 4.410378, 4.301975, 4.176593, 4.034728, 3.87694, 
    3.703852, 3.516146, 3.314563, 3.099899, 2.873002, 2.634766, 2.386132, 
    2.12808, 1.861631, 1.587834, 1.307771, 1.022546, 0.7332866, 0.4411327, 
    0.1472379, -0.1472379, -0.4411327, -0.7332866, -1.022546, -1.307771, 
    -1.587834, -1.861631, -2.12808, -2.386132, -2.634766, -2.873002, 
    -3.099899, -3.314563, -3.516146, -3.703852, -3.87694, -4.034728, 
    -4.176593, -4.301975, -4.410378, -4.501377, -4.57461, -4.629789, 
    -4.666697, -4.685187, -4.685187, -4.666697, -4.629789, -4.57461, 
    -4.501377, -4.410378, -4.301975, -4.176593, -4.034728, -3.87694, 
    -3.703852, -3.516146, -3.314563, -3.099899, -2.873002, -2.634766, 
    -2.386132, -2.12808, -1.861631, -1.587834, -1.307771, -1.022546, 
    -0.7332866, -0.4411327, -0.1472379,
  // z(63, 0-99)
    0.1456046, 0.4362391, 0.725152, 1.011203, 1.293263, 1.57022, 1.840979, 
    2.104473, 2.359662, 2.605537, 2.841131, 3.065511, 3.277793, 3.47714, 
    3.662764, 3.833932, 3.98997, 4.130261, 4.254251, 4.361453, 4.451441, 
    4.523862, 4.578429, 4.614927, 4.633213, 4.633213, 4.614927, 4.578429, 
    4.523862, 4.451441, 4.361453, 4.254251, 4.130261, 3.98997, 3.833932, 
    3.662764, 3.47714, 3.277793, 3.065511, 2.841131, 2.605537, 2.359662, 
    2.104473, 1.840979, 1.57022, 1.293263, 1.011203, 0.725152, 0.4362391, 
    0.1456046, -0.1456046, -0.4362391, -0.725152, -1.011203, -1.293263, 
    -1.57022, -1.840979, -2.104473, -2.359662, -2.605537, -2.841131, 
    -3.065511, -3.277793, -3.47714, -3.662764, -3.833932, -3.98997, 
    -4.130261, -4.254251, -4.361453, -4.451441, -4.523862, -4.578429, 
    -4.614927, -4.633213, -4.633213, -4.614927, -4.578429, -4.523862, 
    -4.451441, -4.361453, -4.254251, -4.130261, -3.98997, -3.833932, 
    -3.662764, -3.47714, -3.277793, -3.065511, -2.841131, -2.605537, 
    -2.359662, -2.104473, -1.840979, -1.57022, -1.293263, -1.011203, 
    -0.725152, -0.4362391, -0.1456046,
  // z(64, 0-99)
    0.1438456, 0.430969, 0.7163916, 0.998987, 1.27764, 1.55125, 1.818739, 
    2.07905, 2.331155, 2.574061, 2.806808, 3.028478, 3.238195, 3.435134, 
    3.618515, 3.787616, 3.941768, 4.080364, 4.202857, 4.308764, 4.397665, 
    4.469211, 4.523119, 4.559176, 4.57724, 4.57724, 4.559176, 4.523119, 
    4.469211, 4.397665, 4.308764, 4.202857, 4.080364, 3.941768, 3.787616, 
    3.618515, 3.435134, 3.238195, 3.028478, 2.806808, 2.574061, 2.331155, 
    2.07905, 1.818739, 1.55125, 1.27764, 0.998987, 0.7163916, 0.430969, 
    0.1438456, -0.1438456, -0.430969, -0.7163916, -0.998987, -1.27764, 
    -1.55125, -1.818739, -2.07905, -2.331155, -2.574061, -2.806808, 
    -3.028478, -3.238195, -3.435134, -3.618515, -3.787616, -3.941768, 
    -4.080364, -4.202857, -4.308764, -4.397665, -4.469211, -4.523119, 
    -4.559176, -4.57724, -4.57724, -4.559176, -4.523119, -4.469211, 
    -4.397665, -4.308764, -4.202857, -4.080364, -3.941768, -3.787616, 
    -3.618515, -3.435134, -3.238195, -3.028478, -2.806808, -2.574061, 
    -2.331155, -2.07905, -1.818739, -1.55125, -1.27764, -0.998987, 
    -0.7163916, -0.430969, -0.1438456,
  // z(65, 0-99)
    0.1419609, 0.4253225, 0.7070056, 0.9858984, 1.2609, 1.530926, 1.79491, 
    2.05181, 2.300613, 2.540336, 2.770033, 2.988799, 3.195769, 3.390127, 
    3.571105, 3.737991, 3.890124, 4.026904, 4.147792, 4.252311, 4.340047, 
    4.410656, 4.463858, 4.499442, 4.51727, 4.51727, 4.499442, 4.463858, 
    4.410656, 4.340047, 4.252311, 4.147792, 4.026904, 3.890124, 3.737991, 
    3.571105, 3.390127, 3.195769, 2.988799, 2.770033, 2.540336, 2.300613, 
    2.05181, 1.79491, 1.530926, 1.2609, 0.9858984, 0.7070056, 0.4253225, 
    0.1419609, -0.1419609, -0.4253225, -0.7070056, -0.9858984, -1.2609, 
    -1.530926, -1.79491, -2.05181, -2.300613, -2.540336, -2.770033, 
    -2.988799, -3.195769, -3.390127, -3.571105, -3.737991, -3.890124, 
    -4.026904, -4.147792, -4.252311, -4.340047, -4.410656, -4.463858, 
    -4.499442, -4.51727, -4.51727, -4.499442, -4.463858, -4.410656, 
    -4.340047, -4.252311, -4.147792, -4.026904, -3.890124, -3.737991, 
    -3.571105, -3.390127, -3.195769, -2.988799, -2.770033, -2.540336, 
    -2.300613, -2.05181, -1.79491, -1.530926, -1.2609, -0.9858984, 
    -0.7070056, -0.4253225, -0.1419609,
  // z(66, 0-99)
    0.1399506, 0.4192996, 0.6969938, 0.9719372, 1.243045, 1.509247, 1.769492, 
    2.022755, 2.268034, 2.504363, 2.730807, 2.946475, 3.150514, 3.34212, 
    3.520536, 3.685057, 3.835036, 3.96988, 4.089056, 4.192094, 4.278588, 
    4.348197, 4.400645, 4.435726, 4.453301, 4.453301, 4.435726, 4.400645, 
    4.348197, 4.278588, 4.192094, 4.089056, 3.96988, 3.835036, 3.685057, 
    3.520536, 3.34212, 3.150514, 2.946475, 2.730807, 2.504363, 2.268034, 
    2.022755, 1.769492, 1.509247, 1.243045, 0.9719372, 0.6969938, 0.4192996, 
    0.1399506, -0.1399506, -0.4192996, -0.6969938, -0.9719372, -1.243045, 
    -1.509247, -1.769492, -2.022755, -2.268034, -2.504363, -2.730807, 
    -2.946475, -3.150514, -3.34212, -3.520536, -3.685057, -3.835036, 
    -3.96988, -4.089056, -4.192094, -4.278588, -4.348197, -4.400645, 
    -4.435726, -4.453301, -4.453301, -4.435726, -4.400645, -4.348197, 
    -4.278588, -4.192094, -4.089056, -3.96988, -3.835036, -3.685057, 
    -3.520536, -3.34212, -3.150514, -2.946475, -2.730807, -2.504363, 
    -2.268034, -2.022755, -1.769492, -1.509247, -1.243045, -0.9719372, 
    -0.6969938, -0.4192996, -0.1399506,
  // z(67, 0-99)
    0.1378147, 0.4129002, 0.6863562, 0.9571035, 1.224074, 1.486213, 1.742486, 
    1.991883, 2.233419, 2.466141, 2.68913, 2.901506, 3.102431, 3.291112, 
    3.466805, 3.628816, 3.776506, 3.909291, 4.026649, 4.128114, 4.213289, 
    4.281835, 4.333483, 4.368028, 4.385335, 4.385335, 4.368028, 4.333483, 
    4.281835, 4.213289, 4.128114, 4.026649, 3.909291, 3.776506, 3.628816, 
    3.466805, 3.291112, 3.102431, 2.901506, 2.68913, 2.466141, 2.233419, 
    1.991883, 1.742486, 1.486213, 1.224074, 0.9571035, 0.6863562, 0.4129002, 
    0.1378147, -0.1378147, -0.4129002, -0.6863562, -0.9571035, -1.224074, 
    -1.486213, -1.742486, -1.991883, -2.233419, -2.466141, -2.68913, 
    -2.901506, -3.102431, -3.291112, -3.466805, -3.628816, -3.776506, 
    -3.909291, -4.026649, -4.128114, -4.213289, -4.281835, -4.333483, 
    -4.368028, -4.385335, -4.385335, -4.368028, -4.333483, -4.281835, 
    -4.213289, -4.128114, -4.026649, -3.909291, -3.776506, -3.628816, 
    -3.466805, -3.291112, -3.102431, -2.901506, -2.68913, -2.466141, 
    -2.233419, -1.991883, -1.742486, -1.486213, -1.224074, -0.9571035, 
    -0.6863562, -0.4129002, -0.1378147,
  // z(68, 0-99)
    0.1355531, 0.4061244, 0.6750929, 0.9413971, 1.203986, 1.461823, 1.713892, 
    1.959196, 2.196768, 2.425671, 2.645, 2.853891, 3.051519, 3.237104, 
    3.409914, 3.569266, 3.714532, 3.845139, 3.96057, 4.060371, 4.144147, 
    4.211569, 4.262369, 4.296348, 4.313371, 4.313371, 4.296348, 4.262369, 
    4.211569, 4.144147, 4.060371, 3.96057, 3.845139, 3.714532, 3.569266, 
    3.409914, 3.237104, 3.051519, 2.853891, 2.645, 2.425671, 2.196768, 
    1.959196, 1.713892, 1.461823, 1.203986, 0.9413971, 0.6750929, 0.4061244, 
    0.1355531, -0.1355531, -0.4061244, -0.6750929, -0.9413971, -1.203986, 
    -1.461823, -1.713892, -1.959196, -2.196768, -2.425671, -2.645, -2.853891, 
    -3.051519, -3.237104, -3.409914, -3.569266, -3.714532, -3.845139, 
    -3.96057, -4.060371, -4.144147, -4.211569, -4.262369, -4.296348, 
    -4.313371, -4.313371, -4.296348, -4.262369, -4.211569, -4.144147, 
    -4.060371, -3.96057, -3.845139, -3.714532, -3.569266, -3.409914, 
    -3.237104, -3.051519, -2.853891, -2.645, -2.425671, -2.196768, -1.959196, 
    -1.713892, -1.461823, -1.203986, -0.9413971, -0.6750929, -0.4061244, 
    -0.1355531,
  // z(69, 0-99)
    0.1331659, 0.3989722, 0.6632039, 0.9248183, 1.182783, 1.436079, 1.683708, 
    1.924693, 2.158081, 2.382952, 2.598419, 2.803632, 2.997779, 3.180096, 
    3.349862, 3.506408, 3.649116, 3.777422, 3.890821, 3.988864, 4.071165, 
    4.137399, 4.187304, 4.220685, 4.237408, 4.237408, 4.220685, 4.187304, 
    4.137399, 4.071165, 3.988864, 3.890821, 3.777422, 3.649116, 3.506408, 
    3.349862, 3.180096, 2.997779, 2.803632, 2.598419, 2.382952, 2.158081, 
    1.924693, 1.683708, 1.436079, 1.182783, 0.9248183, 0.6632039, 0.3989722, 
    0.1331659, -0.1331659, -0.3989722, -0.6632039, -0.9248183, -1.182783, 
    -1.436079, -1.683708, -1.924693, -2.158081, -2.382952, -2.598419, 
    -2.803632, -2.997779, -3.180096, -3.349862, -3.506408, -3.649116, 
    -3.777422, -3.890821, -3.988864, -4.071165, -4.137399, -4.187304, 
    -4.220685, -4.237408, -4.237408, -4.220685, -4.187304, -4.137399, 
    -4.071165, -3.988864, -3.890821, -3.777422, -3.649116, -3.506408, 
    -3.349862, -3.180096, -2.997779, -2.803632, -2.598419, -2.382952, 
    -2.158081, -1.924693, -1.683708, -1.436079, -1.182783, -0.9248183, 
    -0.6632039, -0.3989722, -0.1331659,
  // z(70, 0-99)
    0.1306531, 0.3914435, 0.6506892, 0.9073668, 1.160463, 1.40898, 1.651937, 
    1.888373, 2.117358, 2.337986, 2.549387, 2.750727, 2.941211, 3.120087, 
    3.28665, 3.440242, 3.580256, 3.706142, 3.8174, 3.913594, 3.994342, 
    4.059326, 4.10829, 4.14104, 4.157447, 4.157447, 4.14104, 4.10829, 
    4.059326, 3.994342, 3.913594, 3.8174, 3.706142, 3.580256, 3.440242, 
    3.28665, 3.120087, 2.941211, 2.750727, 2.549387, 2.337986, 2.117358, 
    1.888373, 1.651937, 1.40898, 1.160463, 0.9073668, 0.6506892, 0.3914435, 
    0.1306531, -0.1306531, -0.3914435, -0.6506892, -0.9073668, -1.160463, 
    -1.40898, -1.651937, -1.888373, -2.117358, -2.337986, -2.549387, 
    -2.750727, -2.941211, -3.120087, -3.28665, -3.440242, -3.580256, 
    -3.706142, -3.8174, -3.913594, -3.994342, -4.059326, -4.10829, -4.14104, 
    -4.157447, -4.157447, -4.14104, -4.10829, -4.059326, -3.994342, 
    -3.913594, -3.8174, -3.706142, -3.580256, -3.440242, -3.28665, -3.120087, 
    -2.941211, -2.750727, -2.549387, -2.337986, -2.117358, -1.888373, 
    -1.651937, -1.40898, -1.160463, -0.9073668, -0.6506892, -0.3914435, 
    -0.1306531,
  // z(71, 0-99)
    0.1280145, 0.3835384, 0.6375487, 0.8890428, 1.137028, 1.380526, 1.618576, 
    1.850238, 2.074598, 2.290771, 2.497903, 2.695177, 2.881814, 3.057078, 
    3.220277, 3.370767, 3.507954, 3.631297, 3.740309, 3.83456, 3.913677, 
    3.977349, 4.025324, 4.057413, 4.073489, 4.073489, 4.057413, 4.025324, 
    3.977349, 3.913677, 3.83456, 3.740309, 3.631297, 3.507954, 3.370767, 
    3.220277, 3.057078, 2.881814, 2.695177, 2.497903, 2.290771, 2.074598, 
    1.850238, 1.618576, 1.380526, 1.137028, 0.8890428, 0.6375487, 0.3835384, 
    0.1280145, -0.1280145, -0.3835384, -0.6375487, -0.8890428, -1.137028, 
    -1.380526, -1.618576, -1.850238, -2.074598, -2.290771, -2.497903, 
    -2.695177, -2.881814, -3.057078, -3.220277, -3.370767, -3.507954, 
    -3.631297, -3.740309, -3.83456, -3.913677, -3.977349, -4.025324, 
    -4.057413, -4.073489, -4.073489, -4.057413, -4.025324, -3.977349, 
    -3.913677, -3.83456, -3.740309, -3.631297, -3.507954, -3.370767, 
    -3.220277, -3.057078, -2.881814, -2.695177, -2.497903, -2.290771, 
    -2.074598, -1.850238, -1.618576, -1.380526, -1.137028, -0.8890428, 
    -0.6375487, -0.3835384, -0.1280145,
  // z(72, 0-99)
    0.1252504, 0.3752569, 0.6237825, 0.8698462, 1.112477, 1.350717, 1.583627, 
    1.810287, 2.029803, 2.241307, 2.443967, 2.636981, 2.819588, 2.991068, 
    3.150743, 3.297984, 3.432209, 3.552889, 3.659547, 3.751762, 3.829171, 
    3.891468, 3.938407, 3.969803, 3.985533, 3.985533, 3.969803, 3.938407, 
    3.891468, 3.829171, 3.751762, 3.659547, 3.552889, 3.432209, 3.297984, 
    3.150743, 2.991068, 2.819588, 2.636981, 2.443967, 2.241307, 2.029803, 
    1.810287, 1.583627, 1.350717, 1.112477, 0.8698462, 0.6237825, 0.3752569, 
    0.1252504, -0.1252504, -0.3752569, -0.6237825, -0.8698462, -1.112477, 
    -1.350717, -1.583627, -1.810287, -2.029803, -2.241307, -2.443967, 
    -2.636981, -2.819588, -2.991068, -3.150743, -3.297984, -3.432209, 
    -3.552889, -3.659547, -3.751762, -3.829171, -3.891468, -3.938407, 
    -3.969803, -3.985533, -3.985533, -3.969803, -3.938407, -3.891468, 
    -3.829171, -3.751762, -3.659547, -3.552889, -3.432209, -3.297984, 
    -3.150743, -2.991068, -2.819588, -2.636981, -2.443967, -2.241307, 
    -2.029803, -1.810287, -1.583627, -1.350717, -1.112477, -0.8698462, 
    -0.6237825, -0.3752569, -0.1252504,
  // z(73, 0-99)
    0.1223606, 0.3665989, 0.6093904, 0.849777, 1.08681, 1.319554, 1.54709, 
    1.76852, 1.982971, 2.189596, 2.387579, 2.57614, 2.754534, 2.922058, 
    3.078049, 3.221892, 3.353021, 3.470916, 3.575113, 3.665201, 3.740824, 
    3.801684, 3.84754, 3.878212, 3.893578, 3.893578, 3.878212, 3.84754, 
    3.801684, 3.740824, 3.665201, 3.575113, 3.470916, 3.353021, 3.221892, 
    3.078049, 2.922058, 2.754534, 2.57614, 2.387579, 2.189596, 1.982971, 
    1.76852, 1.54709, 1.319554, 1.08681, 0.849777, 0.6093904, 0.3665989, 
    0.1223606, -0.1223606, -0.3665989, -0.6093904, -0.849777, -1.08681, 
    -1.319554, -1.54709, -1.76852, -1.982971, -2.189596, -2.387579, -2.57614, 
    -2.754534, -2.922058, -3.078049, -3.221892, -3.353021, -3.470916, 
    -3.575113, -3.665201, -3.740824, -3.801684, -3.84754, -3.878212, 
    -3.893578, -3.893578, -3.878212, -3.84754, -3.801684, -3.740824, 
    -3.665201, -3.575113, -3.470916, -3.353021, -3.221892, -3.078049, 
    -2.922058, -2.754534, -2.57614, -2.387579, -2.189596, -1.982971, 
    -1.76852, -1.54709, -1.319554, -1.08681, -0.849777, -0.6093904, 
    -0.3665989, -0.1223606,
  // z(74, 0-99)
    0.1193452, 0.3575645, 0.5943727, 0.8288352, 1.060027, 1.287035, 1.508963, 
    1.724937, 1.934103, 2.135636, 2.32874, 2.512655, 2.686652, 2.850047, 
    3.002194, 3.142493, 3.270389, 3.385379, 3.487009, 3.574877, 3.648636, 
    3.707996, 3.752722, 3.782638, 3.797625, 3.797625, 3.782638, 3.752722, 
    3.707996, 3.648636, 3.574877, 3.487009, 3.385379, 3.270389, 3.142493, 
    3.002194, 2.850047, 2.686652, 2.512655, 2.32874, 2.135636, 1.934103, 
    1.724937, 1.508963, 1.287035, 1.060027, 0.8288352, 0.5943727, 0.3575645, 
    0.1193452, -0.1193452, -0.3575645, -0.5943727, -0.8288352, -1.060027, 
    -1.287035, -1.508963, -1.724937, -1.934103, -2.135636, -2.32874, 
    -2.512655, -2.686652, -2.850047, -3.002194, -3.142493, -3.270389, 
    -3.385379, -3.487009, -3.574877, -3.648636, -3.707996, -3.752722, 
    -3.782638, -3.797625, -3.797625, -3.782638, -3.752722, -3.707996, 
    -3.648636, -3.574877, -3.487009, -3.385379, -3.270389, -3.142493, 
    -3.002194, -2.850047, -2.686652, -2.512655, -2.32874, -2.135636, 
    -1.934103, -1.724937, -1.508963, -1.287035, -1.060027, -0.8288352, 
    -0.5943727, -0.3575645, -0.1193452,
  // z(75, 0-99)
    0.1162041, 0.3481537, 0.5787293, 0.8070209, 1.032128, 1.253161, 1.469249, 
    1.679538, 1.883199, 2.079427, 2.26745, 2.446523, 2.615942, 2.775036, 
    2.923178, 3.059785, 3.184315, 3.296279, 3.395233, 3.480788, 3.552607, 
    3.610404, 3.653953, 3.683081, 3.697675, 3.697675, 3.683081, 3.653953, 
    3.610404, 3.552607, 3.480788, 3.395233, 3.296279, 3.184315, 3.059785, 
    2.923178, 2.775036, 2.615942, 2.446523, 2.26745, 2.079427, 1.883199, 
    1.679538, 1.469249, 1.253161, 1.032128, 0.8070209, 0.5787293, 0.3481537, 
    0.1162041, -0.1162041, -0.3481537, -0.5787293, -0.8070209, -1.032128, 
    -1.253161, -1.469249, -1.679538, -1.883199, -2.079427, -2.26745, 
    -2.446523, -2.615942, -2.775036, -2.923178, -3.059785, -3.184315, 
    -3.296279, -3.395233, -3.480788, -3.552607, -3.610404, -3.653953, 
    -3.683081, -3.697675, -3.697675, -3.683081, -3.653953, -3.610404, 
    -3.552607, -3.480788, -3.395233, -3.296279, -3.184315, -3.059785, 
    -2.923178, -2.775036, -2.615942, -2.446523, -2.26745, -2.079427, 
    -1.883199, -1.679538, -1.469249, -1.253161, -1.032128, -0.8070209, 
    -0.5787293, -0.3481537, -0.1162041,
  // z(76, 0-99)
    0.1129374, 0.3383664, 0.5624601, 0.784334, 1.003113, 1.217932, 1.427945, 
    1.632323, 1.830258, 2.020971, 2.203707, 2.377747, 2.542403, 2.697024, 
    2.841002, 2.973768, 3.094798, 3.203614, 3.299787, 3.382937, 3.452736, 
    3.508909, 3.551234, 3.579543, 3.593726, 3.593726, 3.579543, 3.551234, 
    3.508909, 3.452736, 3.382937, 3.299787, 3.203614, 3.094798, 2.973768, 
    2.841002, 2.697024, 2.542403, 2.377747, 2.203707, 2.020971, 1.830258, 
    1.632323, 1.427945, 1.217932, 1.003113, 0.784334, 0.5624601, 0.3383664, 
    0.1129374, -0.1129374, -0.3383664, -0.5624601, -0.784334, -1.003113, 
    -1.217932, -1.427945, -1.632323, -1.830258, -2.020971, -2.203707, 
    -2.377747, -2.542403, -2.697024, -2.841002, -2.973768, -3.094798, 
    -3.203614, -3.299787, -3.382937, -3.452736, -3.508909, -3.551234, 
    -3.579543, -3.593726, -3.593726, -3.579543, -3.551234, -3.508909, 
    -3.452736, -3.382937, -3.299787, -3.203614, -3.094798, -2.973768, 
    -2.841002, -2.697024, -2.542403, -2.377747, -2.203707, -2.020971, 
    -1.830258, -1.632323, -1.427945, -1.217932, -1.003113, -0.784334, 
    -0.5624601, -0.3383664, -0.1129374,
  // z(77, 0-99)
    0.109545, 0.3282028, 0.5455652, 0.7607746, 0.9729815, 1.181348, 1.385053, 
    1.583292, 1.775282, 1.960266, 2.137513, 2.306325, 2.466035, 2.616012, 
    2.755666, 2.884444, 3.001838, 3.107385, 3.200669, 3.281322, 3.349024, 
    3.40351, 3.444563, 3.472022, 3.485779, 3.485779, 3.472022, 3.444563, 
    3.40351, 3.349024, 3.281322, 3.200669, 3.107385, 3.001838, 2.884444, 
    2.755666, 2.616012, 2.466035, 2.306325, 2.137513, 1.960266, 1.775282, 
    1.583292, 1.385053, 1.181348, 0.9729815, 0.7607746, 0.5455652, 0.3282028, 
    0.109545, -0.109545, -0.3282028, -0.5455652, -0.7607746, -0.9729815, 
    -1.181348, -1.385053, -1.583292, -1.775282, -1.960266, -2.137513, 
    -2.306325, -2.466035, -2.616012, -2.755666, -2.884444, -3.001838, 
    -3.107385, -3.200669, -3.281322, -3.349024, -3.40351, -3.444563, 
    -3.472022, -3.485779, -3.485779, -3.472022, -3.444563, -3.40351, 
    -3.349024, -3.281322, -3.200669, -3.107385, -3.001838, -2.884444, 
    -2.755666, -2.616012, -2.466035, -2.306325, -2.137513, -1.960266, 
    -1.775282, -1.583292, -1.385053, -1.181348, -0.9729815, -0.7607746, 
    -0.5455652, -0.3282028, -0.109545,
  // z(78, 0-99)
    0.106027, 0.3176626, 0.5280445, 0.7363425, 0.9417345, 1.14341, 1.340573, 
    1.532445, 1.718269, 1.897312, 2.068868, 2.232258, 2.386839, 2.532, 
    2.667168, 2.791811, 2.905435, 3.007592, 3.097881, 3.175943, 3.241471, 
    3.294207, 3.333942, 3.360519, 3.373834, 3.373834, 3.360519, 3.333942, 
    3.294207, 3.241471, 3.175943, 3.097881, 3.007592, 2.905435, 2.791811, 
    2.667168, 2.532, 2.386839, 2.232258, 2.068868, 1.897312, 1.718269, 
    1.532445, 1.340573, 1.14341, 0.9417345, 0.7363425, 0.5280445, 0.3176626, 
    0.106027, -0.106027, -0.3176626, -0.5280445, -0.7363425, -0.9417345, 
    -1.14341, -1.340573, -1.532445, -1.718269, -1.897312, -2.068868, 
    -2.232258, -2.386839, -2.532, -2.667168, -2.791811, -2.905435, -3.007592, 
    -3.097881, -3.175943, -3.241471, -3.294207, -3.333942, -3.360519, 
    -3.373834, -3.373834, -3.360519, -3.333942, -3.294207, -3.241471, 
    -3.175943, -3.097881, -3.007592, -2.905435, -2.791811, -2.667168, -2.532, 
    -2.386839, -2.232258, -2.068868, -1.897312, -1.718269, -1.532445, 
    -1.340573, -1.14341, -0.9417345, -0.7363425, -0.5280445, -0.3176626, 
    -0.106027,
  // z(79, 0-99)
    0.1023834, 0.306746, 0.5098981, 0.7110379, 0.9093715, 1.104116, 1.294504, 
    1.479782, 1.65922, 1.832111, 1.997771, 2.155546, 2.304815, 2.444987, 
    2.57551, 2.695869, 2.805589, 2.904236, 2.991421, 3.066801, 3.130077, 
    3.181001, 3.21937, 3.245034, 3.257892, 3.257892, 3.245034, 3.21937, 
    3.181001, 3.130077, 3.066801, 2.991421, 2.904236, 2.805589, 2.695869, 
    2.57551, 2.444987, 2.304815, 2.155546, 1.997771, 1.832111, 1.65922, 
    1.479782, 1.294504, 1.104116, 0.9093715, 0.7110379, 0.5098981, 0.306746, 
    0.1023834, -0.1023834, -0.306746, -0.5098981, -0.7110379, -0.9093715, 
    -1.104116, -1.294504, -1.479782, -1.65922, -1.832111, -1.997771, 
    -2.155546, -2.304815, -2.444987, -2.57551, -2.695869, -2.805589, 
    -2.904236, -2.991421, -3.066801, -3.130077, -3.181001, -3.21937, 
    -3.245034, -3.257892, -3.257892, -3.245034, -3.21937, -3.181001, 
    -3.130077, -3.066801, -2.991421, -2.904236, -2.805589, -2.695869, 
    -2.57551, -2.444987, -2.304815, -2.155546, -1.997771, -1.832111, 
    -1.65922, -1.479782, -1.294504, -1.104116, -0.9093715, -0.7110379, 
    -0.5098981, -0.306746, -0.1023834,
  // z(80, 0-99)
    0.09861408, 0.295453, 0.491126, 0.6848607, 0.8758926, 1.063468, 1.246846, 
    1.425303, 1.598135, 1.764661, 1.924222, 2.076189, 2.219962, 2.354974, 
    2.480692, 2.596619, 2.7023, 2.797315, 2.881291, 2.953895, 3.014842, 
    3.063891, 3.100847, 3.125567, 3.137951, 3.137951, 3.125567, 3.100847, 
    3.063891, 3.014842, 2.953895, 2.881291, 2.797315, 2.7023, 2.596619, 
    2.480692, 2.354974, 2.219962, 2.076189, 1.924222, 1.764661, 1.598135, 
    1.425303, 1.246846, 1.063468, 0.8758926, 0.6848607, 0.491126, 0.295453, 
    0.09861408, -0.09861408, -0.295453, -0.491126, -0.6848607, -0.8758926, 
    -1.063468, -1.246846, -1.425303, -1.598135, -1.764661, -1.924222, 
    -2.076189, -2.219962, -2.354974, -2.480692, -2.596619, -2.7023, 
    -2.797315, -2.881291, -2.953895, -3.014842, -3.063891, -3.100847, 
    -3.125567, -3.137951, -3.137951, -3.125567, -3.100847, -3.063891, 
    -3.014842, -2.953895, -2.881291, -2.797315, -2.7023, -2.596619, 
    -2.480692, -2.354974, -2.219962, -2.076189, -1.924222, -1.764661, 
    -1.598135, -1.425303, -1.246846, -1.063468, -0.8758926, -0.6848607, 
    -0.491126, -0.295453, -0.09861408,
  // z(81, 0-99)
    0.09471914, 0.2837836, 0.4717281, 0.6578109, 0.8412977, 1.021464, 
    1.197599, 1.369008, 1.535014, 1.694962, 1.848221, 1.994186, 2.132281, 
    2.26196, 2.382712, 2.494061, 2.595567, 2.68683, 2.767489, 2.837226, 
    2.895766, 2.942877, 2.978374, 3.002117, 3.014012, 3.014012, 3.002117, 
    2.978374, 2.942877, 2.895766, 2.837226, 2.767489, 2.68683, 2.595567, 
    2.494061, 2.382712, 2.26196, 2.132281, 1.994186, 1.848221, 1.694962, 
    1.535014, 1.369008, 1.197599, 1.021464, 0.8412977, 0.6578109, 0.4717281, 
    0.2837836, 0.09471914, -0.09471914, -0.2837836, -0.4717281, -0.6578109, 
    -0.8412977, -1.021464, -1.197599, -1.369008, -1.535014, -1.694962, 
    -1.848221, -1.994186, -2.132281, -2.26196, -2.382712, -2.494061, 
    -2.595567, -2.68683, -2.767489, -2.837226, -2.895766, -2.942877, 
    -2.978374, -3.002117, -3.014012, -3.014012, -3.002117, -2.978374, 
    -2.942877, -2.895766, -2.837226, -2.767489, -2.68683, -2.595567, 
    -2.494061, -2.382712, -2.26196, -2.132281, -1.994186, -1.848221, 
    -1.694962, -1.535014, -1.369008, -1.197599, -1.021464, -0.8412977, 
    -0.6578109, -0.4717281, -0.2837836, -0.09471914,
  // z(82, 0-99)
    0.09069857, 0.2717378, 0.4517045, 0.6298886, 0.8055868, 0.9781057, 
    1.146765, 1.310898, 1.469857, 1.623016, 1.769769, 1.909538, 2.041771, 
    2.165946, 2.281573, 2.388195, 2.485393, 2.572781, 2.650017, 2.716793, 
    2.772848, 2.81796, 2.85195, 2.874685, 2.886075, 2.886075, 2.874685, 
    2.85195, 2.81796, 2.772848, 2.716793, 2.650017, 2.572781, 2.485393, 
    2.388195, 2.281573, 2.165946, 2.041771, 1.909538, 1.769769, 1.623016, 
    1.469857, 1.310898, 1.146765, 0.9781057, 0.8055868, 0.6298886, 0.4517045, 
    0.2717378, 0.09069857, -0.09069857, -0.2717378, -0.4517045, -0.6298886, 
    -0.8055868, -0.9781057, -1.146765, -1.310898, -1.469857, -1.623016, 
    -1.769769, -1.909538, -2.041771, -2.165946, -2.281573, -2.388195, 
    -2.485393, -2.572781, -2.650017, -2.716793, -2.772848, -2.81796, 
    -2.85195, -2.874685, -2.886075, -2.886075, -2.874685, -2.85195, -2.81796, 
    -2.772848, -2.716793, -2.650017, -2.572781, -2.485393, -2.388195, 
    -2.281573, -2.165946, -2.041771, -1.909538, -1.769769, -1.623016, 
    -1.469857, -1.310898, -1.146765, -0.9781057, -0.8055868, -0.6298886, 
    -0.4517045, -0.2717378, -0.09069857,
  // z(83, 0-99)
    0.08655234, 0.2593155, 0.4310552, 0.6010937, 0.76876, 0.9333923, 
    1.094341, 1.250971, 1.402664, 1.548821, 1.688865, 1.822245, 1.948433, 
    2.066931, 2.177272, 2.279021, 2.371775, 2.455168, 2.528873, 2.592597, 
    2.646089, 2.689139, 2.721575, 2.743271, 2.75414, 2.75414, 2.743271, 
    2.721575, 2.689139, 2.646089, 2.592597, 2.528873, 2.455168, 2.371775, 
    2.279021, 2.177272, 2.066931, 1.948433, 1.822245, 1.688865, 1.548821, 
    1.402664, 1.250971, 1.094341, 0.9333923, 0.76876, 0.6010937, 0.4310552, 
    0.2593155, 0.08655234, -0.08655234, -0.2593155, -0.4310552, -0.6010937, 
    -0.76876, -0.9333923, -1.094341, -1.250971, -1.402664, -1.548821, 
    -1.688865, -1.822245, -1.948433, -2.066931, -2.177272, -2.279021, 
    -2.371775, -2.455168, -2.528873, -2.592597, -2.646089, -2.689139, 
    -2.721575, -2.743271, -2.75414, -2.75414, -2.743271, -2.721575, 
    -2.689139, -2.646089, -2.592597, -2.528873, -2.455168, -2.371775, 
    -2.279021, -2.177272, -2.066931, -1.948433, -1.822245, -1.688865, 
    -1.548821, -1.402664, -1.250971, -1.094341, -0.9333923, -0.76876, 
    -0.6010937, -0.4310552, -0.2593155, -0.08655234,
  // z(84, 0-99)
    0.08228049, 0.2465167, 0.4097801, 0.5714262, 0.7308172, 0.887324, 
    1.040329, 1.189228, 1.333434, 1.472377, 1.60551, 1.732306, 1.852266, 
    1.964916, 2.069811, 2.166538, 2.254714, 2.333992, 2.404058, 2.464637, 
    2.515489, 2.556414, 2.58725, 2.607875, 2.618207, 2.618207, 2.607875, 
    2.58725, 2.556414, 2.515489, 2.464637, 2.404058, 2.333992, 2.254714, 
    2.166538, 2.069811, 1.964916, 1.852266, 1.732306, 1.60551, 1.472377, 
    1.333434, 1.189228, 1.040329, 0.887324, 0.7308172, 0.5714262, 0.4097801, 
    0.2465167, 0.08228049, -0.08228049, -0.2465167, -0.4097801, -0.5714262, 
    -0.7308172, -0.887324, -1.040329, -1.189228, -1.333434, -1.472377, 
    -1.60551, -1.732306, -1.852266, -1.964916, -2.069811, -2.166538, 
    -2.254714, -2.333992, -2.404058, -2.464637, -2.515489, -2.556414, 
    -2.58725, -2.607875, -2.618207, -2.618207, -2.607875, -2.58725, 
    -2.556414, -2.515489, -2.464637, -2.404058, -2.333992, -2.254714, 
    -2.166538, -2.069811, -1.964916, -1.852266, -1.732306, -1.60551, 
    -1.472377, -1.333434, -1.189228, -1.040329, -0.887324, -0.7308172, 
    -0.5714262, -0.4097801, -0.2465167, -0.08228049,
  // z(85, 0-99)
    0.07788298, 0.2333416, 0.3878793, 0.5408862, 0.6917585, 0.8399007, 
    0.9847282, 1.125669, 1.262168, 1.393686, 1.519703, 1.639723, 1.753271, 
    1.8599, 1.959189, 2.050746, 2.13421, 2.209251, 2.275573, 2.332914, 
    2.381048, 2.419785, 2.448973, 2.468496, 2.478276, 2.478276, 2.468496, 
    2.448973, 2.419785, 2.381048, 2.332914, 2.275573, 2.209251, 2.13421, 
    2.050746, 1.959189, 1.8599, 1.753271, 1.639723, 1.519703, 1.393686, 
    1.262168, 1.125669, 0.9847282, 0.8399007, 0.6917585, 0.5408862, 
    0.3878793, 0.2333416, 0.07788298, -0.07788298, -0.2333416, -0.3878793, 
    -0.5408862, -0.6917585, -0.8399007, -0.9847282, -1.125669, -1.262168, 
    -1.393686, -1.519703, -1.639723, -1.753271, -1.8599, -1.959189, 
    -2.050746, -2.13421, -2.209251, -2.275573, -2.332914, -2.381048, 
    -2.419785, -2.448973, -2.468496, -2.478276, -2.478276, -2.468496, 
    -2.448973, -2.419785, -2.381048, -2.332914, -2.275573, -2.209251, 
    -2.13421, -2.050746, -1.959189, -1.8599, -1.753271, -1.639723, -1.519703, 
    -1.393686, -1.262168, -1.125669, -0.9847282, -0.8399007, -0.6917585, 
    -0.5408862, -0.3878793, -0.2333416, -0.07788298,
  // z(86, 0-99)
    0.07335982, 0.21979, 0.3653527, 0.5094736, 0.6515837, 0.7911224, 
    0.9275389, 1.060295, 1.188866, 1.312746, 1.431444, 1.544494, 1.651448, 
    1.751884, 1.845407, 1.931647, 2.010263, 2.080946, 2.143416, 2.197427, 
    2.242766, 2.279253, 2.306746, 2.325135, 2.334347, 2.334347, 2.325135, 
    2.306746, 2.279253, 2.242766, 2.197427, 2.143416, 2.080946, 2.010263, 
    1.931647, 1.845407, 1.751884, 1.651448, 1.544494, 1.431444, 1.312746, 
    1.188866, 1.060295, 0.9275389, 0.7911224, 0.6515837, 0.5094736, 
    0.3653527, 0.21979, 0.07335982, -0.07335982, -0.21979, -0.3653527, 
    -0.5094736, -0.6515837, -0.7911224, -0.9275389, -1.060295, -1.188866, 
    -1.312746, -1.431444, -1.544494, -1.651448, -1.751884, -1.845407, 
    -1.931647, -2.010263, -2.080946, -2.143416, -2.197427, -2.242766, 
    -2.279253, -2.306746, -2.325135, -2.334347, -2.334347, -2.325135, 
    -2.306746, -2.279253, -2.242766, -2.197427, -2.143416, -2.080946, 
    -2.010263, -1.931647, -1.845407, -1.751884, -1.651448, -1.544494, 
    -1.431444, -1.312746, -1.188866, -1.060295, -0.9275389, -0.7911224, 
    -0.6515837, -0.5094736, -0.3653527, -0.21979, -0.07335982,
  // z(87, 0-99)
    0.06871103, 0.2058619, 0.3422004, 0.4771883, 0.610293, 0.7409892, 
    0.868761, 0.9931042, 1.113528, 1.229557, 1.340734, 1.44662, 1.546796, 
    1.640868, 1.728464, 1.809239, 1.882873, 1.949077, 2.007588, 2.058177, 
    2.100642, 2.134818, 2.160568, 2.177792, 2.186421, 2.186421, 2.177792, 
    2.160568, 2.134818, 2.100642, 2.058177, 2.007588, 1.949077, 1.882873, 
    1.809239, 1.728464, 1.640868, 1.546796, 1.44662, 1.340734, 1.229557, 
    1.113528, 0.9931042, 0.868761, 0.7409892, 0.610293, 0.4771883, 0.3422004, 
    0.2058619, 0.06871103, -0.06871103, -0.2058619, -0.3422004, -0.4771883, 
    -0.610293, -0.7409892, -0.868761, -0.9931042, -1.113528, -1.229557, 
    -1.340734, -1.44662, -1.546796, -1.640868, -1.728464, -1.809239, 
    -1.882873, -1.949077, -2.007588, -2.058177, -2.100642, -2.134818, 
    -2.160568, -2.177792, -2.186421, -2.186421, -2.177792, -2.160568, 
    -2.134818, -2.100642, -2.058177, -2.007588, -1.949077, -1.882873, 
    -1.809239, -1.728464, -1.640868, -1.546796, -1.44662, -1.340734, 
    -1.229557, -1.113528, -0.9931042, -0.868761, -0.7409892, -0.610293, 
    -0.4771883, -0.3422004, -0.2058619, -0.06871103,
  // z(88, 0-99)
    0.0639366, 0.1915575, 0.3184223, 0.4440306, 0.5678864, 0.689501, 
    0.8083946, 0.9240977, 1.036154, 1.144121, 1.247572, 1.3461, 1.439316, 
    1.526851, 1.608361, 1.683522, 1.75204, 1.813644, 1.86809, 1.915163, 
    1.954678, 1.986479, 2.01044, 2.026466, 2.034496, 2.034496, 2.026466, 
    2.01044, 1.986479, 1.954678, 1.915163, 1.86809, 1.813644, 1.75204, 
    1.683522, 1.608361, 1.526851, 1.439316, 1.3461, 1.247572, 1.144121, 
    1.036154, 0.9240977, 0.8083946, 0.689501, 0.5678864, 0.4440306, 
    0.3184223, 0.1915575, 0.0639366, -0.0639366, -0.1915575, -0.3184223, 
    -0.4440306, -0.5678864, -0.689501, -0.8083946, -0.9240977, -1.036154, 
    -1.144121, -1.247572, -1.3461, -1.439316, -1.526851, -1.608361, 
    -1.683522, -1.75204, -1.813644, -1.86809, -1.915163, -1.954678, 
    -1.986479, -2.01044, -2.026466, -2.034496, -2.034496, -2.026466, 
    -2.01044, -1.986479, -1.954678, -1.915163, -1.86809, -1.813644, -1.75204, 
    -1.683522, -1.608361, -1.526851, -1.439316, -1.3461, -1.247572, 
    -1.144121, -1.036154, -0.9240977, -0.8083946, -0.689501, -0.5678864, 
    -0.4440306, -0.3184223, -0.1915575, -0.0639366,
  // z(89, 0-99)
    0.05903652, 0.1768766, 0.2940186, 0.4100002, 0.5243638, 0.6366579, 
    0.7464395, 0.8532751, 0.9567434, 1.056436, 1.151959, 1.242936, 1.329007, 
    1.409834, 1.485096, 1.554498, 1.617765, 1.674647, 1.72492, 1.768385, 
    1.804872, 1.834236, 1.85636, 1.871159, 1.878573, 1.878573, 1.871159, 
    1.85636, 1.834236, 1.804872, 1.768385, 1.72492, 1.674647, 1.617765, 
    1.554498, 1.485096, 1.409834, 1.329007, 1.242936, 1.151959, 1.056436, 
    0.9567434, 0.8532751, 0.7464395, 0.6366579, 0.5243638, 0.4100002, 
    0.2940186, 0.1768766, 0.05903652, -0.05903652, -0.1768766, -0.2940186, 
    -0.4100002, -0.5243638, -0.6366579, -0.7464395, -0.8532751, -0.9567434, 
    -1.056436, -1.151959, -1.242936, -1.329007, -1.409834, -1.485096, 
    -1.554498, -1.617765, -1.674647, -1.72492, -1.768385, -1.804872, 
    -1.834236, -1.85636, -1.871159, -1.878573, -1.878573, -1.871159, 
    -1.85636, -1.834236, -1.804872, -1.768385, -1.72492, -1.674647, 
    -1.617765, -1.554498, -1.485096, -1.409834, -1.329007, -1.242936, 
    -1.151959, -1.056436, -0.9567434, -0.8532751, -0.7464395, -0.6366579, 
    -0.5243638, -0.4100002, -0.2940186, -0.1768766, -0.05903652,
  // z(90, 0-99)
    0.0540108, 0.1618192, 0.2689891, 0.3750973, 0.4797252, 0.5824599, 
    0.6828958, 0.7806367, 0.8752967, 0.9665024, 1.053894, 1.137126, 1.21587, 
    1.289816, 1.358672, 1.422165, 1.480046, 1.532086, 1.578079, 1.617844, 
    1.651225, 1.678089, 1.69833, 1.711869, 1.718652, 1.718652, 1.711869, 
    1.69833, 1.678089, 1.651225, 1.617844, 1.578079, 1.532086, 1.480046, 
    1.422165, 1.358672, 1.289816, 1.21587, 1.137126, 1.053894, 0.9665024, 
    0.8752967, 0.7806367, 0.6828958, 0.5824599, 0.4797252, 0.3750973, 
    0.2689891, 0.1618192, 0.0540108, -0.0540108, -0.1618192, -0.2689891, 
    -0.3750973, -0.4797252, -0.5824599, -0.6828958, -0.7806367, -0.8752967, 
    -0.9665024, -1.053894, -1.137126, -1.21587, -1.289816, -1.358672, 
    -1.422165, -1.480046, -1.532086, -1.578079, -1.617844, -1.651225, 
    -1.678089, -1.69833, -1.711869, -1.718652, -1.718652, -1.711869, 
    -1.69833, -1.678089, -1.651225, -1.617844, -1.578079, -1.532086, 
    -1.480046, -1.422165, -1.358672, -1.289816, -1.21587, -1.137126, 
    -1.053894, -0.9665024, -0.8752967, -0.7806367, -0.6828958, -0.5824599, 
    -0.4797252, -0.3750973, -0.2689891, -0.1618192, -0.0540108,
  // z(91, 0-99)
    0.04885944, 0.1463855, 0.2433338, 0.3393218, 0.4339707, 0.5269068, 
    0.6177635, 0.7061822, 0.7918139, 0.8743207, 0.9533769, 1.028671, 
    1.099905, 1.166798, 1.229086, 1.286524, 1.338884, 1.385961, 1.427567, 
    1.46354, 1.493737, 1.518039, 1.536349, 1.548597, 1.554732, 1.554732, 
    1.548597, 1.536349, 1.518039, 1.493737, 1.46354, 1.427567, 1.385961, 
    1.338884, 1.286524, 1.229086, 1.166798, 1.099905, 1.028671, 0.9533769, 
    0.8743207, 0.7918139, 0.7061822, 0.6177635, 0.5269068, 0.4339707, 
    0.3393218, 0.2433338, 0.1463855, 0.04885944, -0.04885944, -0.1463855, 
    -0.2433338, -0.3393218, -0.4339707, -0.5269068, -0.6177635, -0.7061822, 
    -0.7918139, -0.8743207, -0.9533769, -1.028671, -1.099905, -1.166798, 
    -1.229086, -1.286524, -1.338884, -1.385961, -1.427567, -1.46354, 
    -1.493737, -1.518039, -1.536349, -1.548597, -1.554732, -1.554732, 
    -1.548597, -1.536349, -1.518039, -1.493737, -1.46354, -1.427567, 
    -1.385961, -1.338884, -1.286524, -1.229086, -1.166798, -1.099905, 
    -1.028671, -0.9533769, -0.8743207, -0.7918139, -0.7061822, -0.6177635, 
    -0.5269068, -0.4339707, -0.3393218, -0.2433338, -0.1463855, -0.04885944,
  // z(92, 0-99)
    0.04358243, 0.1305753, 0.2170528, 0.3026738, 0.3871002, 0.4699989, 
    0.5510427, 0.6299118, 0.706295, 0.7798907, 0.8504086, 0.9175702, 
    0.9811106, 1.040779, 1.09634, 1.147574, 1.19428, 1.236272, 1.273385, 
    1.305472, 1.332407, 1.354084, 1.370418, 1.381342, 1.386815, 1.386815, 
    1.381342, 1.370418, 1.354084, 1.332407, 1.305472, 1.273385, 1.236272, 
    1.19428, 1.147574, 1.09634, 1.040779, 0.9811106, 0.9175702, 0.8504086, 
    0.7798907, 0.706295, 0.6299118, 0.5510427, 0.4699989, 0.3871002, 
    0.3026738, 0.2170528, 0.1305753, 0.04358243, -0.04358243, -0.1305753, 
    -0.2170528, -0.3026738, -0.3871002, -0.4699989, -0.5510427, -0.6299118, 
    -0.706295, -0.7798907, -0.8504086, -0.9175702, -0.9811106, -1.040779, 
    -1.09634, -1.147574, -1.19428, -1.236272, -1.273385, -1.305472, 
    -1.332407, -1.354084, -1.370418, -1.381342, -1.386815, -1.386815, 
    -1.381342, -1.370418, -1.354084, -1.332407, -1.305472, -1.273385, 
    -1.236272, -1.19428, -1.147574, -1.09634, -1.040779, -0.9811106, 
    -0.9175702, -0.8504086, -0.7798907, -0.706295, -0.6299118, -0.5510427, 
    -0.4699989, -0.3871002, -0.3026738, -0.2170528, -0.1305753, -0.04358243,
  // z(93, 0-99)
    0.03817978, 0.1143887, 0.1901461, 0.2651531, 0.3391137, 0.411736, 
    0.4827332, 0.5518255, 0.6187398, 0.6832123, 0.7449885, 0.8038245, 
    0.8594883, 0.91176, 0.9604334, 1.005316, 1.046232, 1.083018, 1.115531, 
    1.143641, 1.167237, 1.186227, 1.200535, 1.210106, 1.2149, 1.2149, 
    1.210106, 1.200535, 1.186227, 1.167237, 1.143641, 1.115531, 1.083018, 
    1.046232, 1.005316, 0.9604334, 0.91176, 0.8594883, 0.8038245, 0.7449885, 
    0.6832123, 0.6187398, 0.5518255, 0.4827332, 0.411736, 0.3391137, 
    0.2651531, 0.1901461, 0.1143887, 0.03817978, -0.03817978, -0.1143887, 
    -0.1901461, -0.2651531, -0.3391137, -0.411736, -0.4827332, -0.5518255, 
    -0.6187398, -0.6832123, -0.7449885, -0.8038245, -0.8594883, -0.91176, 
    -0.9604334, -1.005316, -1.046232, -1.083018, -1.115531, -1.143641, 
    -1.167237, -1.186227, -1.200535, -1.210106, -1.2149, -1.2149, -1.210106, 
    -1.200535, -1.186227, -1.167237, -1.143641, -1.115531, -1.083018, 
    -1.046232, -1.005316, -0.9604334, -0.91176, -0.8594883, -0.8038245, 
    -0.7449885, -0.6832123, -0.6187398, -0.5518255, -0.4827332, -0.411736, 
    -0.3391137, -0.2651531, -0.1901461, -0.1143887, -0.03817978,
  // z(94, 0-99)
    0.03265148, 0.09782559, 0.1626136, 0.2267599, 0.2900113, 0.3521181, 
    0.4128352, 0.4719231, 0.5291486, 0.5842857, 0.6371169, 0.6874337, 
    0.7350375, 0.7797405, 0.8213661, 0.8597503, 0.8947414, 0.9262013, 
    0.954006, 0.9780456, 0.9982253, 1.014465, 1.026702, 1.034887, 1.038987, 
    1.038987, 1.034887, 1.026702, 1.014465, 0.9982253, 0.9780456, 0.954006, 
    0.9262013, 0.8947414, 0.8597503, 0.8213661, 0.7797405, 0.7350375, 
    0.6874337, 0.6371169, 0.5842857, 0.5291486, 0.4719231, 0.4128352, 
    0.3521181, 0.2900113, 0.2267599, 0.1626136, 0.09782559, 0.03265148, 
    -0.03265148, -0.09782559, -0.1626136, -0.2267599, -0.2900113, -0.3521181, 
    -0.4128352, -0.4719231, -0.5291486, -0.5842857, -0.6371169, -0.6874337, 
    -0.7350375, -0.7797405, -0.8213661, -0.8597503, -0.8947414, -0.9262013, 
    -0.954006, -0.9780456, -0.9982253, -1.014465, -1.026702, -1.034887, 
    -1.038987, -1.038987, -1.034887, -1.026702, -1.014465, -0.9982253, 
    -0.9780456, -0.954006, -0.9262013, -0.8947414, -0.8597503, -0.8213661, 
    -0.7797405, -0.7350375, -0.6874337, -0.6371169, -0.5842857, -0.5291486, 
    -0.4719231, -0.4128352, -0.3521181, -0.2900113, -0.2267599, -0.1626136, 
    -0.09782559, -0.03265148,
  // z(95, 0-99)
    0.02699755, 0.0808861, 0.1344554, 0.1874941, 0.2397929, 0.2911452, 
    0.3413486, 0.3902048, 0.4375211, 0.4831107, 0.5267936, 0.5683975, 
    0.6077583, 0.6447204, 0.6791382, 0.7108757, 0.7398078, 0.7658201, 
    0.7888101, 0.808687, 0.8253724, 0.8388004, 0.8489181, 0.8556855, 
    0.8590759, 0.8590759, 0.8556855, 0.8489181, 0.8388004, 0.8253724, 
    0.808687, 0.7888101, 0.7658201, 0.7398078, 0.7108757, 0.6791382, 
    0.6447204, 0.6077583, 0.5683975, 0.5267936, 0.4831107, 0.4375211, 
    0.3902048, 0.3413486, 0.2911452, 0.2397929, 0.1874941, 0.1344554, 
    0.0808861, 0.02699755, -0.02699755, -0.0808861, -0.1344554, -0.1874941, 
    -0.2397929, -0.2911452, -0.3413486, -0.3902048, -0.4375211, -0.4831107, 
    -0.5267936, -0.5683975, -0.6077583, -0.6447204, -0.6791382, -0.7108757, 
    -0.7398078, -0.7658201, -0.7888101, -0.808687, -0.8253724, -0.8388004, 
    -0.8489181, -0.8556855, -0.8590759, -0.8590759, -0.8556855, -0.8489181, 
    -0.8388004, -0.8253724, -0.808687, -0.7888101, -0.7658201, -0.7398078, 
    -0.7108757, -0.6791382, -0.6447204, -0.6077583, -0.5683975, -0.5267936, 
    -0.4831107, -0.4375211, -0.3902048, -0.3413486, -0.2911452, -0.2397929, 
    -0.1874941, -0.1344554, -0.0808861, -0.02699755,
  // z(96, 0-99)
    0.02121797, 0.06357016, 0.1056715, 0.1473558, 0.1884585, 0.2288175, 
    0.2682734, 0.3066706, 0.3438575, 0.3796873, 0.4140187, 0.4467162, 
    0.4776506, 0.5067, 0.5337497, 0.5586929, 0.5814312, 0.6018749, 0.6199433, 
    0.635565, 0.6486784, 0.6592318, 0.6671835, 0.6725021, 0.6751667, 
    0.6751667, 0.6725021, 0.6671835, 0.6592318, 0.6486784, 0.635565, 
    0.6199433, 0.6018749, 0.5814312, 0.5586929, 0.5337497, 0.5067, 0.4776506, 
    0.4467162, 0.4140187, 0.3796873, 0.3438575, 0.3066706, 0.2682734, 
    0.2288175, 0.1884585, 0.1473558, 0.1056715, 0.06357016, 0.02121797, 
    -0.02121797, -0.06357016, -0.1056715, -0.1473558, -0.1884585, -0.2288175, 
    -0.2682734, -0.3066706, -0.3438575, -0.3796873, -0.4140187, -0.4467162, 
    -0.4776506, -0.5067, -0.5337497, -0.5586929, -0.5814312, -0.6018749, 
    -0.6199433, -0.635565, -0.6486784, -0.6592318, -0.6671835, -0.6725021, 
    -0.6751667, -0.6751667, -0.6725021, -0.6671835, -0.6592318, -0.6486784, 
    -0.635565, -0.6199433, -0.6018749, -0.5814312, -0.5586929, -0.5337497, 
    -0.5067, -0.4776506, -0.4467162, -0.4140187, -0.3796873, -0.3438575, 
    -0.3066706, -0.2682734, -0.2288175, -0.1884585, -0.1473558, -0.1056715, 
    -0.06357016, -0.02121797,
  // z(97, 0-99)
    0.01531275, 0.0458778, 0.0762618, 0.1063448, 0.1360082, 0.1651347, 
    0.1936096, 0.2213204, 0.2481577, 0.2740156, 0.2987922, 0.3223895, 
    0.3447146, 0.3656791, 0.3852006, 0.4032018, 0.4196118, 0.4343657, 
    0.4474054, 0.4586794, 0.4681432, 0.4757594, 0.4814981, 0.4853365, 
    0.4872594, 0.4872594, 0.4853365, 0.4814981, 0.4757594, 0.4681432, 
    0.4586794, 0.4474054, 0.4343657, 0.4196118, 0.4032018, 0.3852006, 
    0.3656791, 0.3447146, 0.3223895, 0.2987922, 0.2740156, 0.2481577, 
    0.2213204, 0.1936096, 0.1651347, 0.1360082, 0.1063448, 0.0762618, 
    0.0458778, 0.01531275, -0.01531275, -0.0458778, -0.0762618, -0.1063448, 
    -0.1360082, -0.1651347, -0.1936096, -0.2213204, -0.2481577, -0.2740156, 
    -0.2987922, -0.3223895, -0.3447146, -0.3656791, -0.3852006, -0.4032018, 
    -0.4196118, -0.4343657, -0.4474054, -0.4586794, -0.4681432, -0.4757594, 
    -0.4814981, -0.4853365, -0.4872594, -0.4872594, -0.4853365, -0.4814981, 
    -0.4757594, -0.4681432, -0.4586794, -0.4474054, -0.4343657, -0.4196118, 
    -0.4032018, -0.3852006, -0.3656791, -0.3447146, -0.3223895, -0.2987922, 
    -0.2740156, -0.2481577, -0.2213204, -0.1936096, -0.1651347, -0.1360082, 
    -0.1063448, -0.0762618, -0.0458778, -0.01531275,
  // z(98, 0-99)
    0.009281879, 0.02780901, 0.04622639, 0.06446133, 0.08244187, 0.1000971, 
    0.1173572, 0.1341542, 0.1504217, 0.1660956, 0.181114, 0.1954177, 
    0.2089501, 0.2216578, 0.2334908, 0.2444023, 0.2543493, 0.2632924, 
    0.2711965, 0.2780303, 0.2837668, 0.2883834, 0.2918619, 0.2941886, 
    0.2953542, 0.2953542, 0.2941886, 0.2918619, 0.2883834, 0.2837668, 
    0.2780303, 0.2711965, 0.2632924, 0.2543493, 0.2444023, 0.2334908, 
    0.2216578, 0.2089501, 0.1954177, 0.181114, 0.1660956, 0.1504217, 
    0.1341542, 0.1173572, 0.1000971, 0.08244187, 0.06446133, 0.04622639, 
    0.02780901, 0.009281879, -0.009281879, -0.02780901, -0.04622639, 
    -0.06446133, -0.08244187, -0.1000971, -0.1173572, -0.1341542, -0.1504217, 
    -0.1660956, -0.181114, -0.1954177, -0.2089501, -0.2216578, -0.2334908, 
    -0.2444023, -0.2543493, -0.2632924, -0.2711965, -0.2780303, -0.2837668, 
    -0.2883834, -0.2918619, -0.2941886, -0.2953542, -0.2953542, -0.2941886, 
    -0.2918619, -0.2883834, -0.2837668, -0.2780303, -0.2711965, -0.2632924, 
    -0.2543493, -0.2444023, -0.2334908, -0.2216578, -0.2089501, -0.1954177, 
    -0.181114, -0.1660956, -0.1504217, -0.1341542, -0.1173572, -0.1000971, 
    -0.08244187, -0.06446133, -0.04622639, -0.02780901, -0.009281879,
  // z(99, 0-99)
    0.00312537, 0.009363777, 0.01556523, 0.02170525, 0.02775962, 0.03370442, 
    0.03951621, 0.04517205, 0.05064962, 0.0559273, 0.06098425, 0.06580053, 
    0.07035712, 0.07463605, 0.07862043, 0.08229452, 0.08564384, 0.08865515, 
    0.09131659, 0.09361763, 0.09554922, 0.09710371, 0.09827499, 0.09905841, 
    0.0994509, 0.0994509, 0.09905841, 0.09827499, 0.09710371, 0.09554922, 
    0.09361763, 0.09131659, 0.08865515, 0.08564384, 0.08229452, 0.07862043, 
    0.07463605, 0.07035712, 0.06580053, 0.06098425, 0.0559273, 0.05064962, 
    0.04517205, 0.03951621, 0.03370442, 0.02775962, 0.02170525, 0.01556523, 
    0.009363777, 0.00312537, -0.00312537, -0.009363777, -0.01556523, 
    -0.02170525, -0.02775962, -0.03370442, -0.03951621, -0.04517205, 
    -0.05064962, -0.0559273, -0.06098425, -0.06580053, -0.07035712, 
    -0.07463605, -0.07862043, -0.08229452, -0.08564384, -0.08865515, 
    -0.09131659, -0.09361763, -0.09554922, -0.09710371, -0.09827499, 
    -0.09905841, -0.0994509, -0.0994509, -0.09905841, -0.09827499, 
    -0.09710371, -0.09554922, -0.09361763, -0.09131659, -0.08865515, 
    -0.08564384, -0.08229452, -0.07862043, -0.07463605, -0.07035712, 
    -0.06580053, -0.06098425, -0.0559273, -0.05064962, -0.04517205, 
    -0.03951621, -0.03370442, -0.02775962, -0.02170525, -0.01556523, 
    -0.009363777, -0.00312537 ;
}
