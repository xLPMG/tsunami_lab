netcdf tsunamiNetCdf {
dimensions:
	x = 10 ;
	y = 10 ;
variables:
	float x(x) ;
		x:units = "meters" ;
		x:axis = "X" ;
	float y(y) ;
		y:units = "meters" ;
		y:axis = "Y" ;
	float bathymetry(x, y) ;
        bathymetry:units = "meters" ;
data:

 x = 0, 1, 2, 3, 4, 5, 6, 7, 8, 9 ;

 y = 0, 1, 2, 3, 4, 5, 6, 7, 8, 9 ;

 bathymetry =
  // bathymetry(0, 0-9)
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1,
  // bathymetry(1, 0-9)
    -2, -2, -2, -2, -2, -2, -2, -2, -2, -2,
  // bathymetry(2, 0-9)
    -3, -3, -3, -3, -3, -3, -3, -3, -3, -3,
  // bathymetry(3, 0-9)
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1,
  // bathymetry(4, 0-9)
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1,
  // bathymetry(5, 0-9)
    -1, -1, 23, -1, -1, -1, -1, -1, -1, -1,
  // bathymetry(6, 0-9)
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1,
  // bathymetry(7, 0-9)
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1,
  // bathymetry(8, 0-9)
    -1, -1, -1, -1, -1, -1, 99, -1, -1, -1,
  // bathymetry(9, 0-9)
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1 ;
}