netcdf netCdfTest {
dimensions:
	time = UNLIMITED ; // (1 currently)
	x = 10 ;
	y = 10 ;
variables:
	float time(time) ;
		time:units = "seconds since the earthquake event" ;
	float x(x) ;
		x:units = "meters" ;
		x:axis = "X" ;
	float y(y) ;
		y:units = "meters" ;
		y:axis = "Y" ;
	float height(time, x, y) ;
		height:units = "meters" ;
	float totalHeight(time, x, y) ;
		totalHeight:units = "meters" ;
	float bathymetry(x, y) ;
	float momentumX(time, x, y) ;
		momentumX:units = "square meters per second" ;
	float momentumY(time, x, y) ;
		momentumY:units = "square meters per second" ;
data:

 time = 0 ;

 x = 0.5, 1.5, 2.5, 3.5, 4.5, 5.5, 6.5, 7.5, 8.5, 9.5 ;

 y = 0.5, 1.5, 2.5, 3.5, 4.5, 5.5, 6.5, 7.5, 8.5, 9.5 ;

 height =
  // height(0,0, 0-9)
    -100, -200, -300, -400, -500, -600, -700, -800, -900, -1000,
  // height(0,1, 0-9)
    -100, -200, -300, -400, -500, -600, -700, -800, -900, -1000,
  // height(0,2, 0-9)
    -100, -200, -300, -400, -500, -600, -700, -800, -900, -1000,
  // height(0,3, 0-9)
    -100, -200, -300, -400, -500, -600, -700, -800, -900, -1000,
  // height(0,4, 0-9)
    -100, -200, -300, -400, -500, -600, -700, -800, -900, -1000,
  // height(0,5, 0-9)
    -100, -200, -300, -400, -500, -600, -700, -800, -900, -1000,
  // height(0,6, 0-9)
    -100, -200, -300, -400, -500, -600, -700, -800, -900, -1000,
  // height(0,7, 0-9)
    -100, -200, -300, -400, -500, -600, -700, -800, -900, -1000,
  // height(0,8, 0-9)
    -100, -200, -300, -400, -500, -600, -700, -800, -900, -1000,
  // height(0,9, 0-9)
    -100, -200, -300, -400, -500, -600, -700, -800, -900, -1000 ;

 totalHeight =
  // totalHeight(0,0, 0-9)
    -100, -200, -300, -400, -500, -600, -700, -800, -900, -1000,
  // totalHeight(0,1, 0-9)
    -100, -200, -300, -400, -500, -600, -700, -800, -900, -1000,
  // totalHeight(0,2, 0-9)
    -100, -200, -300, -400, -500, -600, -700, -800, -900, -1000,
  // totalHeight(0,3, 0-9)
    -100, -200, -300, -400, -500, -600, -700, -800, -900, -1000,
  // totalHeight(0,4, 0-9)
    -100, -200, -300, -400, -500, -600, -700, -800, -900, -1000,
  // totalHeight(0,5, 0-9)
    -100, -200, -300, -400, -500, -600, -700, -800, -900, -1000,
  // totalHeight(0,6, 0-9)
    -100, -200, -300, -400, -500, -600, -700, -800, -900, -1000,
  // totalHeight(0,7, 0-9)
    -100, -200, -300, -400, -500, -600, -700, -800, -900, -1000,
  // totalHeight(0,8, 0-9)
    -100, -200, -300, -400, -500, -600, -700, -800, -900, -1000,
  // totalHeight(0,9, 0-9)
    -100, -200, -300, -400, -500, -600, -700, -800, -900, -1000 ;

 bathymetry =
  // bathymetry(0, 0-9)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  // bathymetry(1, 0-9)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  // bathymetry(2, 0-9)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  // bathymetry(3, 0-9)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  // bathymetry(4, 0-9)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  // bathymetry(5, 0-9)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  // bathymetry(6, 0-9)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  // bathymetry(7, 0-9)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  // bathymetry(8, 0-9)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  // bathymetry(9, 0-9)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 momentumX =
  // momentumX(0,0, 0-9)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  // momentumX(0,1, 0-9)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  // momentumX(0,2, 0-9)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  // momentumX(0,3, 0-9)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  // momentumX(0,4, 0-9)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  // momentumX(0,5, 0-9)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  // momentumX(0,6, 0-9)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  // momentumX(0,7, 0-9)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  // momentumX(0,8, 0-9)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  // momentumX(0,9, 0-9)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 momentumY =
  // momentumY(0,0, 0-9)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  // momentumY(0,1, 0-9)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  // momentumY(0,2, 0-9)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  // momentumY(0,3, 0-9)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  // momentumY(0,4, 0-9)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  // momentumY(0,5, 0-9)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  // momentumY(0,6, 0-9)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  // momentumY(0,7, 0-9)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  // momentumY(0,8, 0-9)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  // momentumY(0,9, 0-9)
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;
}
